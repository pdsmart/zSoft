-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"b0",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"bf",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"ac",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"ab",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8f",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"90",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"91",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"92",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"90",
           386 => x"97",
           387 => x"90",
           388 => x"80",
           389 => x"bb",
           390 => x"ee",
           391 => x"90",
           392 => x"80",
           393 => x"bb",
           394 => x"f3",
           395 => x"90",
           396 => x"80",
           397 => x"bb",
           398 => x"e0",
           399 => x"90",
           400 => x"80",
           401 => x"bb",
           402 => x"a3",
           403 => x"90",
           404 => x"80",
           405 => x"bb",
           406 => x"f6",
           407 => x"90",
           408 => x"80",
           409 => x"bb",
           410 => x"86",
           411 => x"90",
           412 => x"80",
           413 => x"bb",
           414 => x"82",
           415 => x"90",
           416 => x"80",
           417 => x"bb",
           418 => x"88",
           419 => x"90",
           420 => x"80",
           421 => x"bb",
           422 => x"a8",
           423 => x"90",
           424 => x"80",
           425 => x"bb",
           426 => x"d1",
           427 => x"90",
           428 => x"80",
           429 => x"bb",
           430 => x"8a",
           431 => x"90",
           432 => x"80",
           433 => x"bb",
           434 => x"d4",
           435 => x"bb",
           436 => x"c0",
           437 => x"84",
           438 => x"80",
           439 => x"84",
           440 => x"80",
           441 => x"04",
           442 => x"0c",
           443 => x"2d",
           444 => x"08",
           445 => x"90",
           446 => x"90",
           447 => x"eb",
           448 => x"90",
           449 => x"80",
           450 => x"bb",
           451 => x"ca",
           452 => x"bb",
           453 => x"c0",
           454 => x"84",
           455 => x"82",
           456 => x"84",
           457 => x"80",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"90",
           463 => x"90",
           464 => x"a5",
           465 => x"90",
           466 => x"80",
           467 => x"bb",
           468 => x"ed",
           469 => x"bb",
           470 => x"c0",
           471 => x"84",
           472 => x"82",
           473 => x"84",
           474 => x"80",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"90",
           480 => x"90",
           481 => x"95",
           482 => x"90",
           483 => x"80",
           484 => x"bb",
           485 => x"f3",
           486 => x"bb",
           487 => x"c0",
           488 => x"84",
           489 => x"82",
           490 => x"84",
           491 => x"80",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"90",
           497 => x"90",
           498 => x"f6",
           499 => x"90",
           500 => x"80",
           501 => x"bb",
           502 => x"8c",
           503 => x"bb",
           504 => x"c0",
           505 => x"84",
           506 => x"82",
           507 => x"84",
           508 => x"80",
           509 => x"04",
           510 => x"0c",
           511 => x"2d",
           512 => x"08",
           513 => x"90",
           514 => x"90",
           515 => x"97",
           516 => x"90",
           517 => x"80",
           518 => x"bb",
           519 => x"e5",
           520 => x"bb",
           521 => x"c0",
           522 => x"84",
           523 => x"82",
           524 => x"84",
           525 => x"80",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"90",
           531 => x"90",
           532 => x"fe",
           533 => x"90",
           534 => x"80",
           535 => x"bb",
           536 => x"97",
           537 => x"bb",
           538 => x"c0",
           539 => x"84",
           540 => x"83",
           541 => x"84",
           542 => x"80",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"90",
           548 => x"90",
           549 => x"c7",
           550 => x"90",
           551 => x"80",
           552 => x"bb",
           553 => x"a5",
           554 => x"bb",
           555 => x"c0",
           556 => x"84",
           557 => x"83",
           558 => x"84",
           559 => x"80",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"90",
           565 => x"90",
           566 => x"ab",
           567 => x"90",
           568 => x"80",
           569 => x"bb",
           570 => x"f6",
           571 => x"bb",
           572 => x"c0",
           573 => x"84",
           574 => x"81",
           575 => x"84",
           576 => x"80",
           577 => x"04",
           578 => x"0c",
           579 => x"2d",
           580 => x"08",
           581 => x"90",
           582 => x"90",
           583 => x"8a",
           584 => x"90",
           585 => x"80",
           586 => x"bb",
           587 => x"d7",
           588 => x"bb",
           589 => x"c0",
           590 => x"84",
           591 => x"b1",
           592 => x"bb",
           593 => x"c0",
           594 => x"84",
           595 => x"81",
           596 => x"84",
           597 => x"80",
           598 => x"04",
           599 => x"0c",
           600 => x"2d",
           601 => x"08",
           602 => x"90",
           603 => x"90",
           604 => x"85",
           605 => x"90",
           606 => x"80",
           607 => x"bb",
           608 => x"d6",
           609 => x"bb",
           610 => x"c0",
           611 => x"3c",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"00",
           621 => x"ff",
           622 => x"06",
           623 => x"83",
           624 => x"10",
           625 => x"fc",
           626 => x"51",
           627 => x"80",
           628 => x"ff",
           629 => x"06",
           630 => x"52",
           631 => x"0a",
           632 => x"38",
           633 => x"51",
           634 => x"84",
           635 => x"f0",
           636 => x"80",
           637 => x"05",
           638 => x"0b",
           639 => x"04",
           640 => x"80",
           641 => x"00",
           642 => x"87",
           643 => x"84",
           644 => x"56",
           645 => x"84",
           646 => x"51",
           647 => x"86",
           648 => x"fa",
           649 => x"7a",
           650 => x"33",
           651 => x"06",
           652 => x"07",
           653 => x"57",
           654 => x"72",
           655 => x"06",
           656 => x"ff",
           657 => x"8a",
           658 => x"70",
           659 => x"2a",
           660 => x"56",
           661 => x"25",
           662 => x"80",
           663 => x"75",
           664 => x"3f",
           665 => x"08",
           666 => x"84",
           667 => x"ae",
           668 => x"84",
           669 => x"81",
           670 => x"ff",
           671 => x"32",
           672 => x"72",
           673 => x"51",
           674 => x"73",
           675 => x"38",
           676 => x"76",
           677 => x"bb",
           678 => x"3d",
           679 => x"0b",
           680 => x"0c",
           681 => x"04",
           682 => x"7d",
           683 => x"84",
           684 => x"34",
           685 => x"0a",
           686 => x"88",
           687 => x"52",
           688 => x"05",
           689 => x"73",
           690 => x"74",
           691 => x"0d",
           692 => x"0d",
           693 => x"05",
           694 => x"75",
           695 => x"85",
           696 => x"f1",
           697 => x"63",
           698 => x"5d",
           699 => x"1f",
           700 => x"33",
           701 => x"81",
           702 => x"55",
           703 => x"54",
           704 => x"09",
           705 => x"d2",
           706 => x"57",
           707 => x"80",
           708 => x"1c",
           709 => x"54",
           710 => x"2e",
           711 => x"d0",
           712 => x"89",
           713 => x"38",
           714 => x"70",
           715 => x"25",
           716 => x"78",
           717 => x"80",
           718 => x"7a",
           719 => x"81",
           720 => x"40",
           721 => x"2e",
           722 => x"82",
           723 => x"7b",
           724 => x"ff",
           725 => x"1d",
           726 => x"84",
           727 => x"91",
           728 => x"7a",
           729 => x"78",
           730 => x"79",
           731 => x"98",
           732 => x"2c",
           733 => x"80",
           734 => x"0a",
           735 => x"2c",
           736 => x"56",
           737 => x"24",
           738 => x"73",
           739 => x"72",
           740 => x"78",
           741 => x"58",
           742 => x"38",
           743 => x"76",
           744 => x"81",
           745 => x"81",
           746 => x"5a",
           747 => x"33",
           748 => x"fe",
           749 => x"9e",
           750 => x"76",
           751 => x"3f",
           752 => x"76",
           753 => x"ff",
           754 => x"83",
           755 => x"06",
           756 => x"8a",
           757 => x"74",
           758 => x"7e",
           759 => x"17",
           760 => x"d8",
           761 => x"72",
           762 => x"cb",
           763 => x"73",
           764 => x"e0",
           765 => x"80",
           766 => x"eb",
           767 => x"76",
           768 => x"3f",
           769 => x"58",
           770 => x"86",
           771 => x"39",
           772 => x"fe",
           773 => x"5a",
           774 => x"05",
           775 => x"83",
           776 => x"5e",
           777 => x"84",
           778 => x"79",
           779 => x"93",
           780 => x"bb",
           781 => x"ff",
           782 => x"84",
           783 => x"05",
           784 => x"89",
           785 => x"84",
           786 => x"b0",
           787 => x"7e",
           788 => x"40",
           789 => x"75",
           790 => x"3f",
           791 => x"08",
           792 => x"84",
           793 => x"7d",
           794 => x"31",
           795 => x"b2",
           796 => x"7e",
           797 => x"38",
           798 => x"80",
           799 => x"80",
           800 => x"2c",
           801 => x"86",
           802 => x"06",
           803 => x"80",
           804 => x"77",
           805 => x"29",
           806 => x"05",
           807 => x"2e",
           808 => x"84",
           809 => x"fc",
           810 => x"53",
           811 => x"58",
           812 => x"70",
           813 => x"55",
           814 => x"9e",
           815 => x"2c",
           816 => x"06",
           817 => x"73",
           818 => x"38",
           819 => x"f7",
           820 => x"2a",
           821 => x"41",
           822 => x"81",
           823 => x"80",
           824 => x"38",
           825 => x"90",
           826 => x"2c",
           827 => x"06",
           828 => x"73",
           829 => x"96",
           830 => x"2a",
           831 => x"73",
           832 => x"7a",
           833 => x"06",
           834 => x"98",
           835 => x"2a",
           836 => x"73",
           837 => x"7e",
           838 => x"73",
           839 => x"7a",
           840 => x"06",
           841 => x"2e",
           842 => x"78",
           843 => x"29",
           844 => x"05",
           845 => x"5a",
           846 => x"74",
           847 => x"7c",
           848 => x"88",
           849 => x"78",
           850 => x"29",
           851 => x"05",
           852 => x"5a",
           853 => x"80",
           854 => x"74",
           855 => x"72",
           856 => x"38",
           857 => x"80",
           858 => x"ff",
           859 => x"98",
           860 => x"55",
           861 => x"9d",
           862 => x"b0",
           863 => x"3f",
           864 => x"80",
           865 => x"ff",
           866 => x"98",
           867 => x"55",
           868 => x"e5",
           869 => x"2a",
           870 => x"5c",
           871 => x"2e",
           872 => x"76",
           873 => x"84",
           874 => x"80",
           875 => x"ca",
           876 => x"d3",
           877 => x"38",
           878 => x"94",
           879 => x"7c",
           880 => x"70",
           881 => x"87",
           882 => x"84",
           883 => x"09",
           884 => x"38",
           885 => x"5b",
           886 => x"fc",
           887 => x"78",
           888 => x"29",
           889 => x"05",
           890 => x"5a",
           891 => x"75",
           892 => x"38",
           893 => x"51",
           894 => x"e2",
           895 => x"07",
           896 => x"07",
           897 => x"5b",
           898 => x"38",
           899 => x"7a",
           900 => x"5b",
           901 => x"90",
           902 => x"05",
           903 => x"83",
           904 => x"5f",
           905 => x"5a",
           906 => x"7f",
           907 => x"77",
           908 => x"06",
           909 => x"70",
           910 => x"07",
           911 => x"80",
           912 => x"80",
           913 => x"2c",
           914 => x"56",
           915 => x"7a",
           916 => x"81",
           917 => x"7a",
           918 => x"77",
           919 => x"80",
           920 => x"80",
           921 => x"2c",
           922 => x"80",
           923 => x"b3",
           924 => x"a0",
           925 => x"3f",
           926 => x"1a",
           927 => x"ff",
           928 => x"79",
           929 => x"2e",
           930 => x"7c",
           931 => x"81",
           932 => x"51",
           933 => x"e2",
           934 => x"70",
           935 => x"06",
           936 => x"83",
           937 => x"fe",
           938 => x"52",
           939 => x"05",
           940 => x"85",
           941 => x"39",
           942 => x"06",
           943 => x"07",
           944 => x"80",
           945 => x"80",
           946 => x"2c",
           947 => x"80",
           948 => x"2a",
           949 => x"5d",
           950 => x"fd",
           951 => x"fb",
           952 => x"84",
           953 => x"70",
           954 => x"56",
           955 => x"82",
           956 => x"83",
           957 => x"5b",
           958 => x"5e",
           959 => x"7a",
           960 => x"33",
           961 => x"f8",
           962 => x"ca",
           963 => x"07",
           964 => x"33",
           965 => x"f7",
           966 => x"ba",
           967 => x"84",
           968 => x"77",
           969 => x"58",
           970 => x"82",
           971 => x"51",
           972 => x"84",
           973 => x"83",
           974 => x"78",
           975 => x"2b",
           976 => x"90",
           977 => x"87",
           978 => x"c0",
           979 => x"58",
           980 => x"be",
           981 => x"39",
           982 => x"05",
           983 => x"81",
           984 => x"41",
           985 => x"cf",
           986 => x"87",
           987 => x"bb",
           988 => x"ff",
           989 => x"71",
           990 => x"54",
           991 => x"7a",
           992 => x"7c",
           993 => x"76",
           994 => x"f7",
           995 => x"78",
           996 => x"29",
           997 => x"05",
           998 => x"5a",
           999 => x"74",
          1000 => x"38",
          1001 => x"51",
          1002 => x"e2",
          1003 => x"b0",
          1004 => x"3f",
          1005 => x"09",
          1006 => x"e3",
          1007 => x"76",
          1008 => x"3f",
          1009 => x"81",
          1010 => x"80",
          1011 => x"38",
          1012 => x"75",
          1013 => x"71",
          1014 => x"70",
          1015 => x"83",
          1016 => x"5a",
          1017 => x"fa",
          1018 => x"a2",
          1019 => x"ad",
          1020 => x"3f",
          1021 => x"54",
          1022 => x"fa",
          1023 => x"ad",
          1024 => x"75",
          1025 => x"82",
          1026 => x"81",
          1027 => x"80",
          1028 => x"38",
          1029 => x"78",
          1030 => x"2b",
          1031 => x"5a",
          1032 => x"39",
          1033 => x"51",
          1034 => x"c8",
          1035 => x"a0",
          1036 => x"3f",
          1037 => x"78",
          1038 => x"88",
          1039 => x"bb",
          1040 => x"ff",
          1041 => x"71",
          1042 => x"54",
          1043 => x"39",
          1044 => x"7e",
          1045 => x"ff",
          1046 => x"57",
          1047 => x"39",
          1048 => x"84",
          1049 => x"53",
          1050 => x"51",
          1051 => x"84",
          1052 => x"fa",
          1053 => x"55",
          1054 => x"e6",
          1055 => x"11",
          1056 => x"2a",
          1057 => x"81",
          1058 => x"58",
          1059 => x"56",
          1060 => x"09",
          1061 => x"d5",
          1062 => x"81",
          1063 => x"53",
          1064 => x"b0",
          1065 => x"e8",
          1066 => x"51",
          1067 => x"53",
          1068 => x"bb",
          1069 => x"2e",
          1070 => x"57",
          1071 => x"05",
          1072 => x"72",
          1073 => x"38",
          1074 => x"08",
          1075 => x"84",
          1076 => x"54",
          1077 => x"08",
          1078 => x"90",
          1079 => x"74",
          1080 => x"84",
          1081 => x"83",
          1082 => x"76",
          1083 => x"bb",
          1084 => x"3d",
          1085 => x"3d",
          1086 => x"56",
          1087 => x"85",
          1088 => x"81",
          1089 => x"70",
          1090 => x"55",
          1091 => x"56",
          1092 => x"09",
          1093 => x"38",
          1094 => x"05",
          1095 => x"72",
          1096 => x"81",
          1097 => x"76",
          1098 => x"bb",
          1099 => x"3d",
          1100 => x"70",
          1101 => x"33",
          1102 => x"2e",
          1103 => x"52",
          1104 => x"15",
          1105 => x"2d",
          1106 => x"08",
          1107 => x"38",
          1108 => x"81",
          1109 => x"54",
          1110 => x"38",
          1111 => x"3d",
          1112 => x"e8",
          1113 => x"51",
          1114 => x"3d",
          1115 => x"3d",
          1116 => x"85",
          1117 => x"81",
          1118 => x"81",
          1119 => x"56",
          1120 => x"72",
          1121 => x"82",
          1122 => x"54",
          1123 => x"ac",
          1124 => x"08",
          1125 => x"16",
          1126 => x"38",
          1127 => x"76",
          1128 => x"08",
          1129 => x"0c",
          1130 => x"53",
          1131 => x"16",
          1132 => x"75",
          1133 => x"0c",
          1134 => x"04",
          1135 => x"81",
          1136 => x"90",
          1137 => x"73",
          1138 => x"84",
          1139 => x"e3",
          1140 => x"08",
          1141 => x"16",
          1142 => x"d7",
          1143 => x"0d",
          1144 => x"33",
          1145 => x"06",
          1146 => x"81",
          1147 => x"56",
          1148 => x"71",
          1149 => x"86",
          1150 => x"52",
          1151 => x"72",
          1152 => x"06",
          1153 => x"2e",
          1154 => x"75",
          1155 => x"53",
          1156 => x"2e",
          1157 => x"81",
          1158 => x"8c",
          1159 => x"05",
          1160 => x"71",
          1161 => x"54",
          1162 => x"84",
          1163 => x"0d",
          1164 => x"bf",
          1165 => x"85",
          1166 => x"16",
          1167 => x"8c",
          1168 => x"16",
          1169 => x"84",
          1170 => x"0d",
          1171 => x"94",
          1172 => x"74",
          1173 => x"84",
          1174 => x"bb",
          1175 => x"25",
          1176 => x"85",
          1177 => x"90",
          1178 => x"84",
          1179 => x"ff",
          1180 => x"71",
          1181 => x"72",
          1182 => x"ff",
          1183 => x"bb",
          1184 => x"3d",
          1185 => x"a0",
          1186 => x"85",
          1187 => x"54",
          1188 => x"3d",
          1189 => x"71",
          1190 => x"71",
          1191 => x"53",
          1192 => x"f7",
          1193 => x"52",
          1194 => x"05",
          1195 => x"70",
          1196 => x"05",
          1197 => x"f0",
          1198 => x"bb",
          1199 => x"3d",
          1200 => x"3d",
          1201 => x"71",
          1202 => x"52",
          1203 => x"2e",
          1204 => x"72",
          1205 => x"70",
          1206 => x"38",
          1207 => x"05",
          1208 => x"70",
          1209 => x"34",
          1210 => x"70",
          1211 => x"84",
          1212 => x"86",
          1213 => x"70",
          1214 => x"75",
          1215 => x"70",
          1216 => x"53",
          1217 => x"13",
          1218 => x"33",
          1219 => x"11",
          1220 => x"2e",
          1221 => x"13",
          1222 => x"53",
          1223 => x"34",
          1224 => x"70",
          1225 => x"39",
          1226 => x"74",
          1227 => x"71",
          1228 => x"53",
          1229 => x"f7",
          1230 => x"70",
          1231 => x"bb",
          1232 => x"84",
          1233 => x"fd",
          1234 => x"77",
          1235 => x"54",
          1236 => x"05",
          1237 => x"70",
          1238 => x"05",
          1239 => x"f0",
          1240 => x"bb",
          1241 => x"3d",
          1242 => x"3d",
          1243 => x"71",
          1244 => x"52",
          1245 => x"2e",
          1246 => x"70",
          1247 => x"33",
          1248 => x"05",
          1249 => x"11",
          1250 => x"38",
          1251 => x"84",
          1252 => x"0d",
          1253 => x"0d",
          1254 => x"55",
          1255 => x"80",
          1256 => x"73",
          1257 => x"81",
          1258 => x"52",
          1259 => x"2e",
          1260 => x"9a",
          1261 => x"54",
          1262 => x"b7",
          1263 => x"53",
          1264 => x"80",
          1265 => x"bb",
          1266 => x"3d",
          1267 => x"80",
          1268 => x"73",
          1269 => x"51",
          1270 => x"e9",
          1271 => x"33",
          1272 => x"71",
          1273 => x"38",
          1274 => x"84",
          1275 => x"86",
          1276 => x"71",
          1277 => x"0c",
          1278 => x"04",
          1279 => x"77",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"08",
          1284 => x"55",
          1285 => x"3f",
          1286 => x"08",
          1287 => x"84",
          1288 => x"9b",
          1289 => x"84",
          1290 => x"80",
          1291 => x"53",
          1292 => x"bb",
          1293 => x"fe",
          1294 => x"bb",
          1295 => x"73",
          1296 => x"0c",
          1297 => x"04",
          1298 => x"75",
          1299 => x"54",
          1300 => x"71",
          1301 => x"38",
          1302 => x"05",
          1303 => x"70",
          1304 => x"38",
          1305 => x"71",
          1306 => x"81",
          1307 => x"ff",
          1308 => x"31",
          1309 => x"84",
          1310 => x"85",
          1311 => x"fd",
          1312 => x"77",
          1313 => x"53",
          1314 => x"80",
          1315 => x"72",
          1316 => x"05",
          1317 => x"11",
          1318 => x"38",
          1319 => x"84",
          1320 => x"0d",
          1321 => x"0d",
          1322 => x"54",
          1323 => x"80",
          1324 => x"76",
          1325 => x"3f",
          1326 => x"08",
          1327 => x"53",
          1328 => x"8d",
          1329 => x"80",
          1330 => x"84",
          1331 => x"31",
          1332 => x"72",
          1333 => x"cb",
          1334 => x"72",
          1335 => x"c3",
          1336 => x"74",
          1337 => x"72",
          1338 => x"2b",
          1339 => x"55",
          1340 => x"76",
          1341 => x"72",
          1342 => x"2a",
          1343 => x"77",
          1344 => x"31",
          1345 => x"2c",
          1346 => x"7b",
          1347 => x"71",
          1348 => x"5c",
          1349 => x"55",
          1350 => x"74",
          1351 => x"10",
          1352 => x"71",
          1353 => x"0c",
          1354 => x"04",
          1355 => x"76",
          1356 => x"80",
          1357 => x"70",
          1358 => x"25",
          1359 => x"90",
          1360 => x"71",
          1361 => x"fe",
          1362 => x"30",
          1363 => x"83",
          1364 => x"31",
          1365 => x"70",
          1366 => x"70",
          1367 => x"25",
          1368 => x"71",
          1369 => x"2a",
          1370 => x"1b",
          1371 => x"06",
          1372 => x"80",
          1373 => x"71",
          1374 => x"2a",
          1375 => x"81",
          1376 => x"06",
          1377 => x"74",
          1378 => x"19",
          1379 => x"84",
          1380 => x"54",
          1381 => x"56",
          1382 => x"55",
          1383 => x"56",
          1384 => x"58",
          1385 => x"86",
          1386 => x"fd",
          1387 => x"77",
          1388 => x"53",
          1389 => x"94",
          1390 => x"84",
          1391 => x"74",
          1392 => x"bb",
          1393 => x"85",
          1394 => x"fa",
          1395 => x"7a",
          1396 => x"53",
          1397 => x"8b",
          1398 => x"fe",
          1399 => x"bb",
          1400 => x"e0",
          1401 => x"80",
          1402 => x"73",
          1403 => x"3f",
          1404 => x"84",
          1405 => x"73",
          1406 => x"26",
          1407 => x"80",
          1408 => x"2e",
          1409 => x"12",
          1410 => x"a0",
          1411 => x"71",
          1412 => x"54",
          1413 => x"74",
          1414 => x"38",
          1415 => x"9f",
          1416 => x"10",
          1417 => x"72",
          1418 => x"9f",
          1419 => x"06",
          1420 => x"75",
          1421 => x"1c",
          1422 => x"52",
          1423 => x"53",
          1424 => x"72",
          1425 => x"0c",
          1426 => x"04",
          1427 => x"78",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"9f",
          1431 => x"73",
          1432 => x"74",
          1433 => x"75",
          1434 => x"56",
          1435 => x"fc",
          1436 => x"bb",
          1437 => x"32",
          1438 => x"bb",
          1439 => x"3d",
          1440 => x"3d",
          1441 => x"5b",
          1442 => x"7b",
          1443 => x"70",
          1444 => x"59",
          1445 => x"09",
          1446 => x"38",
          1447 => x"78",
          1448 => x"55",
          1449 => x"2e",
          1450 => x"ad",
          1451 => x"38",
          1452 => x"81",
          1453 => x"14",
          1454 => x"77",
          1455 => x"db",
          1456 => x"80",
          1457 => x"27",
          1458 => x"80",
          1459 => x"89",
          1460 => x"70",
          1461 => x"55",
          1462 => x"70",
          1463 => x"51",
          1464 => x"27",
          1465 => x"13",
          1466 => x"06",
          1467 => x"73",
          1468 => x"38",
          1469 => x"81",
          1470 => x"76",
          1471 => x"16",
          1472 => x"70",
          1473 => x"56",
          1474 => x"ff",
          1475 => x"80",
          1476 => x"75",
          1477 => x"7a",
          1478 => x"75",
          1479 => x"0c",
          1480 => x"04",
          1481 => x"70",
          1482 => x"33",
          1483 => x"73",
          1484 => x"81",
          1485 => x"38",
          1486 => x"78",
          1487 => x"55",
          1488 => x"e2",
          1489 => x"90",
          1490 => x"f8",
          1491 => x"81",
          1492 => x"27",
          1493 => x"14",
          1494 => x"88",
          1495 => x"27",
          1496 => x"75",
          1497 => x"0c",
          1498 => x"04",
          1499 => x"15",
          1500 => x"70",
          1501 => x"80",
          1502 => x"39",
          1503 => x"bb",
          1504 => x"3d",
          1505 => x"3d",
          1506 => x"5b",
          1507 => x"7b",
          1508 => x"70",
          1509 => x"59",
          1510 => x"09",
          1511 => x"38",
          1512 => x"78",
          1513 => x"55",
          1514 => x"2e",
          1515 => x"ad",
          1516 => x"38",
          1517 => x"81",
          1518 => x"14",
          1519 => x"77",
          1520 => x"db",
          1521 => x"80",
          1522 => x"27",
          1523 => x"80",
          1524 => x"89",
          1525 => x"70",
          1526 => x"55",
          1527 => x"70",
          1528 => x"51",
          1529 => x"27",
          1530 => x"13",
          1531 => x"06",
          1532 => x"73",
          1533 => x"38",
          1534 => x"81",
          1535 => x"76",
          1536 => x"16",
          1537 => x"70",
          1538 => x"56",
          1539 => x"ff",
          1540 => x"80",
          1541 => x"75",
          1542 => x"7a",
          1543 => x"75",
          1544 => x"0c",
          1545 => x"04",
          1546 => x"70",
          1547 => x"33",
          1548 => x"73",
          1549 => x"81",
          1550 => x"38",
          1551 => x"78",
          1552 => x"55",
          1553 => x"e2",
          1554 => x"90",
          1555 => x"f8",
          1556 => x"81",
          1557 => x"27",
          1558 => x"14",
          1559 => x"88",
          1560 => x"27",
          1561 => x"75",
          1562 => x"0c",
          1563 => x"04",
          1564 => x"15",
          1565 => x"70",
          1566 => x"80",
          1567 => x"39",
          1568 => x"bb",
          1569 => x"3d",
          1570 => x"d8",
          1571 => x"bb",
          1572 => x"ff",
          1573 => x"84",
          1574 => x"3d",
          1575 => x"71",
          1576 => x"38",
          1577 => x"83",
          1578 => x"52",
          1579 => x"83",
          1580 => x"ef",
          1581 => x"3d",
          1582 => x"cf",
          1583 => x"b3",
          1584 => x"0d",
          1585 => x"d4",
          1586 => x"3f",
          1587 => x"04",
          1588 => x"51",
          1589 => x"83",
          1590 => x"83",
          1591 => x"ef",
          1592 => x"3d",
          1593 => x"d0",
          1594 => x"87",
          1595 => x"0d",
          1596 => x"b4",
          1597 => x"3f",
          1598 => x"04",
          1599 => x"51",
          1600 => x"83",
          1601 => x"83",
          1602 => x"ee",
          1603 => x"3d",
          1604 => x"d1",
          1605 => x"db",
          1606 => x"0d",
          1607 => x"9c",
          1608 => x"3f",
          1609 => x"04",
          1610 => x"51",
          1611 => x"83",
          1612 => x"83",
          1613 => x"ee",
          1614 => x"3d",
          1615 => x"d1",
          1616 => x"af",
          1617 => x"0d",
          1618 => x"f4",
          1619 => x"3f",
          1620 => x"04",
          1621 => x"51",
          1622 => x"83",
          1623 => x"83",
          1624 => x"ee",
          1625 => x"3d",
          1626 => x"d2",
          1627 => x"83",
          1628 => x"0d",
          1629 => x"b8",
          1630 => x"3f",
          1631 => x"04",
          1632 => x"51",
          1633 => x"83",
          1634 => x"83",
          1635 => x"ed",
          1636 => x"3d",
          1637 => x"ec",
          1638 => x"97",
          1639 => x"84",
          1640 => x"05",
          1641 => x"80",
          1642 => x"3d",
          1643 => x"70",
          1644 => x"25",
          1645 => x"59",
          1646 => x"87",
          1647 => x"38",
          1648 => x"77",
          1649 => x"ff",
          1650 => x"93",
          1651 => x"e2",
          1652 => x"77",
          1653 => x"70",
          1654 => x"97",
          1655 => x"bb",
          1656 => x"84",
          1657 => x"80",
          1658 => x"38",
          1659 => x"af",
          1660 => x"30",
          1661 => x"80",
          1662 => x"70",
          1663 => x"06",
          1664 => x"58",
          1665 => x"aa",
          1666 => x"98",
          1667 => x"74",
          1668 => x"80",
          1669 => x"52",
          1670 => x"29",
          1671 => x"3f",
          1672 => x"08",
          1673 => x"84",
          1674 => x"83",
          1675 => x"df",
          1676 => x"84",
          1677 => x"81",
          1678 => x"04",
          1679 => x"08",
          1680 => x"88",
          1681 => x"84",
          1682 => x"96",
          1683 => x"05",
          1684 => x"53",
          1685 => x"51",
          1686 => x"3f",
          1687 => x"08",
          1688 => x"84",
          1689 => x"38",
          1690 => x"80",
          1691 => x"38",
          1692 => x"17",
          1693 => x"39",
          1694 => x"74",
          1695 => x"3f",
          1696 => x"08",
          1697 => x"f4",
          1698 => x"bb",
          1699 => x"83",
          1700 => x"78",
          1701 => x"e0",
          1702 => x"3f",
          1703 => x"f8",
          1704 => x"02",
          1705 => x"05",
          1706 => x"ff",
          1707 => x"7b",
          1708 => x"fd",
          1709 => x"bb",
          1710 => x"38",
          1711 => x"91",
          1712 => x"2e",
          1713 => x"84",
          1714 => x"8a",
          1715 => x"78",
          1716 => x"e4",
          1717 => x"60",
          1718 => x"84",
          1719 => x"7e",
          1720 => x"84",
          1721 => x"84",
          1722 => x"8a",
          1723 => x"f3",
          1724 => x"61",
          1725 => x"05",
          1726 => x"33",
          1727 => x"68",
          1728 => x"5c",
          1729 => x"78",
          1730 => x"82",
          1731 => x"83",
          1732 => x"dd",
          1733 => x"d3",
          1734 => x"ec",
          1735 => x"73",
          1736 => x"38",
          1737 => x"81",
          1738 => x"a0",
          1739 => x"38",
          1740 => x"72",
          1741 => x"a7",
          1742 => x"52",
          1743 => x"51",
          1744 => x"81",
          1745 => x"e8",
          1746 => x"a0",
          1747 => x"3f",
          1748 => x"dc",
          1749 => x"a0",
          1750 => x"3f",
          1751 => x"79",
          1752 => x"38",
          1753 => x"33",
          1754 => x"55",
          1755 => x"83",
          1756 => x"80",
          1757 => x"27",
          1758 => x"53",
          1759 => x"70",
          1760 => x"56",
          1761 => x"2e",
          1762 => x"fe",
          1763 => x"ee",
          1764 => x"e8",
          1765 => x"51",
          1766 => x"81",
          1767 => x"76",
          1768 => x"83",
          1769 => x"e9",
          1770 => x"18",
          1771 => x"58",
          1772 => x"c8",
          1773 => x"84",
          1774 => x"70",
          1775 => x"54",
          1776 => x"81",
          1777 => x"9b",
          1778 => x"38",
          1779 => x"76",
          1780 => x"b9",
          1781 => x"84",
          1782 => x"8f",
          1783 => x"83",
          1784 => x"dc",
          1785 => x"14",
          1786 => x"08",
          1787 => x"51",
          1788 => x"78",
          1789 => x"b8",
          1790 => x"39",
          1791 => x"51",
          1792 => x"82",
          1793 => x"e8",
          1794 => x"a0",
          1795 => x"3f",
          1796 => x"fe",
          1797 => x"18",
          1798 => x"27",
          1799 => x"22",
          1800 => x"ac",
          1801 => x"3f",
          1802 => x"e6",
          1803 => x"54",
          1804 => x"ba",
          1805 => x"26",
          1806 => x"99",
          1807 => x"b4",
          1808 => x"3f",
          1809 => x"e6",
          1810 => x"54",
          1811 => x"9e",
          1812 => x"27",
          1813 => x"73",
          1814 => x"7a",
          1815 => x"72",
          1816 => x"d3",
          1817 => x"a0",
          1818 => x"84",
          1819 => x"53",
          1820 => x"e9",
          1821 => x"74",
          1822 => x"fd",
          1823 => x"e6",
          1824 => x"73",
          1825 => x"3f",
          1826 => x"fe",
          1827 => x"d0",
          1828 => x"bb",
          1829 => x"ff",
          1830 => x"59",
          1831 => x"fc",
          1832 => x"59",
          1833 => x"2e",
          1834 => x"fc",
          1835 => x"59",
          1836 => x"80",
          1837 => x"3f",
          1838 => x"08",
          1839 => x"98",
          1840 => x"32",
          1841 => x"9b",
          1842 => x"70",
          1843 => x"75",
          1844 => x"55",
          1845 => x"58",
          1846 => x"25",
          1847 => x"80",
          1848 => x"3f",
          1849 => x"08",
          1850 => x"98",
          1851 => x"32",
          1852 => x"9b",
          1853 => x"70",
          1854 => x"75",
          1855 => x"55",
          1856 => x"58",
          1857 => x"24",
          1858 => x"fd",
          1859 => x"0b",
          1860 => x"0c",
          1861 => x"04",
          1862 => x"87",
          1863 => x"08",
          1864 => x"3f",
          1865 => x"8d",
          1866 => x"d0",
          1867 => x"3f",
          1868 => x"81",
          1869 => x"2a",
          1870 => x"51",
          1871 => x"b7",
          1872 => x"2a",
          1873 => x"51",
          1874 => x"89",
          1875 => x"2a",
          1876 => x"51",
          1877 => x"db",
          1878 => x"2a",
          1879 => x"51",
          1880 => x"ad",
          1881 => x"2a",
          1882 => x"51",
          1883 => x"ff",
          1884 => x"2a",
          1885 => x"51",
          1886 => x"d2",
          1887 => x"2a",
          1888 => x"51",
          1889 => x"38",
          1890 => x"81",
          1891 => x"88",
          1892 => x"3f",
          1893 => x"04",
          1894 => x"99",
          1895 => x"e8",
          1896 => x"3f",
          1897 => x"8d",
          1898 => x"3f",
          1899 => x"04",
          1900 => x"81",
          1901 => x"fc",
          1902 => x"3f",
          1903 => x"f5",
          1904 => x"2a",
          1905 => x"72",
          1906 => x"38",
          1907 => x"51",
          1908 => x"83",
          1909 => x"9b",
          1910 => x"51",
          1911 => x"72",
          1912 => x"81",
          1913 => x"71",
          1914 => x"9c",
          1915 => x"81",
          1916 => x"3f",
          1917 => x"51",
          1918 => x"80",
          1919 => x"3f",
          1920 => x"70",
          1921 => x"52",
          1922 => x"fe",
          1923 => x"be",
          1924 => x"9b",
          1925 => x"d5",
          1926 => x"b1",
          1927 => x"9b",
          1928 => x"85",
          1929 => x"06",
          1930 => x"80",
          1931 => x"38",
          1932 => x"81",
          1933 => x"3f",
          1934 => x"51",
          1935 => x"80",
          1936 => x"3f",
          1937 => x"70",
          1938 => x"52",
          1939 => x"fe",
          1940 => x"bd",
          1941 => x"9a",
          1942 => x"d5",
          1943 => x"ed",
          1944 => x"9a",
          1945 => x"83",
          1946 => x"06",
          1947 => x"80",
          1948 => x"38",
          1949 => x"81",
          1950 => x"3f",
          1951 => x"51",
          1952 => x"80",
          1953 => x"3f",
          1954 => x"70",
          1955 => x"52",
          1956 => x"fd",
          1957 => x"bd",
          1958 => x"0d",
          1959 => x"41",
          1960 => x"de",
          1961 => x"81",
          1962 => x"81",
          1963 => x"84",
          1964 => x"81",
          1965 => x"3d",
          1966 => x"61",
          1967 => x"38",
          1968 => x"51",
          1969 => x"98",
          1970 => x"d6",
          1971 => x"b8",
          1972 => x"80",
          1973 => x"52",
          1974 => x"a3",
          1975 => x"83",
          1976 => x"70",
          1977 => x"5b",
          1978 => x"2e",
          1979 => x"79",
          1980 => x"88",
          1981 => x"ff",
          1982 => x"82",
          1983 => x"38",
          1984 => x"5a",
          1985 => x"83",
          1986 => x"33",
          1987 => x"2e",
          1988 => x"8c",
          1989 => x"70",
          1990 => x"7b",
          1991 => x"38",
          1992 => x"9b",
          1993 => x"7b",
          1994 => x"ef",
          1995 => x"08",
          1996 => x"f4",
          1997 => x"84",
          1998 => x"84",
          1999 => x"53",
          2000 => x"5d",
          2001 => x"84",
          2002 => x"8b",
          2003 => x"33",
          2004 => x"2e",
          2005 => x"81",
          2006 => x"ff",
          2007 => x"9b",
          2008 => x"38",
          2009 => x"5c",
          2010 => x"fe",
          2011 => x"f8",
          2012 => x"e9",
          2013 => x"bb",
          2014 => x"84",
          2015 => x"80",
          2016 => x"38",
          2017 => x"08",
          2018 => x"ff",
          2019 => x"91",
          2020 => x"bb",
          2021 => x"62",
          2022 => x"7a",
          2023 => x"84",
          2024 => x"84",
          2025 => x"80",
          2026 => x"84",
          2027 => x"80",
          2028 => x"0b",
          2029 => x"5b",
          2030 => x"8d",
          2031 => x"82",
          2032 => x"38",
          2033 => x"82",
          2034 => x"54",
          2035 => x"d7",
          2036 => x"51",
          2037 => x"83",
          2038 => x"84",
          2039 => x"7d",
          2040 => x"80",
          2041 => x"0a",
          2042 => x"0a",
          2043 => x"f5",
          2044 => x"bb",
          2045 => x"bb",
          2046 => x"70",
          2047 => x"07",
          2048 => x"5b",
          2049 => x"5a",
          2050 => x"83",
          2051 => x"78",
          2052 => x"78",
          2053 => x"38",
          2054 => x"81",
          2055 => x"5a",
          2056 => x"38",
          2057 => x"61",
          2058 => x"5d",
          2059 => x"38",
          2060 => x"81",
          2061 => x"51",
          2062 => x"3f",
          2063 => x"51",
          2064 => x"7e",
          2065 => x"53",
          2066 => x"51",
          2067 => x"0b",
          2068 => x"f8",
          2069 => x"ff",
          2070 => x"79",
          2071 => x"81",
          2072 => x"a8",
          2073 => x"94",
          2074 => x"8a",
          2075 => x"84",
          2076 => x"38",
          2077 => x"0b",
          2078 => x"34",
          2079 => x"53",
          2080 => x"7e",
          2081 => x"cc",
          2082 => x"84",
          2083 => x"a0",
          2084 => x"84",
          2085 => x"db",
          2086 => x"83",
          2087 => x"70",
          2088 => x"5f",
          2089 => x"2e",
          2090 => x"fc",
          2091 => x"39",
          2092 => x"51",
          2093 => x"3f",
          2094 => x"0b",
          2095 => x"34",
          2096 => x"d6",
          2097 => x"53",
          2098 => x"7e",
          2099 => x"3f",
          2100 => x"5a",
          2101 => x"38",
          2102 => x"1a",
          2103 => x"1b",
          2104 => x"81",
          2105 => x"fc",
          2106 => x"10",
          2107 => x"05",
          2108 => x"04",
          2109 => x"d7",
          2110 => x"51",
          2111 => x"60",
          2112 => x"84",
          2113 => x"82",
          2114 => x"84",
          2115 => x"61",
          2116 => x"06",
          2117 => x"81",
          2118 => x"45",
          2119 => x"aa",
          2120 => x"8c",
          2121 => x"3f",
          2122 => x"94",
          2123 => x"8c",
          2124 => x"9c",
          2125 => x"83",
          2126 => x"80",
          2127 => x"a4",
          2128 => x"d2",
          2129 => x"8f",
          2130 => x"e4",
          2131 => x"39",
          2132 => x"fa",
          2133 => x"52",
          2134 => x"c0",
          2135 => x"ea",
          2136 => x"8e",
          2137 => x"39",
          2138 => x"51",
          2139 => x"80",
          2140 => x"83",
          2141 => x"dd",
          2142 => x"ed",
          2143 => x"39",
          2144 => x"84",
          2145 => x"80",
          2146 => x"fa",
          2147 => x"84",
          2148 => x"fa",
          2149 => x"52",
          2150 => x"51",
          2151 => x"68",
          2152 => x"84",
          2153 => x"80",
          2154 => x"38",
          2155 => x"08",
          2156 => x"80",
          2157 => x"3f",
          2158 => x"b8",
          2159 => x"11",
          2160 => x"05",
          2161 => x"3f",
          2162 => x"08",
          2163 => x"fa",
          2164 => x"83",
          2165 => x"d0",
          2166 => x"59",
          2167 => x"3d",
          2168 => x"53",
          2169 => x"51",
          2170 => x"84",
          2171 => x"80",
          2172 => x"38",
          2173 => x"f0",
          2174 => x"80",
          2175 => x"82",
          2176 => x"84",
          2177 => x"38",
          2178 => x"08",
          2179 => x"83",
          2180 => x"cf",
          2181 => x"e6",
          2182 => x"80",
          2183 => x"51",
          2184 => x"7e",
          2185 => x"59",
          2186 => x"f9",
          2187 => x"9f",
          2188 => x"38",
          2189 => x"70",
          2190 => x"39",
          2191 => x"f4",
          2192 => x"80",
          2193 => x"ba",
          2194 => x"84",
          2195 => x"f8",
          2196 => x"3d",
          2197 => x"53",
          2198 => x"51",
          2199 => x"84",
          2200 => x"86",
          2201 => x"59",
          2202 => x"78",
          2203 => x"c8",
          2204 => x"3f",
          2205 => x"08",
          2206 => x"52",
          2207 => x"a3",
          2208 => x"7e",
          2209 => x"ae",
          2210 => x"38",
          2211 => x"87",
          2212 => x"82",
          2213 => x"59",
          2214 => x"3d",
          2215 => x"53",
          2216 => x"51",
          2217 => x"84",
          2218 => x"80",
          2219 => x"38",
          2220 => x"fc",
          2221 => x"80",
          2222 => x"ca",
          2223 => x"84",
          2224 => x"f8",
          2225 => x"3d",
          2226 => x"53",
          2227 => x"51",
          2228 => x"84",
          2229 => x"80",
          2230 => x"38",
          2231 => x"51",
          2232 => x"68",
          2233 => x"78",
          2234 => x"8d",
          2235 => x"33",
          2236 => x"5c",
          2237 => x"2e",
          2238 => x"55",
          2239 => x"33",
          2240 => x"83",
          2241 => x"cd",
          2242 => x"66",
          2243 => x"19",
          2244 => x"59",
          2245 => x"3d",
          2246 => x"53",
          2247 => x"51",
          2248 => x"84",
          2249 => x"80",
          2250 => x"38",
          2251 => x"fc",
          2252 => x"80",
          2253 => x"ce",
          2254 => x"84",
          2255 => x"f7",
          2256 => x"3d",
          2257 => x"53",
          2258 => x"51",
          2259 => x"84",
          2260 => x"80",
          2261 => x"38",
          2262 => x"51",
          2263 => x"68",
          2264 => x"27",
          2265 => x"65",
          2266 => x"81",
          2267 => x"7c",
          2268 => x"05",
          2269 => x"b8",
          2270 => x"11",
          2271 => x"05",
          2272 => x"3f",
          2273 => x"08",
          2274 => x"be",
          2275 => x"fe",
          2276 => x"ff",
          2277 => x"e7",
          2278 => x"bb",
          2279 => x"38",
          2280 => x"54",
          2281 => x"8c",
          2282 => x"3f",
          2283 => x"08",
          2284 => x"52",
          2285 => x"eb",
          2286 => x"7e",
          2287 => x"ae",
          2288 => x"38",
          2289 => x"84",
          2290 => x"81",
          2291 => x"39",
          2292 => x"80",
          2293 => x"79",
          2294 => x"05",
          2295 => x"fe",
          2296 => x"ff",
          2297 => x"e7",
          2298 => x"bb",
          2299 => x"2e",
          2300 => x"68",
          2301 => x"db",
          2302 => x"34",
          2303 => x"49",
          2304 => x"fc",
          2305 => x"80",
          2306 => x"fa",
          2307 => x"84",
          2308 => x"38",
          2309 => x"b8",
          2310 => x"11",
          2311 => x"05",
          2312 => x"3f",
          2313 => x"08",
          2314 => x"9e",
          2315 => x"fe",
          2316 => x"ff",
          2317 => x"e6",
          2318 => x"bb",
          2319 => x"2e",
          2320 => x"b8",
          2321 => x"11",
          2322 => x"05",
          2323 => x"3f",
          2324 => x"08",
          2325 => x"bb",
          2326 => x"83",
          2327 => x"cb",
          2328 => x"67",
          2329 => x"7a",
          2330 => x"65",
          2331 => x"70",
          2332 => x"0c",
          2333 => x"f5",
          2334 => x"d9",
          2335 => x"ca",
          2336 => x"ff",
          2337 => x"87",
          2338 => x"bb",
          2339 => x"3d",
          2340 => x"52",
          2341 => x"3f",
          2342 => x"bb",
          2343 => x"78",
          2344 => x"3f",
          2345 => x"08",
          2346 => x"9e",
          2347 => x"84",
          2348 => x"e6",
          2349 => x"39",
          2350 => x"84",
          2351 => x"80",
          2352 => x"c2",
          2353 => x"84",
          2354 => x"83",
          2355 => x"5a",
          2356 => x"83",
          2357 => x"f3",
          2358 => x"b8",
          2359 => x"11",
          2360 => x"05",
          2361 => x"3f",
          2362 => x"08",
          2363 => x"f4",
          2364 => x"79",
          2365 => x"8a",
          2366 => x"c4",
          2367 => x"3d",
          2368 => x"53",
          2369 => x"51",
          2370 => x"84",
          2371 => x"80",
          2372 => x"80",
          2373 => x"7a",
          2374 => x"38",
          2375 => x"90",
          2376 => x"70",
          2377 => x"2a",
          2378 => x"5f",
          2379 => x"2e",
          2380 => x"a0",
          2381 => x"88",
          2382 => x"a8",
          2383 => x"3f",
          2384 => x"54",
          2385 => x"52",
          2386 => x"a3",
          2387 => x"b4",
          2388 => x"3f",
          2389 => x"64",
          2390 => x"59",
          2391 => x"45",
          2392 => x"f0",
          2393 => x"80",
          2394 => x"96",
          2395 => x"84",
          2396 => x"f2",
          2397 => x"64",
          2398 => x"64",
          2399 => x"b8",
          2400 => x"11",
          2401 => x"05",
          2402 => x"3f",
          2403 => x"08",
          2404 => x"b6",
          2405 => x"02",
          2406 => x"22",
          2407 => x"05",
          2408 => x"45",
          2409 => x"f0",
          2410 => x"80",
          2411 => x"d2",
          2412 => x"84",
          2413 => x"f2",
          2414 => x"5e",
          2415 => x"05",
          2416 => x"82",
          2417 => x"7d",
          2418 => x"fe",
          2419 => x"ff",
          2420 => x"e1",
          2421 => x"bb",
          2422 => x"b9",
          2423 => x"39",
          2424 => x"fc",
          2425 => x"80",
          2426 => x"9a",
          2427 => x"84",
          2428 => x"81",
          2429 => x"5c",
          2430 => x"05",
          2431 => x"68",
          2432 => x"fb",
          2433 => x"3d",
          2434 => x"53",
          2435 => x"51",
          2436 => x"84",
          2437 => x"80",
          2438 => x"38",
          2439 => x"0c",
          2440 => x"05",
          2441 => x"f7",
          2442 => x"83",
          2443 => x"06",
          2444 => x"7b",
          2445 => x"a0",
          2446 => x"83",
          2447 => x"7c",
          2448 => x"3f",
          2449 => x"7b",
          2450 => x"d9",
          2451 => x"87",
          2452 => x"cc",
          2453 => x"3f",
          2454 => x"b8",
          2455 => x"11",
          2456 => x"05",
          2457 => x"3f",
          2458 => x"08",
          2459 => x"38",
          2460 => x"80",
          2461 => x"79",
          2462 => x"5b",
          2463 => x"f7",
          2464 => x"f4",
          2465 => x"7b",
          2466 => x"cf",
          2467 => x"cc",
          2468 => x"ea",
          2469 => x"89",
          2470 => x"80",
          2471 => x"83",
          2472 => x"49",
          2473 => x"83",
          2474 => x"d3",
          2475 => x"59",
          2476 => x"83",
          2477 => x"d3",
          2478 => x"59",
          2479 => x"83",
          2480 => x"59",
          2481 => x"a5",
          2482 => x"d0",
          2483 => x"8b",
          2484 => x"f8",
          2485 => x"3f",
          2486 => x"83",
          2487 => x"59",
          2488 => x"9b",
          2489 => x"d4",
          2490 => x"92",
          2491 => x"8b",
          2492 => x"80",
          2493 => x"83",
          2494 => x"49",
          2495 => x"83",
          2496 => x"5e",
          2497 => x"9b",
          2498 => x"dc",
          2499 => x"ee",
          2500 => x"86",
          2501 => x"80",
          2502 => x"83",
          2503 => x"49",
          2504 => x"83",
          2505 => x"5d",
          2506 => x"94",
          2507 => x"e4",
          2508 => x"ca",
          2509 => x"f0",
          2510 => x"05",
          2511 => x"39",
          2512 => x"08",
          2513 => x"fb",
          2514 => x"3d",
          2515 => x"84",
          2516 => x"87",
          2517 => x"70",
          2518 => x"87",
          2519 => x"74",
          2520 => x"3f",
          2521 => x"08",
          2522 => x"08",
          2523 => x"84",
          2524 => x"51",
          2525 => x"74",
          2526 => x"08",
          2527 => x"87",
          2528 => x"70",
          2529 => x"87",
          2530 => x"74",
          2531 => x"3f",
          2532 => x"08",
          2533 => x"08",
          2534 => x"84",
          2535 => x"51",
          2536 => x"74",
          2537 => x"08",
          2538 => x"8c",
          2539 => x"87",
          2540 => x"0c",
          2541 => x"0b",
          2542 => x"94",
          2543 => x"ba",
          2544 => x"b9",
          2545 => x"84",
          2546 => x"34",
          2547 => x"e6",
          2548 => x"3d",
          2549 => x"0c",
          2550 => x"84",
          2551 => x"56",
          2552 => x"89",
          2553 => x"98",
          2554 => x"51",
          2555 => x"83",
          2556 => x"83",
          2557 => x"c4",
          2558 => x"f3",
          2559 => x"52",
          2560 => x"3f",
          2561 => x"54",
          2562 => x"53",
          2563 => x"52",
          2564 => x"51",
          2565 => x"8d",
          2566 => x"d3",
          2567 => x"d3",
          2568 => x"83",
          2569 => x"c3",
          2570 => x"80",
          2571 => x"d4",
          2572 => x"d4",
          2573 => x"3f",
          2574 => x"3d",
          2575 => x"08",
          2576 => x"75",
          2577 => x"73",
          2578 => x"38",
          2579 => x"81",
          2580 => x"52",
          2581 => x"09",
          2582 => x"38",
          2583 => x"33",
          2584 => x"06",
          2585 => x"70",
          2586 => x"38",
          2587 => x"06",
          2588 => x"2e",
          2589 => x"74",
          2590 => x"2e",
          2591 => x"80",
          2592 => x"81",
          2593 => x"54",
          2594 => x"2e",
          2595 => x"54",
          2596 => x"8b",
          2597 => x"2e",
          2598 => x"12",
          2599 => x"80",
          2600 => x"06",
          2601 => x"a0",
          2602 => x"06",
          2603 => x"54",
          2604 => x"70",
          2605 => x"25",
          2606 => x"52",
          2607 => x"2e",
          2608 => x"72",
          2609 => x"54",
          2610 => x"0c",
          2611 => x"84",
          2612 => x"87",
          2613 => x"70",
          2614 => x"38",
          2615 => x"ff",
          2616 => x"12",
          2617 => x"33",
          2618 => x"06",
          2619 => x"70",
          2620 => x"38",
          2621 => x"39",
          2622 => x"81",
          2623 => x"72",
          2624 => x"81",
          2625 => x"38",
          2626 => x"3d",
          2627 => x"72",
          2628 => x"80",
          2629 => x"84",
          2630 => x"0d",
          2631 => x"fc",
          2632 => x"51",
          2633 => x"84",
          2634 => x"80",
          2635 => x"74",
          2636 => x"0c",
          2637 => x"04",
          2638 => x"76",
          2639 => x"ff",
          2640 => x"81",
          2641 => x"26",
          2642 => x"83",
          2643 => x"05",
          2644 => x"73",
          2645 => x"8a",
          2646 => x"33",
          2647 => x"70",
          2648 => x"fe",
          2649 => x"33",
          2650 => x"73",
          2651 => x"f2",
          2652 => x"33",
          2653 => x"74",
          2654 => x"e6",
          2655 => x"22",
          2656 => x"74",
          2657 => x"80",
          2658 => x"13",
          2659 => x"52",
          2660 => x"26",
          2661 => x"81",
          2662 => x"98",
          2663 => x"22",
          2664 => x"bc",
          2665 => x"33",
          2666 => x"b8",
          2667 => x"33",
          2668 => x"b4",
          2669 => x"33",
          2670 => x"b0",
          2671 => x"33",
          2672 => x"ac",
          2673 => x"33",
          2674 => x"a8",
          2675 => x"c0",
          2676 => x"73",
          2677 => x"a0",
          2678 => x"87",
          2679 => x"0c",
          2680 => x"84",
          2681 => x"86",
          2682 => x"f3",
          2683 => x"5b",
          2684 => x"9c",
          2685 => x"0c",
          2686 => x"bc",
          2687 => x"7b",
          2688 => x"98",
          2689 => x"7b",
          2690 => x"87",
          2691 => x"08",
          2692 => x"1c",
          2693 => x"98",
          2694 => x"7b",
          2695 => x"87",
          2696 => x"08",
          2697 => x"1c",
          2698 => x"98",
          2699 => x"7b",
          2700 => x"87",
          2701 => x"08",
          2702 => x"1c",
          2703 => x"98",
          2704 => x"79",
          2705 => x"80",
          2706 => x"83",
          2707 => x"59",
          2708 => x"ff",
          2709 => x"1b",
          2710 => x"1b",
          2711 => x"1b",
          2712 => x"1b",
          2713 => x"1b",
          2714 => x"83",
          2715 => x"52",
          2716 => x"51",
          2717 => x"3f",
          2718 => x"04",
          2719 => x"02",
          2720 => x"53",
          2721 => x"a8",
          2722 => x"80",
          2723 => x"84",
          2724 => x"98",
          2725 => x"2c",
          2726 => x"ff",
          2727 => x"06",
          2728 => x"83",
          2729 => x"71",
          2730 => x"0c",
          2731 => x"04",
          2732 => x"e9",
          2733 => x"bb",
          2734 => x"2b",
          2735 => x"51",
          2736 => x"2e",
          2737 => x"df",
          2738 => x"80",
          2739 => x"84",
          2740 => x"98",
          2741 => x"2c",
          2742 => x"ff",
          2743 => x"c7",
          2744 => x"0d",
          2745 => x"52",
          2746 => x"54",
          2747 => x"e8",
          2748 => x"bb",
          2749 => x"2b",
          2750 => x"51",
          2751 => x"2e",
          2752 => x"72",
          2753 => x"54",
          2754 => x"25",
          2755 => x"84",
          2756 => x"85",
          2757 => x"fc",
          2758 => x"9b",
          2759 => x"f3",
          2760 => x"81",
          2761 => x"55",
          2762 => x"2e",
          2763 => x"87",
          2764 => x"08",
          2765 => x"70",
          2766 => x"54",
          2767 => x"2e",
          2768 => x"91",
          2769 => x"06",
          2770 => x"e3",
          2771 => x"32",
          2772 => x"72",
          2773 => x"38",
          2774 => x"81",
          2775 => x"cf",
          2776 => x"ff",
          2777 => x"c0",
          2778 => x"70",
          2779 => x"38",
          2780 => x"90",
          2781 => x"0c",
          2782 => x"84",
          2783 => x"0d",
          2784 => x"2a",
          2785 => x"51",
          2786 => x"38",
          2787 => x"81",
          2788 => x"80",
          2789 => x"71",
          2790 => x"06",
          2791 => x"2e",
          2792 => x"c0",
          2793 => x"70",
          2794 => x"81",
          2795 => x"52",
          2796 => x"d8",
          2797 => x"0d",
          2798 => x"33",
          2799 => x"9f",
          2800 => x"52",
          2801 => x"bc",
          2802 => x"0d",
          2803 => x"0d",
          2804 => x"75",
          2805 => x"52",
          2806 => x"2e",
          2807 => x"81",
          2808 => x"bc",
          2809 => x"ff",
          2810 => x"55",
          2811 => x"80",
          2812 => x"c0",
          2813 => x"70",
          2814 => x"81",
          2815 => x"52",
          2816 => x"8c",
          2817 => x"2a",
          2818 => x"51",
          2819 => x"38",
          2820 => x"81",
          2821 => x"80",
          2822 => x"71",
          2823 => x"06",
          2824 => x"38",
          2825 => x"06",
          2826 => x"94",
          2827 => x"80",
          2828 => x"87",
          2829 => x"52",
          2830 => x"81",
          2831 => x"55",
          2832 => x"9b",
          2833 => x"bb",
          2834 => x"3d",
          2835 => x"91",
          2836 => x"06",
          2837 => x"98",
          2838 => x"32",
          2839 => x"72",
          2840 => x"38",
          2841 => x"81",
          2842 => x"80",
          2843 => x"38",
          2844 => x"84",
          2845 => x"2a",
          2846 => x"53",
          2847 => x"ce",
          2848 => x"ff",
          2849 => x"c0",
          2850 => x"70",
          2851 => x"06",
          2852 => x"80",
          2853 => x"38",
          2854 => x"a4",
          2855 => x"c0",
          2856 => x"9e",
          2857 => x"f3",
          2858 => x"c0",
          2859 => x"83",
          2860 => x"87",
          2861 => x"08",
          2862 => x"0c",
          2863 => x"9c",
          2864 => x"d0",
          2865 => x"9e",
          2866 => x"f3",
          2867 => x"c0",
          2868 => x"83",
          2869 => x"87",
          2870 => x"08",
          2871 => x"0c",
          2872 => x"b4",
          2873 => x"e0",
          2874 => x"9e",
          2875 => x"f3",
          2876 => x"c0",
          2877 => x"83",
          2878 => x"87",
          2879 => x"08",
          2880 => x"0c",
          2881 => x"c4",
          2882 => x"f0",
          2883 => x"9e",
          2884 => x"71",
          2885 => x"23",
          2886 => x"84",
          2887 => x"f8",
          2888 => x"9e",
          2889 => x"f3",
          2890 => x"c0",
          2891 => x"83",
          2892 => x"81",
          2893 => x"84",
          2894 => x"87",
          2895 => x"08",
          2896 => x"0a",
          2897 => x"52",
          2898 => x"38",
          2899 => x"85",
          2900 => x"87",
          2901 => x"08",
          2902 => x"0a",
          2903 => x"52",
          2904 => x"83",
          2905 => x"71",
          2906 => x"34",
          2907 => x"c0",
          2908 => x"70",
          2909 => x"06",
          2910 => x"70",
          2911 => x"38",
          2912 => x"83",
          2913 => x"80",
          2914 => x"9e",
          2915 => x"88",
          2916 => x"51",
          2917 => x"80",
          2918 => x"81",
          2919 => x"f4",
          2920 => x"0b",
          2921 => x"90",
          2922 => x"80",
          2923 => x"52",
          2924 => x"2e",
          2925 => x"52",
          2926 => x"89",
          2927 => x"87",
          2928 => x"08",
          2929 => x"80",
          2930 => x"52",
          2931 => x"83",
          2932 => x"71",
          2933 => x"34",
          2934 => x"c0",
          2935 => x"70",
          2936 => x"06",
          2937 => x"70",
          2938 => x"38",
          2939 => x"83",
          2940 => x"80",
          2941 => x"9e",
          2942 => x"82",
          2943 => x"51",
          2944 => x"80",
          2945 => x"81",
          2946 => x"f4",
          2947 => x"0b",
          2948 => x"90",
          2949 => x"80",
          2950 => x"52",
          2951 => x"2e",
          2952 => x"52",
          2953 => x"8d",
          2954 => x"87",
          2955 => x"08",
          2956 => x"80",
          2957 => x"52",
          2958 => x"83",
          2959 => x"71",
          2960 => x"34",
          2961 => x"c0",
          2962 => x"70",
          2963 => x"51",
          2964 => x"80",
          2965 => x"81",
          2966 => x"f4",
          2967 => x"c0",
          2968 => x"98",
          2969 => x"8a",
          2970 => x"71",
          2971 => x"34",
          2972 => x"c0",
          2973 => x"70",
          2974 => x"51",
          2975 => x"80",
          2976 => x"81",
          2977 => x"f4",
          2978 => x"c0",
          2979 => x"83",
          2980 => x"84",
          2981 => x"71",
          2982 => x"34",
          2983 => x"c0",
          2984 => x"70",
          2985 => x"52",
          2986 => x"2e",
          2987 => x"52",
          2988 => x"93",
          2989 => x"9e",
          2990 => x"06",
          2991 => x"f4",
          2992 => x"3d",
          2993 => x"52",
          2994 => x"fb",
          2995 => x"da",
          2996 => x"b6",
          2997 => x"f4",
          2998 => x"73",
          2999 => x"83",
          3000 => x"c3",
          3001 => x"f4",
          3002 => x"74",
          3003 => x"83",
          3004 => x"54",
          3005 => x"38",
          3006 => x"33",
          3007 => x"9e",
          3008 => x"89",
          3009 => x"84",
          3010 => x"f4",
          3011 => x"73",
          3012 => x"83",
          3013 => x"56",
          3014 => x"38",
          3015 => x"33",
          3016 => x"86",
          3017 => x"91",
          3018 => x"83",
          3019 => x"f4",
          3020 => x"75",
          3021 => x"83",
          3022 => x"54",
          3023 => x"38",
          3024 => x"33",
          3025 => x"89",
          3026 => x"8d",
          3027 => x"82",
          3028 => x"f4",
          3029 => x"73",
          3030 => x"83",
          3031 => x"c2",
          3032 => x"f3",
          3033 => x"83",
          3034 => x"ff",
          3035 => x"83",
          3036 => x"52",
          3037 => x"51",
          3038 => x"3f",
          3039 => x"08",
          3040 => x"9c",
          3041 => x"80",
          3042 => x"c4",
          3043 => x"3f",
          3044 => x"22",
          3045 => x"cc",
          3046 => x"ec",
          3047 => x"f8",
          3048 => x"84",
          3049 => x"51",
          3050 => x"84",
          3051 => x"bd",
          3052 => x"76",
          3053 => x"54",
          3054 => x"08",
          3055 => x"f4",
          3056 => x"c4",
          3057 => x"8b",
          3058 => x"b9",
          3059 => x"86",
          3060 => x"85",
          3061 => x"0d",
          3062 => x"80",
          3063 => x"84",
          3064 => x"51",
          3065 => x"84",
          3066 => x"bd",
          3067 => x"76",
          3068 => x"54",
          3069 => x"08",
          3070 => x"a0",
          3071 => x"88",
          3072 => x"0d",
          3073 => x"fc",
          3074 => x"84",
          3075 => x"51",
          3076 => x"84",
          3077 => x"bd",
          3078 => x"76",
          3079 => x"54",
          3080 => x"08",
          3081 => x"cc",
          3082 => x"dc",
          3083 => x"86",
          3084 => x"80",
          3085 => x"38",
          3086 => x"83",
          3087 => x"c0",
          3088 => x"da",
          3089 => x"ab",
          3090 => x"e8",
          3091 => x"da",
          3092 => x"b3",
          3093 => x"f3",
          3094 => x"83",
          3095 => x"ff",
          3096 => x"83",
          3097 => x"52",
          3098 => x"51",
          3099 => x"3f",
          3100 => x"51",
          3101 => x"3f",
          3102 => x"22",
          3103 => x"cc",
          3104 => x"84",
          3105 => x"f8",
          3106 => x"84",
          3107 => x"51",
          3108 => x"84",
          3109 => x"bd",
          3110 => x"76",
          3111 => x"54",
          3112 => x"08",
          3113 => x"f4",
          3114 => x"dc",
          3115 => x"8b",
          3116 => x"80",
          3117 => x"38",
          3118 => x"83",
          3119 => x"ff",
          3120 => x"83",
          3121 => x"54",
          3122 => x"fd",
          3123 => x"eb",
          3124 => x"88",
          3125 => x"9b",
          3126 => x"8d",
          3127 => x"80",
          3128 => x"38",
          3129 => x"dd",
          3130 => x"bf",
          3131 => x"f4",
          3132 => x"74",
          3133 => x"d1",
          3134 => x"83",
          3135 => x"ff",
          3136 => x"83",
          3137 => x"54",
          3138 => x"fc",
          3139 => x"39",
          3140 => x"33",
          3141 => x"b4",
          3142 => x"ec",
          3143 => x"85",
          3144 => x"80",
          3145 => x"38",
          3146 => x"f4",
          3147 => x"83",
          3148 => x"ff",
          3149 => x"83",
          3150 => x"55",
          3151 => x"fb",
          3152 => x"39",
          3153 => x"33",
          3154 => x"f4",
          3155 => x"b8",
          3156 => x"93",
          3157 => x"80",
          3158 => x"38",
          3159 => x"f3",
          3160 => x"f3",
          3161 => x"54",
          3162 => x"94",
          3163 => x"98",
          3164 => x"8f",
          3165 => x"80",
          3166 => x"38",
          3167 => x"f3",
          3168 => x"f3",
          3169 => x"54",
          3170 => x"b0",
          3171 => x"f8",
          3172 => x"8a",
          3173 => x"80",
          3174 => x"38",
          3175 => x"f3",
          3176 => x"f3",
          3177 => x"54",
          3178 => x"cc",
          3179 => x"d8",
          3180 => x"89",
          3181 => x"80",
          3182 => x"38",
          3183 => x"f3",
          3184 => x"f3",
          3185 => x"54",
          3186 => x"e8",
          3187 => x"b8",
          3188 => x"88",
          3189 => x"80",
          3190 => x"38",
          3191 => x"f3",
          3192 => x"f3",
          3193 => x"54",
          3194 => x"84",
          3195 => x"98",
          3196 => x"8b",
          3197 => x"80",
          3198 => x"38",
          3199 => x"df",
          3200 => x"b0",
          3201 => x"da",
          3202 => x"bc",
          3203 => x"f4",
          3204 => x"74",
          3205 => x"d7",
          3206 => x"ff",
          3207 => x"8e",
          3208 => x"71",
          3209 => x"38",
          3210 => x"83",
          3211 => x"52",
          3212 => x"83",
          3213 => x"ff",
          3214 => x"83",
          3215 => x"83",
          3216 => x"ff",
          3217 => x"83",
          3218 => x"83",
          3219 => x"ff",
          3220 => x"83",
          3221 => x"83",
          3222 => x"ff",
          3223 => x"83",
          3224 => x"83",
          3225 => x"ff",
          3226 => x"83",
          3227 => x"83",
          3228 => x"ff",
          3229 => x"83",
          3230 => x"71",
          3231 => x"04",
          3232 => x"c0",
          3233 => x"04",
          3234 => x"08",
          3235 => x"84",
          3236 => x"3d",
          3237 => x"08",
          3238 => x"5a",
          3239 => x"57",
          3240 => x"83",
          3241 => x"51",
          3242 => x"3f",
          3243 => x"08",
          3244 => x"8b",
          3245 => x"0b",
          3246 => x"08",
          3247 => x"f8",
          3248 => x"82",
          3249 => x"84",
          3250 => x"80",
          3251 => x"76",
          3252 => x"3f",
          3253 => x"08",
          3254 => x"55",
          3255 => x"bb",
          3256 => x"8e",
          3257 => x"84",
          3258 => x"70",
          3259 => x"80",
          3260 => x"09",
          3261 => x"72",
          3262 => x"51",
          3263 => x"76",
          3264 => x"73",
          3265 => x"83",
          3266 => x"8c",
          3267 => x"51",
          3268 => x"3f",
          3269 => x"08",
          3270 => x"76",
          3271 => x"77",
          3272 => x"0c",
          3273 => x"04",
          3274 => x"51",
          3275 => x"3f",
          3276 => x"09",
          3277 => x"38",
          3278 => x"51",
          3279 => x"79",
          3280 => x"e4",
          3281 => x"08",
          3282 => x"84",
          3283 => x"76",
          3284 => x"e4",
          3285 => x"b0",
          3286 => x"84",
          3287 => x"a9",
          3288 => x"d8",
          3289 => x"3d",
          3290 => x"08",
          3291 => x"72",
          3292 => x"5a",
          3293 => x"2e",
          3294 => x"80",
          3295 => x"59",
          3296 => x"10",
          3297 => x"f8",
          3298 => x"52",
          3299 => x"98",
          3300 => x"84",
          3301 => x"52",
          3302 => x"ff",
          3303 => x"84",
          3304 => x"90",
          3305 => x"33",
          3306 => x"2e",
          3307 => x"73",
          3308 => x"38",
          3309 => x"81",
          3310 => x"54",
          3311 => x"c1",
          3312 => x"73",
          3313 => x"0c",
          3314 => x"04",
          3315 => x"aa",
          3316 => x"11",
          3317 => x"05",
          3318 => x"3f",
          3319 => x"08",
          3320 => x"38",
          3321 => x"78",
          3322 => x"fd",
          3323 => x"bb",
          3324 => x"ff",
          3325 => x"80",
          3326 => x"81",
          3327 => x"ff",
          3328 => x"82",
          3329 => x"f9",
          3330 => x"39",
          3331 => x"05",
          3332 => x"27",
          3333 => x"81",
          3334 => x"70",
          3335 => x"73",
          3336 => x"81",
          3337 => x"38",
          3338 => x"eb",
          3339 => x"8d",
          3340 => x"fe",
          3341 => x"84",
          3342 => x"53",
          3343 => x"08",
          3344 => x"84",
          3345 => x"bb",
          3346 => x"d0",
          3347 => x"ec",
          3348 => x"f8",
          3349 => x"82",
          3350 => x"84",
          3351 => x"80",
          3352 => x"77",
          3353 => x"c0",
          3354 => x"84",
          3355 => x"0b",
          3356 => x"08",
          3357 => x"84",
          3358 => x"ff",
          3359 => x"58",
          3360 => x"34",
          3361 => x"52",
          3362 => x"e3",
          3363 => x"ff",
          3364 => x"74",
          3365 => x"81",
          3366 => x"38",
          3367 => x"bb",
          3368 => x"3d",
          3369 => x"3d",
          3370 => x"08",
          3371 => x"ba",
          3372 => x"3d",
          3373 => x"08",
          3374 => x"42",
          3375 => x"b5",
          3376 => x"f4",
          3377 => x"75",
          3378 => x"34",
          3379 => x"08",
          3380 => x"38",
          3381 => x"ff",
          3382 => x"74",
          3383 => x"ed",
          3384 => x"2e",
          3385 => x"81",
          3386 => x"5a",
          3387 => x"8b",
          3388 => x"2e",
          3389 => x"94",
          3390 => x"40",
          3391 => x"ea",
          3392 => x"bb",
          3393 => x"2b",
          3394 => x"5b",
          3395 => x"2e",
          3396 => x"79",
          3397 => x"84",
          3398 => x"70",
          3399 => x"98",
          3400 => x"bc",
          3401 => x"2b",
          3402 => x"71",
          3403 => x"70",
          3404 => x"df",
          3405 => x"08",
          3406 => x"51",
          3407 => x"5a",
          3408 => x"5c",
          3409 => x"74",
          3410 => x"cd",
          3411 => x"27",
          3412 => x"75",
          3413 => x"29",
          3414 => x"05",
          3415 => x"57",
          3416 => x"24",
          3417 => x"75",
          3418 => x"82",
          3419 => x"80",
          3420 => x"e4",
          3421 => x"57",
          3422 => x"91",
          3423 => x"e0",
          3424 => x"70",
          3425 => x"78",
          3426 => x"b6",
          3427 => x"2e",
          3428 => x"84",
          3429 => x"81",
          3430 => x"2e",
          3431 => x"81",
          3432 => x"2b",
          3433 => x"84",
          3434 => x"70",
          3435 => x"97",
          3436 => x"2c",
          3437 => x"2b",
          3438 => x"11",
          3439 => x"5e",
          3440 => x"57",
          3441 => x"2e",
          3442 => x"76",
          3443 => x"34",
          3444 => x"a8",
          3445 => x"84",
          3446 => x"70",
          3447 => x"57",
          3448 => x"09",
          3449 => x"ab",
          3450 => x"2e",
          3451 => x"7d",
          3452 => x"39",
          3453 => x"ff",
          3454 => x"81",
          3455 => x"81",
          3456 => x"70",
          3457 => x"81",
          3458 => x"57",
          3459 => x"26",
          3460 => x"75",
          3461 => x"82",
          3462 => x"80",
          3463 => x"e4",
          3464 => x"57",
          3465 => x"ce",
          3466 => x"e0",
          3467 => x"70",
          3468 => x"78",
          3469 => x"bc",
          3470 => x"2e",
          3471 => x"fe",
          3472 => x"57",
          3473 => x"fe",
          3474 => x"c6",
          3475 => x"fd",
          3476 => x"57",
          3477 => x"38",
          3478 => x"c0",
          3479 => x"e2",
          3480 => x"7f",
          3481 => x"0c",
          3482 => x"95",
          3483 => x"38",
          3484 => x"83",
          3485 => x"57",
          3486 => x"83",
          3487 => x"08",
          3488 => x"0b",
          3489 => x"34",
          3490 => x"e2",
          3491 => x"39",
          3492 => x"33",
          3493 => x"2e",
          3494 => x"84",
          3495 => x"52",
          3496 => x"b5",
          3497 => x"e2",
          3498 => x"05",
          3499 => x"e2",
          3500 => x"c9",
          3501 => x"c8",
          3502 => x"ff",
          3503 => x"c4",
          3504 => x"55",
          3505 => x"fc",
          3506 => x"e6",
          3507 => x"81",
          3508 => x"84",
          3509 => x"7b",
          3510 => x"52",
          3511 => x"8e",
          3512 => x"39",
          3513 => x"90",
          3514 => x"92",
          3515 => x"7c",
          3516 => x"f4",
          3517 => x"08",
          3518 => x"8f",
          3519 => x"0b",
          3520 => x"34",
          3521 => x"84",
          3522 => x"84",
          3523 => x"56",
          3524 => x"2e",
          3525 => x"e6",
          3526 => x"88",
          3527 => x"ce",
          3528 => x"e8",
          3529 => x"51",
          3530 => x"3f",
          3531 => x"08",
          3532 => x"ff",
          3533 => x"84",
          3534 => x"ff",
          3535 => x"84",
          3536 => x"78",
          3537 => x"55",
          3538 => x"7b",
          3539 => x"b8",
          3540 => x"e2",
          3541 => x"a5",
          3542 => x"38",
          3543 => x"08",
          3544 => x"f1",
          3545 => x"70",
          3546 => x"58",
          3547 => x"26",
          3548 => x"10",
          3549 => x"98",
          3550 => x"57",
          3551 => x"bc",
          3552 => x"26",
          3553 => x"7c",
          3554 => x"f4",
          3555 => x"08",
          3556 => x"80",
          3557 => x"38",
          3558 => x"b7",
          3559 => x"bb",
          3560 => x"e2",
          3561 => x"bb",
          3562 => x"ff",
          3563 => x"53",
          3564 => x"51",
          3565 => x"3f",
          3566 => x"33",
          3567 => x"33",
          3568 => x"80",
          3569 => x"38",
          3570 => x"08",
          3571 => x"ff",
          3572 => x"84",
          3573 => x"52",
          3574 => x"b3",
          3575 => x"e6",
          3576 => x"88",
          3577 => x"86",
          3578 => x"c8",
          3579 => x"55",
          3580 => x"c8",
          3581 => x"ff",
          3582 => x"39",
          3583 => x"33",
          3584 => x"06",
          3585 => x"33",
          3586 => x"75",
          3587 => x"ed",
          3588 => x"e8",
          3589 => x"15",
          3590 => x"e2",
          3591 => x"16",
          3592 => x"55",
          3593 => x"3f",
          3594 => x"33",
          3595 => x"06",
          3596 => x"33",
          3597 => x"75",
          3598 => x"c1",
          3599 => x"e8",
          3600 => x"15",
          3601 => x"e2",
          3602 => x"16",
          3603 => x"55",
          3604 => x"3f",
          3605 => x"33",
          3606 => x"06",
          3607 => x"33",
          3608 => x"77",
          3609 => x"a9",
          3610 => x"39",
          3611 => x"33",
          3612 => x"33",
          3613 => x"76",
          3614 => x"38",
          3615 => x"7a",
          3616 => x"34",
          3617 => x"70",
          3618 => x"81",
          3619 => x"57",
          3620 => x"24",
          3621 => x"84",
          3622 => x"52",
          3623 => x"b1",
          3624 => x"e2",
          3625 => x"98",
          3626 => x"2c",
          3627 => x"33",
          3628 => x"56",
          3629 => x"f8",
          3630 => x"e6",
          3631 => x"88",
          3632 => x"aa",
          3633 => x"80",
          3634 => x"80",
          3635 => x"98",
          3636 => x"c4",
          3637 => x"59",
          3638 => x"f8",
          3639 => x"e6",
          3640 => x"88",
          3641 => x"86",
          3642 => x"80",
          3643 => x"80",
          3644 => x"98",
          3645 => x"c4",
          3646 => x"59",
          3647 => x"ff",
          3648 => x"f9",
          3649 => x"58",
          3650 => x"78",
          3651 => x"e8",
          3652 => x"33",
          3653 => x"d6",
          3654 => x"80",
          3655 => x"80",
          3656 => x"98",
          3657 => x"c4",
          3658 => x"55",
          3659 => x"fe",
          3660 => x"16",
          3661 => x"33",
          3662 => x"e6",
          3663 => x"77",
          3664 => x"b0",
          3665 => x"81",
          3666 => x"81",
          3667 => x"70",
          3668 => x"e2",
          3669 => x"57",
          3670 => x"24",
          3671 => x"fe",
          3672 => x"e2",
          3673 => x"74",
          3674 => x"91",
          3675 => x"e8",
          3676 => x"51",
          3677 => x"3f",
          3678 => x"33",
          3679 => x"76",
          3680 => x"34",
          3681 => x"06",
          3682 => x"84",
          3683 => x"7c",
          3684 => x"61",
          3685 => x"e8",
          3686 => x"51",
          3687 => x"3f",
          3688 => x"52",
          3689 => x"bb",
          3690 => x"84",
          3691 => x"06",
          3692 => x"da",
          3693 => x"c4",
          3694 => x"80",
          3695 => x"38",
          3696 => x"33",
          3697 => x"83",
          3698 => x"70",
          3699 => x"56",
          3700 => x"38",
          3701 => x"87",
          3702 => x"f4",
          3703 => x"18",
          3704 => x"59",
          3705 => x"3f",
          3706 => x"08",
          3707 => x"f4",
          3708 => x"10",
          3709 => x"9c",
          3710 => x"54",
          3711 => x"94",
          3712 => x"a0",
          3713 => x"f4",
          3714 => x"10",
          3715 => x"9c",
          3716 => x"57",
          3717 => x"8b",
          3718 => x"f4",
          3719 => x"75",
          3720 => x"38",
          3721 => x"33",
          3722 => x"2e",
          3723 => x"80",
          3724 => x"c8",
          3725 => x"84",
          3726 => x"7b",
          3727 => x"0c",
          3728 => x"04",
          3729 => x"33",
          3730 => x"2e",
          3731 => x"e6",
          3732 => x"88",
          3733 => x"96",
          3734 => x"e8",
          3735 => x"51",
          3736 => x"3f",
          3737 => x"08",
          3738 => x"ff",
          3739 => x"84",
          3740 => x"ff",
          3741 => x"84",
          3742 => x"61",
          3743 => x"55",
          3744 => x"83",
          3745 => x"ff",
          3746 => x"80",
          3747 => x"c8",
          3748 => x"84",
          3749 => x"f4",
          3750 => x"e2",
          3751 => x"81",
          3752 => x"56",
          3753 => x"f4",
          3754 => x"e2",
          3755 => x"05",
          3756 => x"e2",
          3757 => x"16",
          3758 => x"e2",
          3759 => x"e6",
          3760 => x"88",
          3761 => x"a6",
          3762 => x"c8",
          3763 => x"2b",
          3764 => x"84",
          3765 => x"5a",
          3766 => x"76",
          3767 => x"ef",
          3768 => x"e8",
          3769 => x"51",
          3770 => x"3f",
          3771 => x"33",
          3772 => x"70",
          3773 => x"e2",
          3774 => x"57",
          3775 => x"79",
          3776 => x"38",
          3777 => x"08",
          3778 => x"ff",
          3779 => x"74",
          3780 => x"29",
          3781 => x"05",
          3782 => x"84",
          3783 => x"5c",
          3784 => x"7a",
          3785 => x"38",
          3786 => x"08",
          3787 => x"ff",
          3788 => x"74",
          3789 => x"29",
          3790 => x"05",
          3791 => x"84",
          3792 => x"5c",
          3793 => x"75",
          3794 => x"38",
          3795 => x"7b",
          3796 => x"17",
          3797 => x"84",
          3798 => x"52",
          3799 => x"ff",
          3800 => x"75",
          3801 => x"29",
          3802 => x"05",
          3803 => x"84",
          3804 => x"44",
          3805 => x"62",
          3806 => x"38",
          3807 => x"81",
          3808 => x"34",
          3809 => x"08",
          3810 => x"51",
          3811 => x"3f",
          3812 => x"0a",
          3813 => x"0a",
          3814 => x"2c",
          3815 => x"33",
          3816 => x"61",
          3817 => x"a7",
          3818 => x"39",
          3819 => x"80",
          3820 => x"34",
          3821 => x"33",
          3822 => x"2e",
          3823 => x"e6",
          3824 => x"88",
          3825 => x"a6",
          3826 => x"e8",
          3827 => x"51",
          3828 => x"3f",
          3829 => x"08",
          3830 => x"ff",
          3831 => x"84",
          3832 => x"ff",
          3833 => x"84",
          3834 => x"7c",
          3835 => x"55",
          3836 => x"83",
          3837 => x"ff",
          3838 => x"80",
          3839 => x"c8",
          3840 => x"84",
          3841 => x"7b",
          3842 => x"0c",
          3843 => x"04",
          3844 => x"33",
          3845 => x"06",
          3846 => x"61",
          3847 => x"38",
          3848 => x"33",
          3849 => x"27",
          3850 => x"98",
          3851 => x"2c",
          3852 => x"76",
          3853 => x"7b",
          3854 => x"33",
          3855 => x"75",
          3856 => x"29",
          3857 => x"05",
          3858 => x"84",
          3859 => x"52",
          3860 => x"78",
          3861 => x"81",
          3862 => x"84",
          3863 => x"77",
          3864 => x"7c",
          3865 => x"3d",
          3866 => x"84",
          3867 => x"57",
          3868 => x"8b",
          3869 => x"56",
          3870 => x"c4",
          3871 => x"84",
          3872 => x"70",
          3873 => x"29",
          3874 => x"05",
          3875 => x"79",
          3876 => x"45",
          3877 => x"61",
          3878 => x"90",
          3879 => x"2b",
          3880 => x"78",
          3881 => x"5b",
          3882 => x"79",
          3883 => x"38",
          3884 => x"08",
          3885 => x"ff",
          3886 => x"75",
          3887 => x"29",
          3888 => x"05",
          3889 => x"84",
          3890 => x"57",
          3891 => x"75",
          3892 => x"38",
          3893 => x"08",
          3894 => x"ff",
          3895 => x"75",
          3896 => x"29",
          3897 => x"05",
          3898 => x"84",
          3899 => x"57",
          3900 => x"76",
          3901 => x"38",
          3902 => x"84",
          3903 => x"e2",
          3904 => x"bb",
          3905 => x"f4",
          3906 => x"bb",
          3907 => x"83",
          3908 => x"ff",
          3909 => x"83",
          3910 => x"55",
          3911 => x"38",
          3912 => x"f0",
          3913 => x"cf",
          3914 => x"39",
          3915 => x"08",
          3916 => x"70",
          3917 => x"ff",
          3918 => x"75",
          3919 => x"29",
          3920 => x"05",
          3921 => x"84",
          3922 => x"52",
          3923 => x"76",
          3924 => x"84",
          3925 => x"70",
          3926 => x"98",
          3927 => x"ff",
          3928 => x"5b",
          3929 => x"25",
          3930 => x"fe",
          3931 => x"f4",
          3932 => x"2e",
          3933 => x"83",
          3934 => x"93",
          3935 => x"55",
          3936 => x"ff",
          3937 => x"58",
          3938 => x"25",
          3939 => x"0b",
          3940 => x"34",
          3941 => x"08",
          3942 => x"2e",
          3943 => x"74",
          3944 => x"e5",
          3945 => x"ec",
          3946 => x"db",
          3947 => x"0b",
          3948 => x"0c",
          3949 => x"3d",
          3950 => x"c1",
          3951 => x"80",
          3952 => x"80",
          3953 => x"16",
          3954 => x"56",
          3955 => x"ff",
          3956 => x"ba",
          3957 => x"ff",
          3958 => x"84",
          3959 => x"84",
          3960 => x"84",
          3961 => x"81",
          3962 => x"05",
          3963 => x"7b",
          3964 => x"f6",
          3965 => x"84",
          3966 => x"84",
          3967 => x"57",
          3968 => x"80",
          3969 => x"38",
          3970 => x"08",
          3971 => x"ff",
          3972 => x"84",
          3973 => x"52",
          3974 => x"a6",
          3975 => x"e6",
          3976 => x"88",
          3977 => x"c6",
          3978 => x"c8",
          3979 => x"59",
          3980 => x"c8",
          3981 => x"ff",
          3982 => x"39",
          3983 => x"a9",
          3984 => x"bb",
          3985 => x"e2",
          3986 => x"bb",
          3987 => x"ff",
          3988 => x"53",
          3989 => x"51",
          3990 => x"3f",
          3991 => x"c4",
          3992 => x"c8",
          3993 => x"5d",
          3994 => x"f1",
          3995 => x"e6",
          3996 => x"88",
          3997 => x"f6",
          3998 => x"e8",
          3999 => x"51",
          4000 => x"3f",
          4001 => x"08",
          4002 => x"ff",
          4003 => x"84",
          4004 => x"ff",
          4005 => x"84",
          4006 => x"76",
          4007 => x"55",
          4008 => x"51",
          4009 => x"3f",
          4010 => x"08",
          4011 => x"34",
          4012 => x"08",
          4013 => x"81",
          4014 => x"52",
          4015 => x"a9",
          4016 => x"1d",
          4017 => x"06",
          4018 => x"33",
          4019 => x"33",
          4020 => x"56",
          4021 => x"f0",
          4022 => x"e6",
          4023 => x"88",
          4024 => x"8a",
          4025 => x"e8",
          4026 => x"51",
          4027 => x"3f",
          4028 => x"08",
          4029 => x"ff",
          4030 => x"84",
          4031 => x"ff",
          4032 => x"84",
          4033 => x"7a",
          4034 => x"55",
          4035 => x"7c",
          4036 => x"84",
          4037 => x"80",
          4038 => x"c4",
          4039 => x"bb",
          4040 => x"3d",
          4041 => x"f4",
          4042 => x"75",
          4043 => x"ce",
          4044 => x"ff",
          4045 => x"84",
          4046 => x"84",
          4047 => x"84",
          4048 => x"81",
          4049 => x"05",
          4050 => x"7b",
          4051 => x"9a",
          4052 => x"c4",
          4053 => x"c8",
          4054 => x"74",
          4055 => x"eb",
          4056 => x"e8",
          4057 => x"51",
          4058 => x"3f",
          4059 => x"08",
          4060 => x"ff",
          4061 => x"84",
          4062 => x"52",
          4063 => x"a3",
          4064 => x"e2",
          4065 => x"05",
          4066 => x"e2",
          4067 => x"81",
          4068 => x"c7",
          4069 => x"80",
          4070 => x"83",
          4071 => x"70",
          4072 => x"fc",
          4073 => x"9c",
          4074 => x"70",
          4075 => x"56",
          4076 => x"3f",
          4077 => x"08",
          4078 => x"f4",
          4079 => x"10",
          4080 => x"9c",
          4081 => x"54",
          4082 => x"94",
          4083 => x"94",
          4084 => x"f4",
          4085 => x"10",
          4086 => x"9c",
          4087 => x"57",
          4088 => x"80",
          4089 => x"38",
          4090 => x"52",
          4091 => x"a6",
          4092 => x"f4",
          4093 => x"05",
          4094 => x"06",
          4095 => x"75",
          4096 => x"38",
          4097 => x"f4",
          4098 => x"39",
          4099 => x"f8",
          4100 => x"53",
          4101 => x"51",
          4102 => x"3f",
          4103 => x"08",
          4104 => x"82",
          4105 => x"83",
          4106 => x"51",
          4107 => x"3f",
          4108 => x"e2",
          4109 => x"0b",
          4110 => x"34",
          4111 => x"84",
          4112 => x"0d",
          4113 => x"77",
          4114 => x"81",
          4115 => x"84",
          4116 => x"82",
          4117 => x"bb",
          4118 => x"3d",
          4119 => x"f4",
          4120 => x"80",
          4121 => x"51",
          4122 => x"3f",
          4123 => x"08",
          4124 => x"84",
          4125 => x"09",
          4126 => x"f5",
          4127 => x"84",
          4128 => x"a5",
          4129 => x"bb",
          4130 => x"80",
          4131 => x"84",
          4132 => x"fb",
          4133 => x"84",
          4134 => x"70",
          4135 => x"80",
          4136 => x"81",
          4137 => x"f4",
          4138 => x"10",
          4139 => x"9c",
          4140 => x"58",
          4141 => x"74",
          4142 => x"75",
          4143 => x"fc",
          4144 => x"9c",
          4145 => x"70",
          4146 => x"80",
          4147 => x"84",
          4148 => x"7f",
          4149 => x"f4",
          4150 => x"10",
          4151 => x"05",
          4152 => x"56",
          4153 => x"52",
          4154 => x"9c",
          4155 => x"f4",
          4156 => x"10",
          4157 => x"05",
          4158 => x"41",
          4159 => x"38",
          4160 => x"81",
          4161 => x"56",
          4162 => x"83",
          4163 => x"76",
          4164 => x"81",
          4165 => x"38",
          4166 => x"38",
          4167 => x"75",
          4168 => x"74",
          4169 => x"c2",
          4170 => x"f4",
          4171 => x"70",
          4172 => x"5b",
          4173 => x"27",
          4174 => x"80",
          4175 => x"f4",
          4176 => x"39",
          4177 => x"d4",
          4178 => x"f4",
          4179 => x"82",
          4180 => x"06",
          4181 => x"05",
          4182 => x"54",
          4183 => x"80",
          4184 => x"84",
          4185 => x"7f",
          4186 => x"f4",
          4187 => x"10",
          4188 => x"05",
          4189 => x"56",
          4190 => x"52",
          4191 => x"88",
          4192 => x"f4",
          4193 => x"10",
          4194 => x"05",
          4195 => x"41",
          4196 => x"2e",
          4197 => x"ff",
          4198 => x"83",
          4199 => x"fe",
          4200 => x"83",
          4201 => x"f0",
          4202 => x"e2",
          4203 => x"9d",
          4204 => x"e6",
          4205 => x"b6",
          4206 => x"0d",
          4207 => x"05",
          4208 => x"05",
          4209 => x"33",
          4210 => x"83",
          4211 => x"38",
          4212 => x"81",
          4213 => x"73",
          4214 => x"38",
          4215 => x"82",
          4216 => x"c7",
          4217 => x"86",
          4218 => x"70",
          4219 => x"56",
          4220 => x"79",
          4221 => x"38",
          4222 => x"b4",
          4223 => x"fa",
          4224 => x"83",
          4225 => x"83",
          4226 => x"70",
          4227 => x"90",
          4228 => x"88",
          4229 => x"07",
          4230 => x"56",
          4231 => x"77",
          4232 => x"80",
          4233 => x"05",
          4234 => x"73",
          4235 => x"55",
          4236 => x"26",
          4237 => x"78",
          4238 => x"83",
          4239 => x"84",
          4240 => x"79",
          4241 => x"55",
          4242 => x"e0",
          4243 => x"74",
          4244 => x"05",
          4245 => x"13",
          4246 => x"38",
          4247 => x"04",
          4248 => x"80",
          4249 => x"b4",
          4250 => x"10",
          4251 => x"b5",
          4252 => x"29",
          4253 => x"5b",
          4254 => x"59",
          4255 => x"80",
          4256 => x"f8",
          4257 => x"ff",
          4258 => x"f7",
          4259 => x"ff",
          4260 => x"b2",
          4261 => x"ff",
          4262 => x"75",
          4263 => x"5d",
          4264 => x"5b",
          4265 => x"26",
          4266 => x"74",
          4267 => x"56",
          4268 => x"06",
          4269 => x"06",
          4270 => x"06",
          4271 => x"ff",
          4272 => x"ff",
          4273 => x"29",
          4274 => x"57",
          4275 => x"74",
          4276 => x"38",
          4277 => x"33",
          4278 => x"05",
          4279 => x"1b",
          4280 => x"83",
          4281 => x"80",
          4282 => x"38",
          4283 => x"53",
          4284 => x"fe",
          4285 => x"73",
          4286 => x"55",
          4287 => x"b0",
          4288 => x"81",
          4289 => x"e8",
          4290 => x"a0",
          4291 => x"c7",
          4292 => x"84",
          4293 => x"70",
          4294 => x"84",
          4295 => x"70",
          4296 => x"83",
          4297 => x"70",
          4298 => x"5b",
          4299 => x"56",
          4300 => x"78",
          4301 => x"38",
          4302 => x"06",
          4303 => x"06",
          4304 => x"18",
          4305 => x"79",
          4306 => x"bb",
          4307 => x"83",
          4308 => x"80",
          4309 => x"b5",
          4310 => x"b0",
          4311 => x"2b",
          4312 => x"07",
          4313 => x"07",
          4314 => x"7f",
          4315 => x"5b",
          4316 => x"fd",
          4317 => x"be",
          4318 => x"e6",
          4319 => x"b4",
          4320 => x"ff",
          4321 => x"10",
          4322 => x"b5",
          4323 => x"29",
          4324 => x"a0",
          4325 => x"57",
          4326 => x"5f",
          4327 => x"80",
          4328 => x"b8",
          4329 => x"81",
          4330 => x"b8",
          4331 => x"81",
          4332 => x"fa",
          4333 => x"83",
          4334 => x"7c",
          4335 => x"05",
          4336 => x"5f",
          4337 => x"5e",
          4338 => x"26",
          4339 => x"7a",
          4340 => x"7d",
          4341 => x"53",
          4342 => x"06",
          4343 => x"06",
          4344 => x"7d",
          4345 => x"06",
          4346 => x"06",
          4347 => x"58",
          4348 => x"5d",
          4349 => x"26",
          4350 => x"75",
          4351 => x"73",
          4352 => x"83",
          4353 => x"79",
          4354 => x"76",
          4355 => x"7b",
          4356 => x"fb",
          4357 => x"78",
          4358 => x"56",
          4359 => x"fb",
          4360 => x"8e",
          4361 => x"ff",
          4362 => x"87",
          4363 => x"73",
          4364 => x"34",
          4365 => x"9c",
          4366 => x"75",
          4367 => x"75",
          4368 => x"80",
          4369 => x"76",
          4370 => x"34",
          4371 => x"94",
          4372 => x"34",
          4373 => x"ff",
          4374 => x"81",
          4375 => x"fa",
          4376 => x"c0",
          4377 => x"08",
          4378 => x"f8",
          4379 => x"81",
          4380 => x"06",
          4381 => x"55",
          4382 => x"73",
          4383 => x"ff",
          4384 => x"07",
          4385 => x"75",
          4386 => x"87",
          4387 => x"77",
          4388 => x"51",
          4389 => x"c0",
          4390 => x"73",
          4391 => x"06",
          4392 => x"72",
          4393 => x"d0",
          4394 => x"f8",
          4395 => x"84",
          4396 => x"87",
          4397 => x"84",
          4398 => x"84",
          4399 => x"04",
          4400 => x"02",
          4401 => x"02",
          4402 => x"05",
          4403 => x"f7",
          4404 => x"56",
          4405 => x"79",
          4406 => x"38",
          4407 => x"33",
          4408 => x"33",
          4409 => x"33",
          4410 => x"12",
          4411 => x"80",
          4412 => x"b2",
          4413 => x"57",
          4414 => x"29",
          4415 => x"ff",
          4416 => x"f9",
          4417 => x"57",
          4418 => x"81",
          4419 => x"38",
          4420 => x"22",
          4421 => x"74",
          4422 => x"23",
          4423 => x"33",
          4424 => x"81",
          4425 => x"81",
          4426 => x"5b",
          4427 => x"26",
          4428 => x"ff",
          4429 => x"83",
          4430 => x"83",
          4431 => x"70",
          4432 => x"06",
          4433 => x"33",
          4434 => x"79",
          4435 => x"89",
          4436 => x"f8",
          4437 => x"29",
          4438 => x"54",
          4439 => x"26",
          4440 => x"99",
          4441 => x"54",
          4442 => x"13",
          4443 => x"16",
          4444 => x"81",
          4445 => x"75",
          4446 => x"57",
          4447 => x"54",
          4448 => x"73",
          4449 => x"73",
          4450 => x"a1",
          4451 => x"b0",
          4452 => x"d6",
          4453 => x"a0",
          4454 => x"14",
          4455 => x"70",
          4456 => x"34",
          4457 => x"9f",
          4458 => x"eb",
          4459 => x"f6",
          4460 => x"56",
          4461 => x"b2",
          4462 => x"78",
          4463 => x"77",
          4464 => x"06",
          4465 => x"73",
          4466 => x"38",
          4467 => x"81",
          4468 => x"f8",
          4469 => x"29",
          4470 => x"75",
          4471 => x"a0",
          4472 => x"c7",
          4473 => x"81",
          4474 => x"81",
          4475 => x"71",
          4476 => x"5c",
          4477 => x"79",
          4478 => x"84",
          4479 => x"54",
          4480 => x"33",
          4481 => x"80",
          4482 => x"70",
          4483 => x"34",
          4484 => x"05",
          4485 => x"70",
          4486 => x"34",
          4487 => x"b8",
          4488 => x"b8",
          4489 => x"71",
          4490 => x"5c",
          4491 => x"75",
          4492 => x"80",
          4493 => x"bb",
          4494 => x"3d",
          4495 => x"83",
          4496 => x"83",
          4497 => x"70",
          4498 => x"06",
          4499 => x"33",
          4500 => x"73",
          4501 => x"f9",
          4502 => x"2e",
          4503 => x"78",
          4504 => x"ff",
          4505 => x"b4",
          4506 => x"72",
          4507 => x"81",
          4508 => x"38",
          4509 => x"81",
          4510 => x"f8",
          4511 => x"29",
          4512 => x"11",
          4513 => x"54",
          4514 => x"fe",
          4515 => x"fa",
          4516 => x"99",
          4517 => x"76",
          4518 => x"56",
          4519 => x"e0",
          4520 => x"75",
          4521 => x"57",
          4522 => x"53",
          4523 => x"fe",
          4524 => x"0b",
          4525 => x"34",
          4526 => x"81",
          4527 => x"ff",
          4528 => x"d8",
          4529 => x"39",
          4530 => x"b8",
          4531 => x"56",
          4532 => x"83",
          4533 => x"33",
          4534 => x"80",
          4535 => x"34",
          4536 => x"33",
          4537 => x"39",
          4538 => x"76",
          4539 => x"9f",
          4540 => x"51",
          4541 => x"9b",
          4542 => x"10",
          4543 => x"05",
          4544 => x"04",
          4545 => x"33",
          4546 => x"27",
          4547 => x"83",
          4548 => x"80",
          4549 => x"84",
          4550 => x"0d",
          4551 => x"83",
          4552 => x"83",
          4553 => x"70",
          4554 => x"54",
          4555 => x"2e",
          4556 => x"12",
          4557 => x"fa",
          4558 => x"0b",
          4559 => x"0c",
          4560 => x"04",
          4561 => x"33",
          4562 => x"70",
          4563 => x"2c",
          4564 => x"55",
          4565 => x"83",
          4566 => x"de",
          4567 => x"b4",
          4568 => x"84",
          4569 => x"ff",
          4570 => x"51",
          4571 => x"83",
          4572 => x"72",
          4573 => x"34",
          4574 => x"bb",
          4575 => x"3d",
          4576 => x"fa",
          4577 => x"73",
          4578 => x"70",
          4579 => x"06",
          4580 => x"55",
          4581 => x"b5",
          4582 => x"84",
          4583 => x"86",
          4584 => x"83",
          4585 => x"72",
          4586 => x"f8",
          4587 => x"55",
          4588 => x"74",
          4589 => x"70",
          4590 => x"fa",
          4591 => x"0b",
          4592 => x"0c",
          4593 => x"04",
          4594 => x"fa",
          4595 => x"fa",
          4596 => x"b8",
          4597 => x"05",
          4598 => x"75",
          4599 => x"38",
          4600 => x"70",
          4601 => x"34",
          4602 => x"ff",
          4603 => x"8f",
          4604 => x"70",
          4605 => x"38",
          4606 => x"83",
          4607 => x"51",
          4608 => x"83",
          4609 => x"70",
          4610 => x"71",
          4611 => x"f0",
          4612 => x"84",
          4613 => x"52",
          4614 => x"80",
          4615 => x"81",
          4616 => x"80",
          4617 => x"fa",
          4618 => x"0b",
          4619 => x"0c",
          4620 => x"04",
          4621 => x"33",
          4622 => x"90",
          4623 => x"83",
          4624 => x"80",
          4625 => x"84",
          4626 => x"0d",
          4627 => x"b0",
          4628 => x"07",
          4629 => x"fa",
          4630 => x"39",
          4631 => x"33",
          4632 => x"86",
          4633 => x"83",
          4634 => x"d7",
          4635 => x"0b",
          4636 => x"34",
          4637 => x"bb",
          4638 => x"3d",
          4639 => x"fa",
          4640 => x"fc",
          4641 => x"51",
          4642 => x"b0",
          4643 => x"39",
          4644 => x"33",
          4645 => x"70",
          4646 => x"34",
          4647 => x"83",
          4648 => x"81",
          4649 => x"07",
          4650 => x"fa",
          4651 => x"93",
          4652 => x"b0",
          4653 => x"06",
          4654 => x"70",
          4655 => x"34",
          4656 => x"83",
          4657 => x"81",
          4658 => x"07",
          4659 => x"fa",
          4660 => x"ef",
          4661 => x"b0",
          4662 => x"06",
          4663 => x"fa",
          4664 => x"df",
          4665 => x"b0",
          4666 => x"06",
          4667 => x"51",
          4668 => x"b0",
          4669 => x"39",
          4670 => x"33",
          4671 => x"b0",
          4672 => x"83",
          4673 => x"fe",
          4674 => x"fa",
          4675 => x"ef",
          4676 => x"07",
          4677 => x"fa",
          4678 => x"a7",
          4679 => x"b0",
          4680 => x"06",
          4681 => x"51",
          4682 => x"b0",
          4683 => x"39",
          4684 => x"33",
          4685 => x"a0",
          4686 => x"83",
          4687 => x"fe",
          4688 => x"fa",
          4689 => x"8f",
          4690 => x"83",
          4691 => x"fd",
          4692 => x"fa",
          4693 => x"fa",
          4694 => x"51",
          4695 => x"b0",
          4696 => x"39",
          4697 => x"02",
          4698 => x"02",
          4699 => x"c3",
          4700 => x"fa",
          4701 => x"fa",
          4702 => x"fa",
          4703 => x"b8",
          4704 => x"41",
          4705 => x"59",
          4706 => x"82",
          4707 => x"82",
          4708 => x"78",
          4709 => x"82",
          4710 => x"b8",
          4711 => x"0b",
          4712 => x"34",
          4713 => x"b4",
          4714 => x"fa",
          4715 => x"83",
          4716 => x"8f",
          4717 => x"78",
          4718 => x"81",
          4719 => x"80",
          4720 => x"fa",
          4721 => x"84",
          4722 => x"82",
          4723 => x"b4",
          4724 => x"83",
          4725 => x"82",
          4726 => x"b2",
          4727 => x"84",
          4728 => x"57",
          4729 => x"33",
          4730 => x"f6",
          4731 => x"54",
          4732 => x"52",
          4733 => x"51",
          4734 => x"3f",
          4735 => x"fa",
          4736 => x"84",
          4737 => x"7a",
          4738 => x"34",
          4739 => x"b2",
          4740 => x"fa",
          4741 => x"3d",
          4742 => x"0b",
          4743 => x"34",
          4744 => x"b8",
          4745 => x"0b",
          4746 => x"34",
          4747 => x"fa",
          4748 => x"0b",
          4749 => x"23",
          4750 => x"33",
          4751 => x"86",
          4752 => x"ba",
          4753 => x"79",
          4754 => x"7c",
          4755 => x"83",
          4756 => x"fe",
          4757 => x"80",
          4758 => x"85",
          4759 => x"79",
          4760 => x"38",
          4761 => x"ba",
          4762 => x"22",
          4763 => x"e5",
          4764 => x"ff",
          4765 => x"1a",
          4766 => x"06",
          4767 => x"33",
          4768 => x"78",
          4769 => x"38",
          4770 => x"51",
          4771 => x"3f",
          4772 => x"fa",
          4773 => x"84",
          4774 => x"7a",
          4775 => x"34",
          4776 => x"b2",
          4777 => x"fa",
          4778 => x"3d",
          4779 => x"0b",
          4780 => x"34",
          4781 => x"b8",
          4782 => x"0b",
          4783 => x"34",
          4784 => x"fa",
          4785 => x"0b",
          4786 => x"23",
          4787 => x"51",
          4788 => x"3f",
          4789 => x"08",
          4790 => x"b0",
          4791 => x"a8",
          4792 => x"83",
          4793 => x"ff",
          4794 => x"78",
          4795 => x"08",
          4796 => x"38",
          4797 => x"19",
          4798 => x"e5",
          4799 => x"fe",
          4800 => x"19",
          4801 => x"06",
          4802 => x"39",
          4803 => x"7a",
          4804 => x"a7",
          4805 => x"b8",
          4806 => x"fa",
          4807 => x"fa",
          4808 => x"71",
          4809 => x"c7",
          4810 => x"83",
          4811 => x"53",
          4812 => x"71",
          4813 => x"70",
          4814 => x"06",
          4815 => x"33",
          4816 => x"55",
          4817 => x"81",
          4818 => x"38",
          4819 => x"81",
          4820 => x"89",
          4821 => x"38",
          4822 => x"83",
          4823 => x"88",
          4824 => x"38",
          4825 => x"33",
          4826 => x"33",
          4827 => x"33",
          4828 => x"05",
          4829 => x"84",
          4830 => x"33",
          4831 => x"80",
          4832 => x"b8",
          4833 => x"fa",
          4834 => x"fa",
          4835 => x"71",
          4836 => x"5a",
          4837 => x"83",
          4838 => x"34",
          4839 => x"33",
          4840 => x"16",
          4841 => x"fa",
          4842 => x"c7",
          4843 => x"34",
          4844 => x"33",
          4845 => x"06",
          4846 => x"22",
          4847 => x"33",
          4848 => x"11",
          4849 => x"55",
          4850 => x"b0",
          4851 => x"d6",
          4852 => x"18",
          4853 => x"06",
          4854 => x"78",
          4855 => x"38",
          4856 => x"33",
          4857 => x"ea",
          4858 => x"53",
          4859 => x"b5",
          4860 => x"fb",
          4861 => x"80",
          4862 => x"84",
          4863 => x"57",
          4864 => x"80",
          4865 => x"0b",
          4866 => x"0c",
          4867 => x"04",
          4868 => x"97",
          4869 => x"24",
          4870 => x"75",
          4871 => x"81",
          4872 => x"38",
          4873 => x"51",
          4874 => x"80",
          4875 => x"b5",
          4876 => x"39",
          4877 => x"15",
          4878 => x"b9",
          4879 => x"74",
          4880 => x"2e",
          4881 => x"fe",
          4882 => x"53",
          4883 => x"51",
          4884 => x"81",
          4885 => x"ff",
          4886 => x"72",
          4887 => x"91",
          4888 => x"a0",
          4889 => x"3f",
          4890 => x"81",
          4891 => x"54",
          4892 => x"d8",
          4893 => x"39",
          4894 => x"b5",
          4895 => x"39",
          4896 => x"51",
          4897 => x"80",
          4898 => x"84",
          4899 => x"0d",
          4900 => x"ff",
          4901 => x"06",
          4902 => x"83",
          4903 => x"70",
          4904 => x"55",
          4905 => x"73",
          4906 => x"53",
          4907 => x"b5",
          4908 => x"a0",
          4909 => x"3f",
          4910 => x"33",
          4911 => x"06",
          4912 => x"53",
          4913 => x"38",
          4914 => x"83",
          4915 => x"fe",
          4916 => x"0b",
          4917 => x"34",
          4918 => x"51",
          4919 => x"fe",
          4920 => x"52",
          4921 => x"d8",
          4922 => x"39",
          4923 => x"02",
          4924 => x"33",
          4925 => x"08",
          4926 => x"81",
          4927 => x"38",
          4928 => x"83",
          4929 => x"8a",
          4930 => x"38",
          4931 => x"82",
          4932 => x"88",
          4933 => x"38",
          4934 => x"88",
          4935 => x"b8",
          4936 => x"fa",
          4937 => x"fa",
          4938 => x"72",
          4939 => x"5e",
          4940 => x"80",
          4941 => x"c7",
          4942 => x"34",
          4943 => x"33",
          4944 => x"33",
          4945 => x"22",
          4946 => x"12",
          4947 => x"40",
          4948 => x"b6",
          4949 => x"fa",
          4950 => x"71",
          4951 => x"40",
          4952 => x"b0",
          4953 => x"c7",
          4954 => x"34",
          4955 => x"33",
          4956 => x"06",
          4957 => x"22",
          4958 => x"33",
          4959 => x"11",
          4960 => x"58",
          4961 => x"b0",
          4962 => x"d6",
          4963 => x"1d",
          4964 => x"06",
          4965 => x"61",
          4966 => x"38",
          4967 => x"33",
          4968 => x"f1",
          4969 => x"56",
          4970 => x"b5",
          4971 => x"84",
          4972 => x"9c",
          4973 => x"78",
          4974 => x"8a",
          4975 => x"25",
          4976 => x"78",
          4977 => x"b3",
          4978 => x"db",
          4979 => x"38",
          4980 => x"ba",
          4981 => x"b8",
          4982 => x"fa",
          4983 => x"fa",
          4984 => x"72",
          4985 => x"40",
          4986 => x"80",
          4987 => x"c7",
          4988 => x"34",
          4989 => x"33",
          4990 => x"33",
          4991 => x"22",
          4992 => x"12",
          4993 => x"56",
          4994 => x"b6",
          4995 => x"fa",
          4996 => x"71",
          4997 => x"57",
          4998 => x"33",
          4999 => x"80",
          5000 => x"b8",
          5001 => x"81",
          5002 => x"fa",
          5003 => x"fa",
          5004 => x"72",
          5005 => x"42",
          5006 => x"83",
          5007 => x"60",
          5008 => x"05",
          5009 => x"58",
          5010 => x"06",
          5011 => x"27",
          5012 => x"77",
          5013 => x"34",
          5014 => x"bb",
          5015 => x"3d",
          5016 => x"9b",
          5017 => x"38",
          5018 => x"83",
          5019 => x"8d",
          5020 => x"06",
          5021 => x"80",
          5022 => x"b5",
          5023 => x"84",
          5024 => x"9c",
          5025 => x"78",
          5026 => x"aa",
          5027 => x"56",
          5028 => x"84",
          5029 => x"ba",
          5030 => x"11",
          5031 => x"84",
          5032 => x"78",
          5033 => x"18",
          5034 => x"ff",
          5035 => x"0b",
          5036 => x"1a",
          5037 => x"84",
          5038 => x"9c",
          5039 => x"78",
          5040 => x"e9",
          5041 => x"84",
          5042 => x"84",
          5043 => x"83",
          5044 => x"83",
          5045 => x"72",
          5046 => x"5e",
          5047 => x"b9",
          5048 => x"86",
          5049 => x"1d",
          5050 => x"f8",
          5051 => x"b5",
          5052 => x"b2",
          5053 => x"29",
          5054 => x"59",
          5055 => x"fa",
          5056 => x"83",
          5057 => x"76",
          5058 => x"5b",
          5059 => x"b0",
          5060 => x"b0",
          5061 => x"84",
          5062 => x"70",
          5063 => x"83",
          5064 => x"83",
          5065 => x"72",
          5066 => x"44",
          5067 => x"59",
          5068 => x"33",
          5069 => x"d6",
          5070 => x"1f",
          5071 => x"39",
          5072 => x"51",
          5073 => x"80",
          5074 => x"b5",
          5075 => x"39",
          5076 => x"33",
          5077 => x"33",
          5078 => x"06",
          5079 => x"33",
          5080 => x"12",
          5081 => x"80",
          5082 => x"b2",
          5083 => x"5d",
          5084 => x"05",
          5085 => x"ff",
          5086 => x"8a",
          5087 => x"59",
          5088 => x"81",
          5089 => x"38",
          5090 => x"06",
          5091 => x"57",
          5092 => x"38",
          5093 => x"83",
          5094 => x"fc",
          5095 => x"0b",
          5096 => x"34",
          5097 => x"ba",
          5098 => x"0b",
          5099 => x"34",
          5100 => x"ba",
          5101 => x"0b",
          5102 => x"0c",
          5103 => x"bb",
          5104 => x"3d",
          5105 => x"fa",
          5106 => x"ba",
          5107 => x"fa",
          5108 => x"ba",
          5109 => x"fa",
          5110 => x"ba",
          5111 => x"0b",
          5112 => x"0c",
          5113 => x"bb",
          5114 => x"3d",
          5115 => x"80",
          5116 => x"81",
          5117 => x"38",
          5118 => x"33",
          5119 => x"33",
          5120 => x"06",
          5121 => x"33",
          5122 => x"06",
          5123 => x"11",
          5124 => x"80",
          5125 => x"b2",
          5126 => x"72",
          5127 => x"70",
          5128 => x"06",
          5129 => x"33",
          5130 => x"5c",
          5131 => x"7d",
          5132 => x"fe",
          5133 => x"ff",
          5134 => x"58",
          5135 => x"38",
          5136 => x"83",
          5137 => x"7b",
          5138 => x"7a",
          5139 => x"78",
          5140 => x"72",
          5141 => x"5f",
          5142 => x"b9",
          5143 => x"c7",
          5144 => x"34",
          5145 => x"33",
          5146 => x"33",
          5147 => x"22",
          5148 => x"12",
          5149 => x"40",
          5150 => x"fa",
          5151 => x"83",
          5152 => x"60",
          5153 => x"05",
          5154 => x"fa",
          5155 => x"c7",
          5156 => x"34",
          5157 => x"33",
          5158 => x"06",
          5159 => x"22",
          5160 => x"33",
          5161 => x"11",
          5162 => x"5e",
          5163 => x"b0",
          5164 => x"99",
          5165 => x"81",
          5166 => x"ff",
          5167 => x"7c",
          5168 => x"ea",
          5169 => x"f9",
          5170 => x"96",
          5171 => x"19",
          5172 => x"fa",
          5173 => x"fa",
          5174 => x"81",
          5175 => x"ff",
          5176 => x"ac",
          5177 => x"2e",
          5178 => x"78",
          5179 => x"d7",
          5180 => x"2e",
          5181 => x"84",
          5182 => x"5f",
          5183 => x"38",
          5184 => x"56",
          5185 => x"84",
          5186 => x"10",
          5187 => x"e0",
          5188 => x"08",
          5189 => x"83",
          5190 => x"80",
          5191 => x"e7",
          5192 => x"0b",
          5193 => x"0c",
          5194 => x"04",
          5195 => x"33",
          5196 => x"33",
          5197 => x"06",
          5198 => x"33",
          5199 => x"06",
          5200 => x"11",
          5201 => x"80",
          5202 => x"b2",
          5203 => x"72",
          5204 => x"70",
          5205 => x"06",
          5206 => x"33",
          5207 => x"5c",
          5208 => x"7f",
          5209 => x"ef",
          5210 => x"7a",
          5211 => x"7a",
          5212 => x"7a",
          5213 => x"72",
          5214 => x"5c",
          5215 => x"b9",
          5216 => x"c7",
          5217 => x"34",
          5218 => x"33",
          5219 => x"33",
          5220 => x"22",
          5221 => x"12",
          5222 => x"56",
          5223 => x"fa",
          5224 => x"83",
          5225 => x"76",
          5226 => x"5a",
          5227 => x"b0",
          5228 => x"b0",
          5229 => x"84",
          5230 => x"70",
          5231 => x"83",
          5232 => x"83",
          5233 => x"72",
          5234 => x"5b",
          5235 => x"59",
          5236 => x"33",
          5237 => x"18",
          5238 => x"05",
          5239 => x"06",
          5240 => x"7a",
          5241 => x"38",
          5242 => x"33",
          5243 => x"fb",
          5244 => x"56",
          5245 => x"b5",
          5246 => x"70",
          5247 => x"5d",
          5248 => x"26",
          5249 => x"83",
          5250 => x"84",
          5251 => x"83",
          5252 => x"72",
          5253 => x"72",
          5254 => x"72",
          5255 => x"72",
          5256 => x"54",
          5257 => x"5b",
          5258 => x"a0",
          5259 => x"a0",
          5260 => x"84",
          5261 => x"83",
          5262 => x"83",
          5263 => x"72",
          5264 => x"5e",
          5265 => x"a0",
          5266 => x"b6",
          5267 => x"fa",
          5268 => x"71",
          5269 => x"5e",
          5270 => x"33",
          5271 => x"80",
          5272 => x"b8",
          5273 => x"81",
          5274 => x"fa",
          5275 => x"fa",
          5276 => x"72",
          5277 => x"44",
          5278 => x"83",
          5279 => x"84",
          5280 => x"34",
          5281 => x"70",
          5282 => x"5b",
          5283 => x"27",
          5284 => x"77",
          5285 => x"34",
          5286 => x"82",
          5287 => x"80",
          5288 => x"84",
          5289 => x"9c",
          5290 => x"83",
          5291 => x"33",
          5292 => x"80",
          5293 => x"34",
          5294 => x"33",
          5295 => x"06",
          5296 => x"56",
          5297 => x"81",
          5298 => x"86",
          5299 => x"84",
          5300 => x"9c",
          5301 => x"83",
          5302 => x"33",
          5303 => x"80",
          5304 => x"34",
          5305 => x"33",
          5306 => x"33",
          5307 => x"33",
          5308 => x"80",
          5309 => x"39",
          5310 => x"42",
          5311 => x"11",
          5312 => x"51",
          5313 => x"3f",
          5314 => x"08",
          5315 => x"f0",
          5316 => x"85",
          5317 => x"57",
          5318 => x"ba",
          5319 => x"10",
          5320 => x"41",
          5321 => x"05",
          5322 => x"ba",
          5323 => x"fb",
          5324 => x"fa",
          5325 => x"5c",
          5326 => x"1c",
          5327 => x"83",
          5328 => x"84",
          5329 => x"83",
          5330 => x"5b",
          5331 => x"e5",
          5332 => x"f8",
          5333 => x"b4",
          5334 => x"b5",
          5335 => x"29",
          5336 => x"5b",
          5337 => x"19",
          5338 => x"c7",
          5339 => x"34",
          5340 => x"33",
          5341 => x"33",
          5342 => x"22",
          5343 => x"12",
          5344 => x"56",
          5345 => x"b6",
          5346 => x"fa",
          5347 => x"71",
          5348 => x"5e",
          5349 => x"33",
          5350 => x"b0",
          5351 => x"84",
          5352 => x"70",
          5353 => x"83",
          5354 => x"83",
          5355 => x"72",
          5356 => x"41",
          5357 => x"5a",
          5358 => x"33",
          5359 => x"1e",
          5360 => x"70",
          5361 => x"5c",
          5362 => x"26",
          5363 => x"84",
          5364 => x"58",
          5365 => x"38",
          5366 => x"75",
          5367 => x"34",
          5368 => x"ba",
          5369 => x"b8",
          5370 => x"7f",
          5371 => x"bd",
          5372 => x"fc",
          5373 => x"f3",
          5374 => x"52",
          5375 => x"e4",
          5376 => x"84",
          5377 => x"9c",
          5378 => x"84",
          5379 => x"83",
          5380 => x"84",
          5381 => x"83",
          5382 => x"84",
          5383 => x"57",
          5384 => x"b2",
          5385 => x"39",
          5386 => x"33",
          5387 => x"34",
          5388 => x"33",
          5389 => x"34",
          5390 => x"33",
          5391 => x"34",
          5392 => x"84",
          5393 => x"5b",
          5394 => x"ff",
          5395 => x"ba",
          5396 => x"7c",
          5397 => x"81",
          5398 => x"38",
          5399 => x"33",
          5400 => x"83",
          5401 => x"81",
          5402 => x"53",
          5403 => x"52",
          5404 => x"52",
          5405 => x"b0",
          5406 => x"fe",
          5407 => x"84",
          5408 => x"81",
          5409 => x"f9",
          5410 => x"76",
          5411 => x"a0",
          5412 => x"38",
          5413 => x"f8",
          5414 => x"fb",
          5415 => x"c0",
          5416 => x"84",
          5417 => x"5b",
          5418 => x"ff",
          5419 => x"7b",
          5420 => x"38",
          5421 => x"ba",
          5422 => x"11",
          5423 => x"75",
          5424 => x"a5",
          5425 => x"10",
          5426 => x"05",
          5427 => x"04",
          5428 => x"33",
          5429 => x"2e",
          5430 => x"83",
          5431 => x"84",
          5432 => x"71",
          5433 => x"09",
          5434 => x"72",
          5435 => x"59",
          5436 => x"83",
          5437 => x"fd",
          5438 => x"ba",
          5439 => x"75",
          5440 => x"e7",
          5441 => x"d9",
          5442 => x"70",
          5443 => x"84",
          5444 => x"5d",
          5445 => x"7b",
          5446 => x"38",
          5447 => x"b5",
          5448 => x"39",
          5449 => x"fa",
          5450 => x"fa",
          5451 => x"81",
          5452 => x"57",
          5453 => x"fd",
          5454 => x"17",
          5455 => x"fa",
          5456 => x"9c",
          5457 => x"83",
          5458 => x"83",
          5459 => x"84",
          5460 => x"ff",
          5461 => x"76",
          5462 => x"84",
          5463 => x"56",
          5464 => x"b4",
          5465 => x"39",
          5466 => x"33",
          5467 => x"2e",
          5468 => x"83",
          5469 => x"84",
          5470 => x"71",
          5471 => x"09",
          5472 => x"72",
          5473 => x"59",
          5474 => x"83",
          5475 => x"fc",
          5476 => x"ba",
          5477 => x"7a",
          5478 => x"c4",
          5479 => x"d8",
          5480 => x"99",
          5481 => x"06",
          5482 => x"84",
          5483 => x"83",
          5484 => x"83",
          5485 => x"72",
          5486 => x"86",
          5487 => x"11",
          5488 => x"22",
          5489 => x"58",
          5490 => x"05",
          5491 => x"ff",
          5492 => x"88",
          5493 => x"fe",
          5494 => x"5a",
          5495 => x"84",
          5496 => x"92",
          5497 => x"0b",
          5498 => x"34",
          5499 => x"84",
          5500 => x"5a",
          5501 => x"fb",
          5502 => x"ba",
          5503 => x"77",
          5504 => x"81",
          5505 => x"38",
          5506 => x"f9",
          5507 => x"d0",
          5508 => x"85",
          5509 => x"80",
          5510 => x"38",
          5511 => x"33",
          5512 => x"33",
          5513 => x"84",
          5514 => x"ff",
          5515 => x"56",
          5516 => x"83",
          5517 => x"76",
          5518 => x"34",
          5519 => x"84",
          5520 => x"57",
          5521 => x"8c",
          5522 => x"ba",
          5523 => x"fa",
          5524 => x"61",
          5525 => x"f7",
          5526 => x"59",
          5527 => x"60",
          5528 => x"75",
          5529 => x"fa",
          5530 => x"f4",
          5531 => x"cc",
          5532 => x"94",
          5533 => x"84",
          5534 => x"57",
          5535 => x"27",
          5536 => x"76",
          5537 => x"d8",
          5538 => x"53",
          5539 => x"ac",
          5540 => x"f4",
          5541 => x"70",
          5542 => x"84",
          5543 => x"58",
          5544 => x"39",
          5545 => x"ba",
          5546 => x"57",
          5547 => x"8d",
          5548 => x"d8",
          5549 => x"83",
          5550 => x"75",
          5551 => x"76",
          5552 => x"51",
          5553 => x"fa",
          5554 => x"ba",
          5555 => x"81",
          5556 => x"b7",
          5557 => x"db",
          5558 => x"70",
          5559 => x"84",
          5560 => x"ff",
          5561 => x"ff",
          5562 => x"f7",
          5563 => x"ff",
          5564 => x"40",
          5565 => x"59",
          5566 => x"7e",
          5567 => x"77",
          5568 => x"fa",
          5569 => x"81",
          5570 => x"18",
          5571 => x"7f",
          5572 => x"77",
          5573 => x"fa",
          5574 => x"b8",
          5575 => x"11",
          5576 => x"60",
          5577 => x"38",
          5578 => x"83",
          5579 => x"f9",
          5580 => x"ba",
          5581 => x"7e",
          5582 => x"ef",
          5583 => x"d9",
          5584 => x"f7",
          5585 => x"7a",
          5586 => x"94",
          5587 => x"b4",
          5588 => x"f8",
          5589 => x"ff",
          5590 => x"b5",
          5591 => x"29",
          5592 => x"a0",
          5593 => x"fa",
          5594 => x"40",
          5595 => x"05",
          5596 => x"ff",
          5597 => x"8a",
          5598 => x"59",
          5599 => x"60",
          5600 => x"f0",
          5601 => x"ff",
          5602 => x"7c",
          5603 => x"80",
          5604 => x"fe",
          5605 => x"f7",
          5606 => x"76",
          5607 => x"38",
          5608 => x"75",
          5609 => x"23",
          5610 => x"06",
          5611 => x"41",
          5612 => x"24",
          5613 => x"84",
          5614 => x"56",
          5615 => x"8d",
          5616 => x"16",
          5617 => x"fa",
          5618 => x"81",
          5619 => x"fa",
          5620 => x"57",
          5621 => x"76",
          5622 => x"75",
          5623 => x"05",
          5624 => x"06",
          5625 => x"5c",
          5626 => x"58",
          5627 => x"80",
          5628 => x"b0",
          5629 => x"ff",
          5630 => x"ff",
          5631 => x"29",
          5632 => x"42",
          5633 => x"27",
          5634 => x"84",
          5635 => x"57",
          5636 => x"33",
          5637 => x"80",
          5638 => x"70",
          5639 => x"34",
          5640 => x"05",
          5641 => x"70",
          5642 => x"34",
          5643 => x"b8",
          5644 => x"b8",
          5645 => x"71",
          5646 => x"40",
          5647 => x"60",
          5648 => x"38",
          5649 => x"33",
          5650 => x"80",
          5651 => x"70",
          5652 => x"34",
          5653 => x"05",
          5654 => x"70",
          5655 => x"34",
          5656 => x"b8",
          5657 => x"b8",
          5658 => x"71",
          5659 => x"40",
          5660 => x"78",
          5661 => x"38",
          5662 => x"84",
          5663 => x"56",
          5664 => x"87",
          5665 => x"52",
          5666 => x"33",
          5667 => x"3f",
          5668 => x"80",
          5669 => x"f8",
          5670 => x"84",
          5671 => x"5d",
          5672 => x"79",
          5673 => x"38",
          5674 => x"22",
          5675 => x"2e",
          5676 => x"8b",
          5677 => x"fa",
          5678 => x"76",
          5679 => x"83",
          5680 => x"79",
          5681 => x"76",
          5682 => x"ed",
          5683 => x"f7",
          5684 => x"60",
          5685 => x"38",
          5686 => x"06",
          5687 => x"26",
          5688 => x"7b",
          5689 => x"7d",
          5690 => x"76",
          5691 => x"7a",
          5692 => x"70",
          5693 => x"05",
          5694 => x"80",
          5695 => x"5d",
          5696 => x"b0",
          5697 => x"83",
          5698 => x"5d",
          5699 => x"38",
          5700 => x"57",
          5701 => x"38",
          5702 => x"33",
          5703 => x"71",
          5704 => x"71",
          5705 => x"71",
          5706 => x"59",
          5707 => x"77",
          5708 => x"38",
          5709 => x"84",
          5710 => x"7d",
          5711 => x"05",
          5712 => x"77",
          5713 => x"84",
          5714 => x"84",
          5715 => x"41",
          5716 => x"ff",
          5717 => x"ff",
          5718 => x"b2",
          5719 => x"29",
          5720 => x"59",
          5721 => x"77",
          5722 => x"76",
          5723 => x"70",
          5724 => x"05",
          5725 => x"76",
          5726 => x"76",
          5727 => x"e0",
          5728 => x"b0",
          5729 => x"d6",
          5730 => x"a0",
          5731 => x"19",
          5732 => x"70",
          5733 => x"34",
          5734 => x"76",
          5735 => x"c0",
          5736 => x"e0",
          5737 => x"79",
          5738 => x"05",
          5739 => x"17",
          5740 => x"27",
          5741 => x"a8",
          5742 => x"70",
          5743 => x"5d",
          5744 => x"39",
          5745 => x"33",
          5746 => x"06",
          5747 => x"80",
          5748 => x"84",
          5749 => x"5d",
          5750 => x"f0",
          5751 => x"06",
          5752 => x"f2",
          5753 => x"b0",
          5754 => x"70",
          5755 => x"59",
          5756 => x"39",
          5757 => x"17",
          5758 => x"b9",
          5759 => x"7c",
          5760 => x"b4",
          5761 => x"f8",
          5762 => x"b2",
          5763 => x"f7",
          5764 => x"5f",
          5765 => x"39",
          5766 => x"33",
          5767 => x"75",
          5768 => x"34",
          5769 => x"81",
          5770 => x"56",
          5771 => x"83",
          5772 => x"81",
          5773 => x"07",
          5774 => x"fa",
          5775 => x"39",
          5776 => x"33",
          5777 => x"83",
          5778 => x"83",
          5779 => x"d4",
          5780 => x"b0",
          5781 => x"06",
          5782 => x"75",
          5783 => x"34",
          5784 => x"fa",
          5785 => x"9f",
          5786 => x"56",
          5787 => x"b0",
          5788 => x"39",
          5789 => x"83",
          5790 => x"81",
          5791 => x"ff",
          5792 => x"f4",
          5793 => x"fa",
          5794 => x"8f",
          5795 => x"83",
          5796 => x"ff",
          5797 => x"fa",
          5798 => x"9f",
          5799 => x"56",
          5800 => x"b0",
          5801 => x"39",
          5802 => x"33",
          5803 => x"80",
          5804 => x"75",
          5805 => x"34",
          5806 => x"83",
          5807 => x"81",
          5808 => x"c0",
          5809 => x"83",
          5810 => x"fe",
          5811 => x"fa",
          5812 => x"af",
          5813 => x"56",
          5814 => x"b0",
          5815 => x"39",
          5816 => x"33",
          5817 => x"86",
          5818 => x"83",
          5819 => x"fe",
          5820 => x"fa",
          5821 => x"fc",
          5822 => x"56",
          5823 => x"b0",
          5824 => x"39",
          5825 => x"33",
          5826 => x"82",
          5827 => x"83",
          5828 => x"fe",
          5829 => x"fa",
          5830 => x"f8",
          5831 => x"83",
          5832 => x"fd",
          5833 => x"fa",
          5834 => x"f0",
          5835 => x"83",
          5836 => x"fd",
          5837 => x"fa",
          5838 => x"f0",
          5839 => x"83",
          5840 => x"fd",
          5841 => x"fa",
          5842 => x"df",
          5843 => x"07",
          5844 => x"fa",
          5845 => x"cc",
          5846 => x"b0",
          5847 => x"06",
          5848 => x"75",
          5849 => x"34",
          5850 => x"80",
          5851 => x"b5",
          5852 => x"81",
          5853 => x"3f",
          5854 => x"84",
          5855 => x"83",
          5856 => x"84",
          5857 => x"83",
          5858 => x"84",
          5859 => x"59",
          5860 => x"b2",
          5861 => x"84",
          5862 => x"e8",
          5863 => x"0b",
          5864 => x"34",
          5865 => x"bb",
          5866 => x"3d",
          5867 => x"83",
          5868 => x"83",
          5869 => x"70",
          5870 => x"58",
          5871 => x"e7",
          5872 => x"ba",
          5873 => x"3d",
          5874 => x"d8",
          5875 => x"f7",
          5876 => x"bb",
          5877 => x"38",
          5878 => x"08",
          5879 => x"0c",
          5880 => x"ba",
          5881 => x"0b",
          5882 => x"0c",
          5883 => x"04",
          5884 => x"b5",
          5885 => x"39",
          5886 => x"33",
          5887 => x"5c",
          5888 => x"85",
          5889 => x"83",
          5890 => x"02",
          5891 => x"22",
          5892 => x"1e",
          5893 => x"84",
          5894 => x"ca",
          5895 => x"83",
          5896 => x"80",
          5897 => x"d1",
          5898 => x"fa",
          5899 => x"81",
          5900 => x"ff",
          5901 => x"d8",
          5902 => x"83",
          5903 => x"80",
          5904 => x"d0",
          5905 => x"98",
          5906 => x"fe",
          5907 => x"ef",
          5908 => x"fa",
          5909 => x"05",
          5910 => x"9f",
          5911 => x"58",
          5912 => x"a6",
          5913 => x"81",
          5914 => x"84",
          5915 => x"40",
          5916 => x"ee",
          5917 => x"83",
          5918 => x"ee",
          5919 => x"fa",
          5920 => x"05",
          5921 => x"9f",
          5922 => x"58",
          5923 => x"e2",
          5924 => x"b4",
          5925 => x"84",
          5926 => x"ff",
          5927 => x"56",
          5928 => x"f3",
          5929 => x"57",
          5930 => x"84",
          5931 => x"70",
          5932 => x"58",
          5933 => x"26",
          5934 => x"83",
          5935 => x"84",
          5936 => x"70",
          5937 => x"83",
          5938 => x"71",
          5939 => x"86",
          5940 => x"05",
          5941 => x"22",
          5942 => x"7e",
          5943 => x"83",
          5944 => x"83",
          5945 => x"5d",
          5946 => x"5f",
          5947 => x"2e",
          5948 => x"79",
          5949 => x"06",
          5950 => x"57",
          5951 => x"84",
          5952 => x"b8",
          5953 => x"76",
          5954 => x"98",
          5955 => x"56",
          5956 => x"b2",
          5957 => x"ff",
          5958 => x"57",
          5959 => x"24",
          5960 => x"84",
          5961 => x"56",
          5962 => x"82",
          5963 => x"16",
          5964 => x"fa",
          5965 => x"81",
          5966 => x"fa",
          5967 => x"57",
          5968 => x"76",
          5969 => x"75",
          5970 => x"05",
          5971 => x"06",
          5972 => x"5c",
          5973 => x"58",
          5974 => x"80",
          5975 => x"b0",
          5976 => x"ff",
          5977 => x"ff",
          5978 => x"29",
          5979 => x"42",
          5980 => x"27",
          5981 => x"84",
          5982 => x"57",
          5983 => x"33",
          5984 => x"80",
          5985 => x"70",
          5986 => x"34",
          5987 => x"05",
          5988 => x"70",
          5989 => x"34",
          5990 => x"b8",
          5991 => x"b8",
          5992 => x"71",
          5993 => x"41",
          5994 => x"76",
          5995 => x"38",
          5996 => x"33",
          5997 => x"80",
          5998 => x"70",
          5999 => x"34",
          6000 => x"05",
          6001 => x"70",
          6002 => x"34",
          6003 => x"b8",
          6004 => x"b8",
          6005 => x"71",
          6006 => x"41",
          6007 => x"78",
          6008 => x"38",
          6009 => x"83",
          6010 => x"33",
          6011 => x"80",
          6012 => x"34",
          6013 => x"33",
          6014 => x"33",
          6015 => x"22",
          6016 => x"33",
          6017 => x"5d",
          6018 => x"76",
          6019 => x"84",
          6020 => x"70",
          6021 => x"ff",
          6022 => x"58",
          6023 => x"83",
          6024 => x"79",
          6025 => x"23",
          6026 => x"06",
          6027 => x"5a",
          6028 => x"83",
          6029 => x"76",
          6030 => x"34",
          6031 => x"33",
          6032 => x"06",
          6033 => x"59",
          6034 => x"27",
          6035 => x"80",
          6036 => x"fa",
          6037 => x"88",
          6038 => x"b5",
          6039 => x"84",
          6040 => x"ff",
          6041 => x"56",
          6042 => x"ef",
          6043 => x"57",
          6044 => x"75",
          6045 => x"81",
          6046 => x"38",
          6047 => x"33",
          6048 => x"06",
          6049 => x"33",
          6050 => x"5d",
          6051 => x"2e",
          6052 => x"f4",
          6053 => x"a1",
          6054 => x"56",
          6055 => x"b4",
          6056 => x"39",
          6057 => x"75",
          6058 => x"23",
          6059 => x"7c",
          6060 => x"75",
          6061 => x"34",
          6062 => x"77",
          6063 => x"77",
          6064 => x"8d",
          6065 => x"70",
          6066 => x"34",
          6067 => x"33",
          6068 => x"05",
          6069 => x"7a",
          6070 => x"38",
          6071 => x"81",
          6072 => x"83",
          6073 => x"77",
          6074 => x"59",
          6075 => x"27",
          6076 => x"d3",
          6077 => x"31",
          6078 => x"fa",
          6079 => x"a8",
          6080 => x"83",
          6081 => x"fc",
          6082 => x"83",
          6083 => x"fc",
          6084 => x"0b",
          6085 => x"23",
          6086 => x"80",
          6087 => x"b4",
          6088 => x"39",
          6089 => x"18",
          6090 => x"b9",
          6091 => x"77",
          6092 => x"83",
          6093 => x"e9",
          6094 => x"3d",
          6095 => x"05",
          6096 => x"fa",
          6097 => x"72",
          6098 => x"38",
          6099 => x"9c",
          6100 => x"84",
          6101 => x"85",
          6102 => x"76",
          6103 => x"d7",
          6104 => x"0b",
          6105 => x"0c",
          6106 => x"04",
          6107 => x"02",
          6108 => x"5c",
          6109 => x"f9",
          6110 => x"81",
          6111 => x"f8",
          6112 => x"58",
          6113 => x"74",
          6114 => x"d6",
          6115 => x"56",
          6116 => x"88",
          6117 => x"78",
          6118 => x"0c",
          6119 => x"04",
          6120 => x"08",
          6121 => x"73",
          6122 => x"38",
          6123 => x"70",
          6124 => x"70",
          6125 => x"2a",
          6126 => x"58",
          6127 => x"e4",
          6128 => x"80",
          6129 => x"2e",
          6130 => x"83",
          6131 => x"7b",
          6132 => x"30",
          6133 => x"76",
          6134 => x"5d",
          6135 => x"85",
          6136 => x"b8",
          6137 => x"fa",
          6138 => x"fa",
          6139 => x"71",
          6140 => x"c7",
          6141 => x"83",
          6142 => x"5b",
          6143 => x"79",
          6144 => x"83",
          6145 => x"83",
          6146 => x"58",
          6147 => x"74",
          6148 => x"8c",
          6149 => x"54",
          6150 => x"80",
          6151 => x"0b",
          6152 => x"88",
          6153 => x"98",
          6154 => x"75",
          6155 => x"38",
          6156 => x"84",
          6157 => x"83",
          6158 => x"34",
          6159 => x"81",
          6160 => x"55",
          6161 => x"27",
          6162 => x"54",
          6163 => x"14",
          6164 => x"ff",
          6165 => x"ae",
          6166 => x"54",
          6167 => x"2e",
          6168 => x"72",
          6169 => x"86",
          6170 => x"83",
          6171 => x"34",
          6172 => x"06",
          6173 => x"ff",
          6174 => x"38",
          6175 => x"c2",
          6176 => x"f8",
          6177 => x"83",
          6178 => x"34",
          6179 => x"81",
          6180 => x"5e",
          6181 => x"ff",
          6182 => x"f8",
          6183 => x"98",
          6184 => x"25",
          6185 => x"75",
          6186 => x"34",
          6187 => x"06",
          6188 => x"81",
          6189 => x"06",
          6190 => x"72",
          6191 => x"e7",
          6192 => x"83",
          6193 => x"73",
          6194 => x"53",
          6195 => x"85",
          6196 => x"0b",
          6197 => x"34",
          6198 => x"f8",
          6199 => x"f8",
          6200 => x"f8",
          6201 => x"83",
          6202 => x"83",
          6203 => x"5d",
          6204 => x"5c",
          6205 => x"f8",
          6206 => x"55",
          6207 => x"2e",
          6208 => x"f8",
          6209 => x"54",
          6210 => x"82",
          6211 => x"f8",
          6212 => x"53",
          6213 => x"2e",
          6214 => x"f8",
          6215 => x"54",
          6216 => x"38",
          6217 => x"06",
          6218 => x"ff",
          6219 => x"83",
          6220 => x"33",
          6221 => x"2e",
          6222 => x"74",
          6223 => x"53",
          6224 => x"2e",
          6225 => x"83",
          6226 => x"33",
          6227 => x"27",
          6228 => x"83",
          6229 => x"87",
          6230 => x"c0",
          6231 => x"54",
          6232 => x"27",
          6233 => x"81",
          6234 => x"98",
          6235 => x"f8",
          6236 => x"81",
          6237 => x"ff",
          6238 => x"89",
          6239 => x"f6",
          6240 => x"f8",
          6241 => x"83",
          6242 => x"fe",
          6243 => x"72",
          6244 => x"8b",
          6245 => x"10",
          6246 => x"05",
          6247 => x"04",
          6248 => x"08",
          6249 => x"2e",
          6250 => x"f4",
          6251 => x"98",
          6252 => x"5e",
          6253 => x"fc",
          6254 => x"0b",
          6255 => x"33",
          6256 => x"81",
          6257 => x"74",
          6258 => x"f9",
          6259 => x"c0",
          6260 => x"83",
          6261 => x"73",
          6262 => x"58",
          6263 => x"94",
          6264 => x"b6",
          6265 => x"84",
          6266 => x"33",
          6267 => x"f0",
          6268 => x"39",
          6269 => x"08",
          6270 => x"2e",
          6271 => x"72",
          6272 => x"f4",
          6273 => x"76",
          6274 => x"54",
          6275 => x"80",
          6276 => x"39",
          6277 => x"57",
          6278 => x"81",
          6279 => x"79",
          6280 => x"81",
          6281 => x"38",
          6282 => x"80",
          6283 => x"81",
          6284 => x"38",
          6285 => x"06",
          6286 => x"27",
          6287 => x"54",
          6288 => x"25",
          6289 => x"80",
          6290 => x"81",
          6291 => x"ff",
          6292 => x"81",
          6293 => x"72",
          6294 => x"2b",
          6295 => x"58",
          6296 => x"24",
          6297 => x"10",
          6298 => x"10",
          6299 => x"83",
          6300 => x"83",
          6301 => x"70",
          6302 => x"54",
          6303 => x"98",
          6304 => x"f8",
          6305 => x"fd",
          6306 => x"59",
          6307 => x"ff",
          6308 => x"81",
          6309 => x"ff",
          6310 => x"59",
          6311 => x"78",
          6312 => x"9f",
          6313 => x"84",
          6314 => x"54",
          6315 => x"2e",
          6316 => x"7b",
          6317 => x"30",
          6318 => x"76",
          6319 => x"56",
          6320 => x"7b",
          6321 => x"81",
          6322 => x"38",
          6323 => x"f9",
          6324 => x"53",
          6325 => x"10",
          6326 => x"05",
          6327 => x"54",
          6328 => x"83",
          6329 => x"13",
          6330 => x"06",
          6331 => x"73",
          6332 => x"84",
          6333 => x"53",
          6334 => x"f9",
          6335 => x"b8",
          6336 => x"74",
          6337 => x"78",
          6338 => x"52",
          6339 => x"d4",
          6340 => x"bb",
          6341 => x"3d",
          6342 => x"76",
          6343 => x"54",
          6344 => x"72",
          6345 => x"92",
          6346 => x"cc",
          6347 => x"05",
          6348 => x"f8",
          6349 => x"fa",
          6350 => x"0b",
          6351 => x"15",
          6352 => x"83",
          6353 => x"34",
          6354 => x"f8",
          6355 => x"fa",
          6356 => x"81",
          6357 => x"72",
          6358 => x"fc",
          6359 => x"f8",
          6360 => x"55",
          6361 => x"fc",
          6362 => x"81",
          6363 => x"73",
          6364 => x"81",
          6365 => x"38",
          6366 => x"08",
          6367 => x"87",
          6368 => x"08",
          6369 => x"73",
          6370 => x"38",
          6371 => x"9c",
          6372 => x"d8",
          6373 => x"ff",
          6374 => x"d7",
          6375 => x"83",
          6376 => x"34",
          6377 => x"72",
          6378 => x"34",
          6379 => x"06",
          6380 => x"9e",
          6381 => x"f8",
          6382 => x"0b",
          6383 => x"33",
          6384 => x"08",
          6385 => x"33",
          6386 => x"e0",
          6387 => x"df",
          6388 => x"42",
          6389 => x"56",
          6390 => x"79",
          6391 => x"81",
          6392 => x"38",
          6393 => x"81",
          6394 => x"38",
          6395 => x"09",
          6396 => x"c0",
          6397 => x"39",
          6398 => x"81",
          6399 => x"98",
          6400 => x"84",
          6401 => x"57",
          6402 => x"38",
          6403 => x"84",
          6404 => x"ff",
          6405 => x"39",
          6406 => x"b8",
          6407 => x"54",
          6408 => x"81",
          6409 => x"b8",
          6410 => x"59",
          6411 => x"81",
          6412 => x"e4",
          6413 => x"f7",
          6414 => x"0b",
          6415 => x"0c",
          6416 => x"84",
          6417 => x"70",
          6418 => x"ff",
          6419 => x"54",
          6420 => x"83",
          6421 => x"74",
          6422 => x"23",
          6423 => x"06",
          6424 => x"53",
          6425 => x"83",
          6426 => x"73",
          6427 => x"34",
          6428 => x"33",
          6429 => x"06",
          6430 => x"53",
          6431 => x"83",
          6432 => x"72",
          6433 => x"34",
          6434 => x"b7",
          6435 => x"83",
          6436 => x"a5",
          6437 => x"f6",
          6438 => x"54",
          6439 => x"84",
          6440 => x"83",
          6441 => x"fe",
          6442 => x"81",
          6443 => x"88",
          6444 => x"e8",
          6445 => x"bb",
          6446 => x"0d",
          6447 => x"ac",
          6448 => x"0d",
          6449 => x"0d",
          6450 => x"f5",
          6451 => x"57",
          6452 => x"33",
          6453 => x"83",
          6454 => x"51",
          6455 => x"34",
          6456 => x"f5",
          6457 => x"56",
          6458 => x"15",
          6459 => x"87",
          6460 => x"34",
          6461 => x"9c",
          6462 => x"90",
          6463 => x"ce",
          6464 => x"87",
          6465 => x"08",
          6466 => x"98",
          6467 => x"70",
          6468 => x"38",
          6469 => x"87",
          6470 => x"08",
          6471 => x"73",
          6472 => x"71",
          6473 => x"db",
          6474 => x"98",
          6475 => x"ff",
          6476 => x"27",
          6477 => x"71",
          6478 => x"2e",
          6479 => x"87",
          6480 => x"08",
          6481 => x"05",
          6482 => x"98",
          6483 => x"87",
          6484 => x"08",
          6485 => x"2e",
          6486 => x"14",
          6487 => x"98",
          6488 => x"52",
          6489 => x"87",
          6490 => x"ff",
          6491 => x"87",
          6492 => x"08",
          6493 => x"26",
          6494 => x"52",
          6495 => x"16",
          6496 => x"06",
          6497 => x"80",
          6498 => x"74",
          6499 => x"52",
          6500 => x"38",
          6501 => x"8a",
          6502 => x"bb",
          6503 => x"3d",
          6504 => x"0b",
          6505 => x"0c",
          6506 => x"04",
          6507 => x"79",
          6508 => x"a3",
          6509 => x"52",
          6510 => x"f5",
          6511 => x"88",
          6512 => x"80",
          6513 => x"75",
          6514 => x"51",
          6515 => x"71",
          6516 => x"72",
          6517 => x"70",
          6518 => x"71",
          6519 => x"75",
          6520 => x"72",
          6521 => x"83",
          6522 => x"52",
          6523 => x"34",
          6524 => x"08",
          6525 => x"71",
          6526 => x"83",
          6527 => x"55",
          6528 => x"81",
          6529 => x"0b",
          6530 => x"e8",
          6531 => x"98",
          6532 => x"f5",
          6533 => x"80",
          6534 => x"53",
          6535 => x"9c",
          6536 => x"c0",
          6537 => x"51",
          6538 => x"f6",
          6539 => x"33",
          6540 => x"9c",
          6541 => x"74",
          6542 => x"38",
          6543 => x"2e",
          6544 => x"c0",
          6545 => x"51",
          6546 => x"73",
          6547 => x"38",
          6548 => x"ff",
          6549 => x"38",
          6550 => x"9c",
          6551 => x"90",
          6552 => x"c0",
          6553 => x"52",
          6554 => x"9c",
          6555 => x"72",
          6556 => x"81",
          6557 => x"c0",
          6558 => x"52",
          6559 => x"27",
          6560 => x"81",
          6561 => x"38",
          6562 => x"a4",
          6563 => x"75",
          6564 => x"ff",
          6565 => x"ff",
          6566 => x"ff",
          6567 => x"75",
          6568 => x"c7",
          6569 => x"ff",
          6570 => x"fe",
          6571 => x"51",
          6572 => x"06",
          6573 => x"38",
          6574 => x"7b",
          6575 => x"55",
          6576 => x"73",
          6577 => x"71",
          6578 => x"53",
          6579 => x"81",
          6580 => x"72",
          6581 => x"38",
          6582 => x"84",
          6583 => x"0d",
          6584 => x"84",
          6585 => x"88",
          6586 => x"ff",
          6587 => x"fa",
          6588 => x"02",
          6589 => x"05",
          6590 => x"80",
          6591 => x"90",
          6592 => x"2b",
          6593 => x"80",
          6594 => x"98",
          6595 => x"55",
          6596 => x"83",
          6597 => x"90",
          6598 => x"84",
          6599 => x"90",
          6600 => x"85",
          6601 => x"86",
          6602 => x"83",
          6603 => x"80",
          6604 => x"80",
          6605 => x"55",
          6606 => x"27",
          6607 => x"70",
          6608 => x"33",
          6609 => x"05",
          6610 => x"71",
          6611 => x"83",
          6612 => x"54",
          6613 => x"34",
          6614 => x"08",
          6615 => x"75",
          6616 => x"83",
          6617 => x"55",
          6618 => x"81",
          6619 => x"0b",
          6620 => x"e8",
          6621 => x"98",
          6622 => x"f5",
          6623 => x"80",
          6624 => x"53",
          6625 => x"9c",
          6626 => x"c0",
          6627 => x"51",
          6628 => x"f6",
          6629 => x"33",
          6630 => x"9c",
          6631 => x"74",
          6632 => x"38",
          6633 => x"2e",
          6634 => x"c0",
          6635 => x"51",
          6636 => x"73",
          6637 => x"38",
          6638 => x"ff",
          6639 => x"38",
          6640 => x"9c",
          6641 => x"90",
          6642 => x"c0",
          6643 => x"52",
          6644 => x"9c",
          6645 => x"72",
          6646 => x"81",
          6647 => x"c0",
          6648 => x"52",
          6649 => x"27",
          6650 => x"81",
          6651 => x"38",
          6652 => x"a4",
          6653 => x"75",
          6654 => x"ff",
          6655 => x"ff",
          6656 => x"ff",
          6657 => x"75",
          6658 => x"38",
          6659 => x"06",
          6660 => x"d5",
          6661 => x"70",
          6662 => x"54",
          6663 => x"83",
          6664 => x"76",
          6665 => x"0c",
          6666 => x"04",
          6667 => x"39",
          6668 => x"83",
          6669 => x"51",
          6670 => x"34",
          6671 => x"f5",
          6672 => x"56",
          6673 => x"16",
          6674 => x"87",
          6675 => x"34",
          6676 => x"9c",
          6677 => x"90",
          6678 => x"ce",
          6679 => x"87",
          6680 => x"08",
          6681 => x"98",
          6682 => x"72",
          6683 => x"38",
          6684 => x"87",
          6685 => x"08",
          6686 => x"74",
          6687 => x"71",
          6688 => x"db",
          6689 => x"98",
          6690 => x"ff",
          6691 => x"27",
          6692 => x"71",
          6693 => x"2e",
          6694 => x"87",
          6695 => x"08",
          6696 => x"05",
          6697 => x"98",
          6698 => x"87",
          6699 => x"08",
          6700 => x"2e",
          6701 => x"15",
          6702 => x"98",
          6703 => x"52",
          6704 => x"87",
          6705 => x"ff",
          6706 => x"87",
          6707 => x"08",
          6708 => x"26",
          6709 => x"52",
          6710 => x"16",
          6711 => x"06",
          6712 => x"80",
          6713 => x"72",
          6714 => x"54",
          6715 => x"38",
          6716 => x"3d",
          6717 => x"88",
          6718 => x"f7",
          6719 => x"0d",
          6720 => x"0d",
          6721 => x"08",
          6722 => x"83",
          6723 => x"ff",
          6724 => x"83",
          6725 => x"70",
          6726 => x"33",
          6727 => x"71",
          6728 => x"77",
          6729 => x"81",
          6730 => x"98",
          6731 => x"2b",
          6732 => x"41",
          6733 => x"57",
          6734 => x"57",
          6735 => x"24",
          6736 => x"72",
          6737 => x"33",
          6738 => x"71",
          6739 => x"83",
          6740 => x"05",
          6741 => x"12",
          6742 => x"2b",
          6743 => x"07",
          6744 => x"52",
          6745 => x"80",
          6746 => x"9e",
          6747 => x"33",
          6748 => x"71",
          6749 => x"83",
          6750 => x"05",
          6751 => x"52",
          6752 => x"74",
          6753 => x"73",
          6754 => x"54",
          6755 => x"34",
          6756 => x"08",
          6757 => x"12",
          6758 => x"33",
          6759 => x"07",
          6760 => x"5c",
          6761 => x"51",
          6762 => x"34",
          6763 => x"34",
          6764 => x"08",
          6765 => x"0b",
          6766 => x"80",
          6767 => x"34",
          6768 => x"08",
          6769 => x"14",
          6770 => x"14",
          6771 => x"f4",
          6772 => x"33",
          6773 => x"71",
          6774 => x"82",
          6775 => x"70",
          6776 => x"58",
          6777 => x"72",
          6778 => x"13",
          6779 => x"0d",
          6780 => x"33",
          6781 => x"71",
          6782 => x"83",
          6783 => x"11",
          6784 => x"85",
          6785 => x"88",
          6786 => x"88",
          6787 => x"54",
          6788 => x"58",
          6789 => x"34",
          6790 => x"34",
          6791 => x"08",
          6792 => x"11",
          6793 => x"33",
          6794 => x"71",
          6795 => x"56",
          6796 => x"72",
          6797 => x"33",
          6798 => x"71",
          6799 => x"70",
          6800 => x"55",
          6801 => x"86",
          6802 => x"87",
          6803 => x"ba",
          6804 => x"70",
          6805 => x"33",
          6806 => x"07",
          6807 => x"06",
          6808 => x"5a",
          6809 => x"76",
          6810 => x"81",
          6811 => x"ba",
          6812 => x"17",
          6813 => x"12",
          6814 => x"2b",
          6815 => x"07",
          6816 => x"33",
          6817 => x"71",
          6818 => x"70",
          6819 => x"ff",
          6820 => x"05",
          6821 => x"54",
          6822 => x"5c",
          6823 => x"52",
          6824 => x"34",
          6825 => x"34",
          6826 => x"08",
          6827 => x"33",
          6828 => x"71",
          6829 => x"83",
          6830 => x"05",
          6831 => x"12",
          6832 => x"2b",
          6833 => x"ff",
          6834 => x"2a",
          6835 => x"55",
          6836 => x"52",
          6837 => x"70",
          6838 => x"84",
          6839 => x"70",
          6840 => x"33",
          6841 => x"71",
          6842 => x"83",
          6843 => x"05",
          6844 => x"12",
          6845 => x"2b",
          6846 => x"07",
          6847 => x"52",
          6848 => x"53",
          6849 => x"fc",
          6850 => x"33",
          6851 => x"71",
          6852 => x"82",
          6853 => x"70",
          6854 => x"59",
          6855 => x"34",
          6856 => x"34",
          6857 => x"08",
          6858 => x"33",
          6859 => x"71",
          6860 => x"83",
          6861 => x"05",
          6862 => x"83",
          6863 => x"88",
          6864 => x"88",
          6865 => x"5c",
          6866 => x"52",
          6867 => x"15",
          6868 => x"15",
          6869 => x"0d",
          6870 => x"0d",
          6871 => x"f4",
          6872 => x"76",
          6873 => x"38",
          6874 => x"86",
          6875 => x"fb",
          6876 => x"3d",
          6877 => x"ff",
          6878 => x"ba",
          6879 => x"80",
          6880 => x"f0",
          6881 => x"80",
          6882 => x"84",
          6883 => x"fe",
          6884 => x"84",
          6885 => x"55",
          6886 => x"81",
          6887 => x"34",
          6888 => x"08",
          6889 => x"15",
          6890 => x"85",
          6891 => x"ba",
          6892 => x"76",
          6893 => x"81",
          6894 => x"34",
          6895 => x"08",
          6896 => x"22",
          6897 => x"80",
          6898 => x"83",
          6899 => x"70",
          6900 => x"51",
          6901 => x"88",
          6902 => x"89",
          6903 => x"ba",
          6904 => x"10",
          6905 => x"ba",
          6906 => x"f8",
          6907 => x"76",
          6908 => x"81",
          6909 => x"34",
          6910 => x"f7",
          6911 => x"52",
          6912 => x"51",
          6913 => x"8e",
          6914 => x"83",
          6915 => x"70",
          6916 => x"06",
          6917 => x"83",
          6918 => x"84",
          6919 => x"84",
          6920 => x"12",
          6921 => x"2b",
          6922 => x"59",
          6923 => x"81",
          6924 => x"75",
          6925 => x"cc",
          6926 => x"10",
          6927 => x"33",
          6928 => x"71",
          6929 => x"70",
          6930 => x"06",
          6931 => x"83",
          6932 => x"70",
          6933 => x"53",
          6934 => x"52",
          6935 => x"8a",
          6936 => x"2e",
          6937 => x"73",
          6938 => x"12",
          6939 => x"33",
          6940 => x"07",
          6941 => x"c1",
          6942 => x"ff",
          6943 => x"38",
          6944 => x"56",
          6945 => x"2b",
          6946 => x"33",
          6947 => x"71",
          6948 => x"70",
          6949 => x"06",
          6950 => x"56",
          6951 => x"79",
          6952 => x"81",
          6953 => x"74",
          6954 => x"8d",
          6955 => x"78",
          6956 => x"85",
          6957 => x"2e",
          6958 => x"74",
          6959 => x"2b",
          6960 => x"82",
          6961 => x"70",
          6962 => x"5c",
          6963 => x"76",
          6964 => x"81",
          6965 => x"ba",
          6966 => x"76",
          6967 => x"53",
          6968 => x"34",
          6969 => x"34",
          6970 => x"08",
          6971 => x"33",
          6972 => x"71",
          6973 => x"70",
          6974 => x"ff",
          6975 => x"05",
          6976 => x"ff",
          6977 => x"2a",
          6978 => x"57",
          6979 => x"75",
          6980 => x"72",
          6981 => x"53",
          6982 => x"34",
          6983 => x"08",
          6984 => x"74",
          6985 => x"15",
          6986 => x"f4",
          6987 => x"86",
          6988 => x"12",
          6989 => x"2b",
          6990 => x"07",
          6991 => x"5c",
          6992 => x"75",
          6993 => x"72",
          6994 => x"84",
          6995 => x"70",
          6996 => x"05",
          6997 => x"87",
          6998 => x"88",
          6999 => x"88",
          7000 => x"58",
          7001 => x"15",
          7002 => x"15",
          7003 => x"f4",
          7004 => x"84",
          7005 => x"12",
          7006 => x"2b",
          7007 => x"07",
          7008 => x"5a",
          7009 => x"75",
          7010 => x"72",
          7011 => x"84",
          7012 => x"70",
          7013 => x"05",
          7014 => x"85",
          7015 => x"88",
          7016 => x"88",
          7017 => x"57",
          7018 => x"15",
          7019 => x"15",
          7020 => x"f4",
          7021 => x"05",
          7022 => x"bb",
          7023 => x"3d",
          7024 => x"14",
          7025 => x"33",
          7026 => x"71",
          7027 => x"79",
          7028 => x"33",
          7029 => x"71",
          7030 => x"70",
          7031 => x"5b",
          7032 => x"52",
          7033 => x"34",
          7034 => x"34",
          7035 => x"08",
          7036 => x"11",
          7037 => x"33",
          7038 => x"71",
          7039 => x"74",
          7040 => x"33",
          7041 => x"71",
          7042 => x"70",
          7043 => x"5d",
          7044 => x"5b",
          7045 => x"86",
          7046 => x"87",
          7047 => x"ba",
          7048 => x"70",
          7049 => x"33",
          7050 => x"07",
          7051 => x"06",
          7052 => x"59",
          7053 => x"75",
          7054 => x"81",
          7055 => x"ba",
          7056 => x"84",
          7057 => x"f1",
          7058 => x"0d",
          7059 => x"f4",
          7060 => x"76",
          7061 => x"38",
          7062 => x"8a",
          7063 => x"bb",
          7064 => x"3d",
          7065 => x"51",
          7066 => x"84",
          7067 => x"84",
          7068 => x"89",
          7069 => x"84",
          7070 => x"84",
          7071 => x"a0",
          7072 => x"ba",
          7073 => x"80",
          7074 => x"52",
          7075 => x"51",
          7076 => x"3f",
          7077 => x"08",
          7078 => x"34",
          7079 => x"16",
          7080 => x"f4",
          7081 => x"84",
          7082 => x"0b",
          7083 => x"84",
          7084 => x"56",
          7085 => x"34",
          7086 => x"17",
          7087 => x"f4",
          7088 => x"f0",
          7089 => x"fe",
          7090 => x"70",
          7091 => x"06",
          7092 => x"58",
          7093 => x"74",
          7094 => x"73",
          7095 => x"84",
          7096 => x"70",
          7097 => x"84",
          7098 => x"05",
          7099 => x"55",
          7100 => x"34",
          7101 => x"15",
          7102 => x"77",
          7103 => x"dd",
          7104 => x"39",
          7105 => x"65",
          7106 => x"80",
          7107 => x"f4",
          7108 => x"41",
          7109 => x"84",
          7110 => x"80",
          7111 => x"38",
          7112 => x"88",
          7113 => x"54",
          7114 => x"8f",
          7115 => x"05",
          7116 => x"05",
          7117 => x"ff",
          7118 => x"73",
          7119 => x"06",
          7120 => x"83",
          7121 => x"ff",
          7122 => x"83",
          7123 => x"70",
          7124 => x"33",
          7125 => x"07",
          7126 => x"70",
          7127 => x"06",
          7128 => x"10",
          7129 => x"83",
          7130 => x"70",
          7131 => x"33",
          7132 => x"07",
          7133 => x"70",
          7134 => x"42",
          7135 => x"53",
          7136 => x"5c",
          7137 => x"5e",
          7138 => x"7a",
          7139 => x"38",
          7140 => x"83",
          7141 => x"88",
          7142 => x"10",
          7143 => x"70",
          7144 => x"33",
          7145 => x"71",
          7146 => x"53",
          7147 => x"56",
          7148 => x"24",
          7149 => x"7a",
          7150 => x"f6",
          7151 => x"58",
          7152 => x"87",
          7153 => x"80",
          7154 => x"38",
          7155 => x"77",
          7156 => x"be",
          7157 => x"59",
          7158 => x"92",
          7159 => x"1e",
          7160 => x"12",
          7161 => x"2b",
          7162 => x"07",
          7163 => x"33",
          7164 => x"71",
          7165 => x"90",
          7166 => x"43",
          7167 => x"57",
          7168 => x"60",
          7169 => x"38",
          7170 => x"11",
          7171 => x"33",
          7172 => x"71",
          7173 => x"7a",
          7174 => x"33",
          7175 => x"71",
          7176 => x"83",
          7177 => x"05",
          7178 => x"85",
          7179 => x"88",
          7180 => x"88",
          7181 => x"48",
          7182 => x"58",
          7183 => x"56",
          7184 => x"34",
          7185 => x"34",
          7186 => x"08",
          7187 => x"11",
          7188 => x"33",
          7189 => x"71",
          7190 => x"74",
          7191 => x"33",
          7192 => x"71",
          7193 => x"70",
          7194 => x"42",
          7195 => x"57",
          7196 => x"86",
          7197 => x"87",
          7198 => x"ba",
          7199 => x"70",
          7200 => x"33",
          7201 => x"07",
          7202 => x"06",
          7203 => x"5a",
          7204 => x"76",
          7205 => x"81",
          7206 => x"ba",
          7207 => x"1f",
          7208 => x"83",
          7209 => x"8b",
          7210 => x"2b",
          7211 => x"73",
          7212 => x"33",
          7213 => x"07",
          7214 => x"41",
          7215 => x"5f",
          7216 => x"79",
          7217 => x"81",
          7218 => x"ba",
          7219 => x"1f",
          7220 => x"12",
          7221 => x"2b",
          7222 => x"07",
          7223 => x"14",
          7224 => x"33",
          7225 => x"07",
          7226 => x"41",
          7227 => x"5f",
          7228 => x"79",
          7229 => x"75",
          7230 => x"84",
          7231 => x"70",
          7232 => x"33",
          7233 => x"71",
          7234 => x"66",
          7235 => x"70",
          7236 => x"52",
          7237 => x"05",
          7238 => x"fe",
          7239 => x"84",
          7240 => x"1e",
          7241 => x"65",
          7242 => x"83",
          7243 => x"5d",
          7244 => x"62",
          7245 => x"38",
          7246 => x"84",
          7247 => x"95",
          7248 => x"84",
          7249 => x"84",
          7250 => x"a0",
          7251 => x"ba",
          7252 => x"80",
          7253 => x"52",
          7254 => x"51",
          7255 => x"3f",
          7256 => x"08",
          7257 => x"34",
          7258 => x"1f",
          7259 => x"f4",
          7260 => x"84",
          7261 => x"0b",
          7262 => x"84",
          7263 => x"5c",
          7264 => x"34",
          7265 => x"1d",
          7266 => x"f4",
          7267 => x"f0",
          7268 => x"fe",
          7269 => x"70",
          7270 => x"06",
          7271 => x"5c",
          7272 => x"78",
          7273 => x"77",
          7274 => x"84",
          7275 => x"70",
          7276 => x"84",
          7277 => x"05",
          7278 => x"56",
          7279 => x"34",
          7280 => x"15",
          7281 => x"f4",
          7282 => x"fa",
          7283 => x"80",
          7284 => x"38",
          7285 => x"80",
          7286 => x"38",
          7287 => x"9b",
          7288 => x"84",
          7289 => x"84",
          7290 => x"0d",
          7291 => x"84",
          7292 => x"71",
          7293 => x"11",
          7294 => x"05",
          7295 => x"12",
          7296 => x"2b",
          7297 => x"ff",
          7298 => x"2a",
          7299 => x"5e",
          7300 => x"34",
          7301 => x"34",
          7302 => x"f4",
          7303 => x"88",
          7304 => x"75",
          7305 => x"7b",
          7306 => x"84",
          7307 => x"70",
          7308 => x"81",
          7309 => x"88",
          7310 => x"83",
          7311 => x"f8",
          7312 => x"64",
          7313 => x"06",
          7314 => x"4a",
          7315 => x"5e",
          7316 => x"63",
          7317 => x"76",
          7318 => x"41",
          7319 => x"05",
          7320 => x"f4",
          7321 => x"63",
          7322 => x"81",
          7323 => x"84",
          7324 => x"05",
          7325 => x"ed",
          7326 => x"54",
          7327 => x"7b",
          7328 => x"83",
          7329 => x"42",
          7330 => x"39",
          7331 => x"ff",
          7332 => x"70",
          7333 => x"06",
          7334 => x"83",
          7335 => x"88",
          7336 => x"10",
          7337 => x"70",
          7338 => x"33",
          7339 => x"71",
          7340 => x"53",
          7341 => x"58",
          7342 => x"73",
          7343 => x"f7",
          7344 => x"39",
          7345 => x"fa",
          7346 => x"7a",
          7347 => x"38",
          7348 => x"ff",
          7349 => x"7b",
          7350 => x"38",
          7351 => x"84",
          7352 => x"84",
          7353 => x"a0",
          7354 => x"ba",
          7355 => x"80",
          7356 => x"52",
          7357 => x"51",
          7358 => x"3f",
          7359 => x"08",
          7360 => x"34",
          7361 => x"1b",
          7362 => x"f4",
          7363 => x"84",
          7364 => x"0b",
          7365 => x"84",
          7366 => x"58",
          7367 => x"34",
          7368 => x"19",
          7369 => x"f4",
          7370 => x"f0",
          7371 => x"fe",
          7372 => x"70",
          7373 => x"06",
          7374 => x"58",
          7375 => x"74",
          7376 => x"34",
          7377 => x"05",
          7378 => x"f0",
          7379 => x"10",
          7380 => x"f4",
          7381 => x"05",
          7382 => x"61",
          7383 => x"81",
          7384 => x"34",
          7385 => x"80",
          7386 => x"de",
          7387 => x"ff",
          7388 => x"61",
          7389 => x"c0",
          7390 => x"39",
          7391 => x"82",
          7392 => x"51",
          7393 => x"7f",
          7394 => x"bb",
          7395 => x"3d",
          7396 => x"1e",
          7397 => x"83",
          7398 => x"8b",
          7399 => x"2b",
          7400 => x"86",
          7401 => x"12",
          7402 => x"2b",
          7403 => x"07",
          7404 => x"14",
          7405 => x"33",
          7406 => x"07",
          7407 => x"43",
          7408 => x"5b",
          7409 => x"5c",
          7410 => x"64",
          7411 => x"7a",
          7412 => x"34",
          7413 => x"08",
          7414 => x"11",
          7415 => x"33",
          7416 => x"71",
          7417 => x"74",
          7418 => x"33",
          7419 => x"71",
          7420 => x"70",
          7421 => x"41",
          7422 => x"59",
          7423 => x"64",
          7424 => x"7a",
          7425 => x"34",
          7426 => x"08",
          7427 => x"81",
          7428 => x"88",
          7429 => x"ff",
          7430 => x"88",
          7431 => x"5a",
          7432 => x"34",
          7433 => x"34",
          7434 => x"08",
          7435 => x"11",
          7436 => x"33",
          7437 => x"71",
          7438 => x"74",
          7439 => x"81",
          7440 => x"88",
          7441 => x"88",
          7442 => x"5e",
          7443 => x"45",
          7444 => x"34",
          7445 => x"34",
          7446 => x"08",
          7447 => x"33",
          7448 => x"71",
          7449 => x"83",
          7450 => x"05",
          7451 => x"83",
          7452 => x"88",
          7453 => x"88",
          7454 => x"40",
          7455 => x"55",
          7456 => x"18",
          7457 => x"18",
          7458 => x"f4",
          7459 => x"82",
          7460 => x"12",
          7461 => x"2b",
          7462 => x"62",
          7463 => x"2b",
          7464 => x"5d",
          7465 => x"05",
          7466 => x"96",
          7467 => x"f4",
          7468 => x"05",
          7469 => x"ff",
          7470 => x"fc",
          7471 => x"ff",
          7472 => x"ba",
          7473 => x"80",
          7474 => x"f0",
          7475 => x"80",
          7476 => x"84",
          7477 => x"fe",
          7478 => x"84",
          7479 => x"56",
          7480 => x"81",
          7481 => x"34",
          7482 => x"08",
          7483 => x"16",
          7484 => x"85",
          7485 => x"ba",
          7486 => x"7f",
          7487 => x"81",
          7488 => x"34",
          7489 => x"08",
          7490 => x"22",
          7491 => x"80",
          7492 => x"83",
          7493 => x"70",
          7494 => x"43",
          7495 => x"88",
          7496 => x"89",
          7497 => x"ba",
          7498 => x"10",
          7499 => x"ba",
          7500 => x"f8",
          7501 => x"7f",
          7502 => x"81",
          7503 => x"34",
          7504 => x"bd",
          7505 => x"fc",
          7506 => x"19",
          7507 => x"33",
          7508 => x"71",
          7509 => x"79",
          7510 => x"33",
          7511 => x"71",
          7512 => x"70",
          7513 => x"48",
          7514 => x"55",
          7515 => x"05",
          7516 => x"85",
          7517 => x"ba",
          7518 => x"1e",
          7519 => x"85",
          7520 => x"8b",
          7521 => x"2b",
          7522 => x"86",
          7523 => x"15",
          7524 => x"2b",
          7525 => x"2a",
          7526 => x"48",
          7527 => x"40",
          7528 => x"05",
          7529 => x"87",
          7530 => x"ba",
          7531 => x"70",
          7532 => x"33",
          7533 => x"07",
          7534 => x"06",
          7535 => x"59",
          7536 => x"75",
          7537 => x"81",
          7538 => x"ba",
          7539 => x"1f",
          7540 => x"12",
          7541 => x"2b",
          7542 => x"07",
          7543 => x"33",
          7544 => x"71",
          7545 => x"70",
          7546 => x"ff",
          7547 => x"05",
          7548 => x"48",
          7549 => x"5d",
          7550 => x"41",
          7551 => x"34",
          7552 => x"34",
          7553 => x"08",
          7554 => x"33",
          7555 => x"71",
          7556 => x"83",
          7557 => x"05",
          7558 => x"12",
          7559 => x"2b",
          7560 => x"ff",
          7561 => x"2a",
          7562 => x"5e",
          7563 => x"5b",
          7564 => x"76",
          7565 => x"34",
          7566 => x"ff",
          7567 => x"b3",
          7568 => x"33",
          7569 => x"71",
          7570 => x"83",
          7571 => x"05",
          7572 => x"85",
          7573 => x"88",
          7574 => x"88",
          7575 => x"5a",
          7576 => x"78",
          7577 => x"79",
          7578 => x"84",
          7579 => x"70",
          7580 => x"33",
          7581 => x"71",
          7582 => x"83",
          7583 => x"05",
          7584 => x"87",
          7585 => x"88",
          7586 => x"88",
          7587 => x"5e",
          7588 => x"55",
          7589 => x"86",
          7590 => x"60",
          7591 => x"84",
          7592 => x"18",
          7593 => x"12",
          7594 => x"2b",
          7595 => x"ff",
          7596 => x"2a",
          7597 => x"55",
          7598 => x"78",
          7599 => x"84",
          7600 => x"70",
          7601 => x"81",
          7602 => x"8b",
          7603 => x"2b",
          7604 => x"70",
          7605 => x"33",
          7606 => x"07",
          7607 => x"8f",
          7608 => x"77",
          7609 => x"2a",
          7610 => x"5f",
          7611 => x"5e",
          7612 => x"17",
          7613 => x"17",
          7614 => x"f4",
          7615 => x"70",
          7616 => x"33",
          7617 => x"71",
          7618 => x"74",
          7619 => x"81",
          7620 => x"88",
          7621 => x"ff",
          7622 => x"88",
          7623 => x"5e",
          7624 => x"5d",
          7625 => x"34",
          7626 => x"34",
          7627 => x"08",
          7628 => x"11",
          7629 => x"33",
          7630 => x"71",
          7631 => x"74",
          7632 => x"33",
          7633 => x"71",
          7634 => x"83",
          7635 => x"05",
          7636 => x"85",
          7637 => x"88",
          7638 => x"88",
          7639 => x"49",
          7640 => x"59",
          7641 => x"57",
          7642 => x"1d",
          7643 => x"1d",
          7644 => x"f4",
          7645 => x"84",
          7646 => x"12",
          7647 => x"2b",
          7648 => x"07",
          7649 => x"14",
          7650 => x"33",
          7651 => x"07",
          7652 => x"5f",
          7653 => x"40",
          7654 => x"77",
          7655 => x"7b",
          7656 => x"84",
          7657 => x"16",
          7658 => x"12",
          7659 => x"2b",
          7660 => x"ff",
          7661 => x"2a",
          7662 => x"59",
          7663 => x"79",
          7664 => x"84",
          7665 => x"70",
          7666 => x"33",
          7667 => x"71",
          7668 => x"83",
          7669 => x"05",
          7670 => x"15",
          7671 => x"2b",
          7672 => x"2a",
          7673 => x"5d",
          7674 => x"55",
          7675 => x"75",
          7676 => x"84",
          7677 => x"70",
          7678 => x"81",
          7679 => x"8b",
          7680 => x"2b",
          7681 => x"82",
          7682 => x"15",
          7683 => x"2b",
          7684 => x"2a",
          7685 => x"5d",
          7686 => x"55",
          7687 => x"34",
          7688 => x"34",
          7689 => x"08",
          7690 => x"11",
          7691 => x"33",
          7692 => x"07",
          7693 => x"56",
          7694 => x"42",
          7695 => x"7e",
          7696 => x"51",
          7697 => x"3f",
          7698 => x"08",
          7699 => x"61",
          7700 => x"70",
          7701 => x"06",
          7702 => x"f1",
          7703 => x"19",
          7704 => x"33",
          7705 => x"71",
          7706 => x"79",
          7707 => x"33",
          7708 => x"71",
          7709 => x"70",
          7710 => x"48",
          7711 => x"55",
          7712 => x"05",
          7713 => x"85",
          7714 => x"ba",
          7715 => x"1e",
          7716 => x"85",
          7717 => x"8b",
          7718 => x"2b",
          7719 => x"86",
          7720 => x"15",
          7721 => x"2b",
          7722 => x"2a",
          7723 => x"48",
          7724 => x"56",
          7725 => x"05",
          7726 => x"87",
          7727 => x"ba",
          7728 => x"70",
          7729 => x"33",
          7730 => x"07",
          7731 => x"06",
          7732 => x"5c",
          7733 => x"78",
          7734 => x"81",
          7735 => x"ba",
          7736 => x"1f",
          7737 => x"12",
          7738 => x"2b",
          7739 => x"07",
          7740 => x"33",
          7741 => x"71",
          7742 => x"70",
          7743 => x"ff",
          7744 => x"05",
          7745 => x"5d",
          7746 => x"58",
          7747 => x"40",
          7748 => x"34",
          7749 => x"34",
          7750 => x"08",
          7751 => x"33",
          7752 => x"71",
          7753 => x"83",
          7754 => x"05",
          7755 => x"12",
          7756 => x"2b",
          7757 => x"ff",
          7758 => x"2a",
          7759 => x"58",
          7760 => x"5b",
          7761 => x"78",
          7762 => x"77",
          7763 => x"06",
          7764 => x"39",
          7765 => x"54",
          7766 => x"84",
          7767 => x"5f",
          7768 => x"08",
          7769 => x"38",
          7770 => x"52",
          7771 => x"08",
          7772 => x"f6",
          7773 => x"df",
          7774 => x"5b",
          7775 => x"ef",
          7776 => x"e9",
          7777 => x"0d",
          7778 => x"84",
          7779 => x"58",
          7780 => x"2e",
          7781 => x"54",
          7782 => x"73",
          7783 => x"0c",
          7784 => x"04",
          7785 => x"d3",
          7786 => x"84",
          7787 => x"bb",
          7788 => x"2e",
          7789 => x"53",
          7790 => x"bb",
          7791 => x"fe",
          7792 => x"73",
          7793 => x"0c",
          7794 => x"04",
          7795 => x"0b",
          7796 => x"0c",
          7797 => x"84",
          7798 => x"82",
          7799 => x"76",
          7800 => x"f4",
          7801 => x"97",
          7802 => x"f4",
          7803 => x"75",
          7804 => x"81",
          7805 => x"ba",
          7806 => x"76",
          7807 => x"81",
          7808 => x"34",
          7809 => x"08",
          7810 => x"17",
          7811 => x"87",
          7812 => x"ba",
          7813 => x"ba",
          7814 => x"05",
          7815 => x"07",
          7816 => x"ff",
          7817 => x"2a",
          7818 => x"56",
          7819 => x"34",
          7820 => x"34",
          7821 => x"22",
          7822 => x"10",
          7823 => x"08",
          7824 => x"55",
          7825 => x"15",
          7826 => x"83",
          7827 => x"54",
          7828 => x"fe",
          7829 => x"cc",
          7830 => x"0d",
          7831 => x"33",
          7832 => x"70",
          7833 => x"38",
          7834 => x"11",
          7835 => x"84",
          7836 => x"83",
          7837 => x"fe",
          7838 => x"93",
          7839 => x"83",
          7840 => x"26",
          7841 => x"51",
          7842 => x"84",
          7843 => x"81",
          7844 => x"72",
          7845 => x"84",
          7846 => x"34",
          7847 => x"12",
          7848 => x"84",
          7849 => x"84",
          7850 => x"f7",
          7851 => x"7e",
          7852 => x"05",
          7853 => x"5a",
          7854 => x"81",
          7855 => x"26",
          7856 => x"bb",
          7857 => x"54",
          7858 => x"54",
          7859 => x"bd",
          7860 => x"85",
          7861 => x"98",
          7862 => x"53",
          7863 => x"51",
          7864 => x"84",
          7865 => x"81",
          7866 => x"74",
          7867 => x"38",
          7868 => x"8c",
          7869 => x"e2",
          7870 => x"26",
          7871 => x"fc",
          7872 => x"54",
          7873 => x"83",
          7874 => x"73",
          7875 => x"bb",
          7876 => x"3d",
          7877 => x"80",
          7878 => x"70",
          7879 => x"5a",
          7880 => x"78",
          7881 => x"38",
          7882 => x"3d",
          7883 => x"60",
          7884 => x"af",
          7885 => x"5c",
          7886 => x"54",
          7887 => x"87",
          7888 => x"80",
          7889 => x"73",
          7890 => x"83",
          7891 => x"38",
          7892 => x"0b",
          7893 => x"8c",
          7894 => x"75",
          7895 => x"d7",
          7896 => x"bb",
          7897 => x"ff",
          7898 => x"80",
          7899 => x"87",
          7900 => x"08",
          7901 => x"38",
          7902 => x"d6",
          7903 => x"80",
          7904 => x"73",
          7905 => x"38",
          7906 => x"55",
          7907 => x"84",
          7908 => x"0d",
          7909 => x"16",
          7910 => x"81",
          7911 => x"55",
          7912 => x"26",
          7913 => x"d5",
          7914 => x"0d",
          7915 => x"05",
          7916 => x"02",
          7917 => x"05",
          7918 => x"55",
          7919 => x"73",
          7920 => x"84",
          7921 => x"33",
          7922 => x"06",
          7923 => x"73",
          7924 => x"0b",
          7925 => x"8c",
          7926 => x"70",
          7927 => x"38",
          7928 => x"ad",
          7929 => x"2e",
          7930 => x"53",
          7931 => x"84",
          7932 => x"0d",
          7933 => x"0a",
          7934 => x"84",
          7935 => x"86",
          7936 => x"81",
          7937 => x"80",
          7938 => x"84",
          7939 => x"0d",
          7940 => x"2b",
          7941 => x"8c",
          7942 => x"70",
          7943 => x"08",
          7944 => x"81",
          7945 => x"70",
          7946 => x"38",
          7947 => x"8c",
          7948 => x"ea",
          7949 => x"98",
          7950 => x"70",
          7951 => x"72",
          7952 => x"92",
          7953 => x"71",
          7954 => x"54",
          7955 => x"ff",
          7956 => x"08",
          7957 => x"73",
          7958 => x"90",
          7959 => x"0d",
          7960 => x"0b",
          7961 => x"71",
          7962 => x"74",
          7963 => x"81",
          7964 => x"77",
          7965 => x"83",
          7966 => x"38",
          7967 => x"52",
          7968 => x"51",
          7969 => x"84",
          7970 => x"80",
          7971 => x"81",
          7972 => x"bb",
          7973 => x"3d",
          7974 => x"54",
          7975 => x"53",
          7976 => x"53",
          7977 => x"52",
          7978 => x"3f",
          7979 => x"bb",
          7980 => x"2e",
          7981 => x"d9",
          7982 => x"84",
          7983 => x"34",
          7984 => x"70",
          7985 => x"31",
          7986 => x"84",
          7987 => x"5c",
          7988 => x"74",
          7989 => x"9b",
          7990 => x"33",
          7991 => x"2e",
          7992 => x"ff",
          7993 => x"54",
          7994 => x"79",
          7995 => x"33",
          7996 => x"3f",
          7997 => x"57",
          7998 => x"2e",
          7999 => x"fe",
          8000 => x"18",
          8001 => x"81",
          8002 => x"06",
          8003 => x"b8",
          8004 => x"80",
          8005 => x"80",
          8006 => x"05",
          8007 => x"17",
          8008 => x"38",
          8009 => x"84",
          8010 => x"ff",
          8011 => x"b7",
          8012 => x"d2",
          8013 => x"d2",
          8014 => x"34",
          8015 => x"ba",
          8016 => x"c1",
          8017 => x"34",
          8018 => x"84",
          8019 => x"80",
          8020 => x"9d",
          8021 => x"c1",
          8022 => x"19",
          8023 => x"0b",
          8024 => x"34",
          8025 => x"55",
          8026 => x"19",
          8027 => x"2a",
          8028 => x"a1",
          8029 => x"90",
          8030 => x"84",
          8031 => x"74",
          8032 => x"7a",
          8033 => x"34",
          8034 => x"5b",
          8035 => x"19",
          8036 => x"2a",
          8037 => x"a5",
          8038 => x"90",
          8039 => x"84",
          8040 => x"7a",
          8041 => x"74",
          8042 => x"34",
          8043 => x"81",
          8044 => x"1a",
          8045 => x"54",
          8046 => x"52",
          8047 => x"51",
          8048 => x"76",
          8049 => x"80",
          8050 => x"81",
          8051 => x"fb",
          8052 => x"bb",
          8053 => x"2e",
          8054 => x"fd",
          8055 => x"3d",
          8056 => x"70",
          8057 => x"56",
          8058 => x"88",
          8059 => x"08",
          8060 => x"38",
          8061 => x"84",
          8062 => x"8f",
          8063 => x"ff",
          8064 => x"58",
          8065 => x"81",
          8066 => x"82",
          8067 => x"38",
          8068 => x"09",
          8069 => x"38",
          8070 => x"16",
          8071 => x"a8",
          8072 => x"5a",
          8073 => x"b4",
          8074 => x"2e",
          8075 => x"17",
          8076 => x"7b",
          8077 => x"06",
          8078 => x"81",
          8079 => x"b8",
          8080 => x"17",
          8081 => x"e3",
          8082 => x"84",
          8083 => x"85",
          8084 => x"81",
          8085 => x"18",
          8086 => x"9a",
          8087 => x"ff",
          8088 => x"11",
          8089 => x"70",
          8090 => x"1b",
          8091 => x"5d",
          8092 => x"17",
          8093 => x"b5",
          8094 => x"83",
          8095 => x"5c",
          8096 => x"7d",
          8097 => x"06",
          8098 => x"81",
          8099 => x"b8",
          8100 => x"17",
          8101 => x"93",
          8102 => x"84",
          8103 => x"85",
          8104 => x"81",
          8105 => x"18",
          8106 => x"ca",
          8107 => x"ff",
          8108 => x"11",
          8109 => x"2b",
          8110 => x"81",
          8111 => x"2a",
          8112 => x"59",
          8113 => x"ae",
          8114 => x"ff",
          8115 => x"84",
          8116 => x"0d",
          8117 => x"2a",
          8118 => x"05",
          8119 => x"08",
          8120 => x"38",
          8121 => x"18",
          8122 => x"5d",
          8123 => x"2e",
          8124 => x"81",
          8125 => x"54",
          8126 => x"17",
          8127 => x"33",
          8128 => x"3f",
          8129 => x"08",
          8130 => x"38",
          8131 => x"5a",
          8132 => x"0c",
          8133 => x"38",
          8134 => x"fe",
          8135 => x"b8",
          8136 => x"33",
          8137 => x"88",
          8138 => x"bb",
          8139 => x"5b",
          8140 => x"04",
          8141 => x"09",
          8142 => x"b8",
          8143 => x"2a",
          8144 => x"05",
          8145 => x"08",
          8146 => x"38",
          8147 => x"18",
          8148 => x"5e",
          8149 => x"2e",
          8150 => x"82",
          8151 => x"54",
          8152 => x"17",
          8153 => x"33",
          8154 => x"3f",
          8155 => x"08",
          8156 => x"38",
          8157 => x"5a",
          8158 => x"0c",
          8159 => x"38",
          8160 => x"83",
          8161 => x"05",
          8162 => x"11",
          8163 => x"33",
          8164 => x"71",
          8165 => x"81",
          8166 => x"72",
          8167 => x"75",
          8168 => x"ff",
          8169 => x"06",
          8170 => x"84",
          8171 => x"5e",
          8172 => x"8f",
          8173 => x"81",
          8174 => x"08",
          8175 => x"70",
          8176 => x"33",
          8177 => x"e2",
          8178 => x"84",
          8179 => x"7b",
          8180 => x"06",
          8181 => x"84",
          8182 => x"83",
          8183 => x"17",
          8184 => x"08",
          8185 => x"84",
          8186 => x"7d",
          8187 => x"27",
          8188 => x"82",
          8189 => x"74",
          8190 => x"81",
          8191 => x"38",
          8192 => x"17",
          8193 => x"08",
          8194 => x"52",
          8195 => x"51",
          8196 => x"7a",
          8197 => x"39",
          8198 => x"17",
          8199 => x"17",
          8200 => x"18",
          8201 => x"f6",
          8202 => x"bb",
          8203 => x"2e",
          8204 => x"82",
          8205 => x"bb",
          8206 => x"18",
          8207 => x"08",
          8208 => x"31",
          8209 => x"18",
          8210 => x"38",
          8211 => x"5e",
          8212 => x"81",
          8213 => x"bb",
          8214 => x"fb",
          8215 => x"54",
          8216 => x"53",
          8217 => x"53",
          8218 => x"52",
          8219 => x"3f",
          8220 => x"bb",
          8221 => x"2e",
          8222 => x"fd",
          8223 => x"bb",
          8224 => x"18",
          8225 => x"08",
          8226 => x"31",
          8227 => x"08",
          8228 => x"a0",
          8229 => x"fd",
          8230 => x"17",
          8231 => x"82",
          8232 => x"06",
          8233 => x"81",
          8234 => x"08",
          8235 => x"05",
          8236 => x"81",
          8237 => x"f4",
          8238 => x"5a",
          8239 => x"81",
          8240 => x"08",
          8241 => x"70",
          8242 => x"33",
          8243 => x"da",
          8244 => x"84",
          8245 => x"7d",
          8246 => x"06",
          8247 => x"84",
          8248 => x"83",
          8249 => x"17",
          8250 => x"08",
          8251 => x"84",
          8252 => x"74",
          8253 => x"27",
          8254 => x"82",
          8255 => x"74",
          8256 => x"81",
          8257 => x"38",
          8258 => x"17",
          8259 => x"08",
          8260 => x"52",
          8261 => x"51",
          8262 => x"7c",
          8263 => x"39",
          8264 => x"17",
          8265 => x"08",
          8266 => x"52",
          8267 => x"51",
          8268 => x"fa",
          8269 => x"5b",
          8270 => x"38",
          8271 => x"f2",
          8272 => x"62",
          8273 => x"59",
          8274 => x"76",
          8275 => x"75",
          8276 => x"27",
          8277 => x"33",
          8278 => x"2e",
          8279 => x"78",
          8280 => x"38",
          8281 => x"82",
          8282 => x"84",
          8283 => x"90",
          8284 => x"75",
          8285 => x"1a",
          8286 => x"80",
          8287 => x"08",
          8288 => x"78",
          8289 => x"38",
          8290 => x"7c",
          8291 => x"7c",
          8292 => x"06",
          8293 => x"81",
          8294 => x"b8",
          8295 => x"19",
          8296 => x"87",
          8297 => x"84",
          8298 => x"85",
          8299 => x"81",
          8300 => x"1a",
          8301 => x"79",
          8302 => x"75",
          8303 => x"06",
          8304 => x"83",
          8305 => x"58",
          8306 => x"1f",
          8307 => x"2a",
          8308 => x"1f",
          8309 => x"83",
          8310 => x"84",
          8311 => x"90",
          8312 => x"74",
          8313 => x"81",
          8314 => x"38",
          8315 => x"a8",
          8316 => x"58",
          8317 => x"1a",
          8318 => x"76",
          8319 => x"e1",
          8320 => x"33",
          8321 => x"7c",
          8322 => x"81",
          8323 => x"38",
          8324 => x"53",
          8325 => x"81",
          8326 => x"f1",
          8327 => x"bb",
          8328 => x"2e",
          8329 => x"58",
          8330 => x"b4",
          8331 => x"58",
          8332 => x"38",
          8333 => x"83",
          8334 => x"05",
          8335 => x"11",
          8336 => x"2b",
          8337 => x"7e",
          8338 => x"07",
          8339 => x"5c",
          8340 => x"7d",
          8341 => x"75",
          8342 => x"7d",
          8343 => x"79",
          8344 => x"7d",
          8345 => x"7a",
          8346 => x"81",
          8347 => x"34",
          8348 => x"75",
          8349 => x"70",
          8350 => x"1b",
          8351 => x"1b",
          8352 => x"5a",
          8353 => x"b7",
          8354 => x"83",
          8355 => x"5e",
          8356 => x"7d",
          8357 => x"06",
          8358 => x"81",
          8359 => x"b8",
          8360 => x"19",
          8361 => x"83",
          8362 => x"84",
          8363 => x"85",
          8364 => x"81",
          8365 => x"1a",
          8366 => x"7b",
          8367 => x"79",
          8368 => x"19",
          8369 => x"1b",
          8370 => x"5f",
          8371 => x"55",
          8372 => x"8f",
          8373 => x"2b",
          8374 => x"77",
          8375 => x"71",
          8376 => x"74",
          8377 => x"0b",
          8378 => x"7d",
          8379 => x"1a",
          8380 => x"80",
          8381 => x"08",
          8382 => x"76",
          8383 => x"38",
          8384 => x"53",
          8385 => x"53",
          8386 => x"52",
          8387 => x"3f",
          8388 => x"bb",
          8389 => x"2e",
          8390 => x"80",
          8391 => x"bb",
          8392 => x"1a",
          8393 => x"08",
          8394 => x"08",
          8395 => x"08",
          8396 => x"08",
          8397 => x"5c",
          8398 => x"8b",
          8399 => x"33",
          8400 => x"2e",
          8401 => x"81",
          8402 => x"76",
          8403 => x"33",
          8404 => x"3f",
          8405 => x"08",
          8406 => x"38",
          8407 => x"58",
          8408 => x"0c",
          8409 => x"38",
          8410 => x"06",
          8411 => x"7b",
          8412 => x"56",
          8413 => x"7a",
          8414 => x"33",
          8415 => x"71",
          8416 => x"56",
          8417 => x"34",
          8418 => x"1a",
          8419 => x"39",
          8420 => x"53",
          8421 => x"53",
          8422 => x"52",
          8423 => x"3f",
          8424 => x"bb",
          8425 => x"2e",
          8426 => x"fc",
          8427 => x"bb",
          8428 => x"1a",
          8429 => x"08",
          8430 => x"08",
          8431 => x"08",
          8432 => x"08",
          8433 => x"5e",
          8434 => x"fb",
          8435 => x"19",
          8436 => x"82",
          8437 => x"06",
          8438 => x"81",
          8439 => x"53",
          8440 => x"19",
          8441 => x"c2",
          8442 => x"fb",
          8443 => x"54",
          8444 => x"19",
          8445 => x"1a",
          8446 => x"ee",
          8447 => x"5c",
          8448 => x"08",
          8449 => x"81",
          8450 => x"38",
          8451 => x"08",
          8452 => x"b4",
          8453 => x"a8",
          8454 => x"a0",
          8455 => x"bb",
          8456 => x"40",
          8457 => x"7e",
          8458 => x"38",
          8459 => x"55",
          8460 => x"09",
          8461 => x"e3",
          8462 => x"7d",
          8463 => x"52",
          8464 => x"51",
          8465 => x"7c",
          8466 => x"39",
          8467 => x"53",
          8468 => x"53",
          8469 => x"52",
          8470 => x"3f",
          8471 => x"bb",
          8472 => x"2e",
          8473 => x"fb",
          8474 => x"bb",
          8475 => x"1a",
          8476 => x"08",
          8477 => x"08",
          8478 => x"08",
          8479 => x"08",
          8480 => x"5e",
          8481 => x"fb",
          8482 => x"19",
          8483 => x"82",
          8484 => x"06",
          8485 => x"81",
          8486 => x"53",
          8487 => x"19",
          8488 => x"86",
          8489 => x"fa",
          8490 => x"54",
          8491 => x"76",
          8492 => x"33",
          8493 => x"3f",
          8494 => x"8b",
          8495 => x"10",
          8496 => x"7a",
          8497 => x"ff",
          8498 => x"5f",
          8499 => x"1f",
          8500 => x"2a",
          8501 => x"1f",
          8502 => x"39",
          8503 => x"88",
          8504 => x"82",
          8505 => x"06",
          8506 => x"11",
          8507 => x"70",
          8508 => x"0a",
          8509 => x"0a",
          8510 => x"58",
          8511 => x"7d",
          8512 => x"88",
          8513 => x"b9",
          8514 => x"90",
          8515 => x"ba",
          8516 => x"98",
          8517 => x"bb",
          8518 => x"cf",
          8519 => x"0d",
          8520 => x"08",
          8521 => x"7a",
          8522 => x"90",
          8523 => x"76",
          8524 => x"f4",
          8525 => x"1a",
          8526 => x"ec",
          8527 => x"08",
          8528 => x"73",
          8529 => x"d7",
          8530 => x"2e",
          8531 => x"76",
          8532 => x"56",
          8533 => x"76",
          8534 => x"82",
          8535 => x"26",
          8536 => x"75",
          8537 => x"f0",
          8538 => x"bb",
          8539 => x"2e",
          8540 => x"80",
          8541 => x"84",
          8542 => x"b1",
          8543 => x"84",
          8544 => x"30",
          8545 => x"80",
          8546 => x"07",
          8547 => x"55",
          8548 => x"38",
          8549 => x"09",
          8550 => x"b5",
          8551 => x"74",
          8552 => x"0c",
          8553 => x"04",
          8554 => x"91",
          8555 => x"84",
          8556 => x"39",
          8557 => x"51",
          8558 => x"81",
          8559 => x"bb",
          8560 => x"db",
          8561 => x"84",
          8562 => x"bb",
          8563 => x"2e",
          8564 => x"19",
          8565 => x"84",
          8566 => x"38",
          8567 => x"dd",
          8568 => x"56",
          8569 => x"76",
          8570 => x"82",
          8571 => x"79",
          8572 => x"3f",
          8573 => x"bb",
          8574 => x"2e",
          8575 => x"84",
          8576 => x"09",
          8577 => x"72",
          8578 => x"70",
          8579 => x"bb",
          8580 => x"51",
          8581 => x"73",
          8582 => x"84",
          8583 => x"80",
          8584 => x"90",
          8585 => x"81",
          8586 => x"a3",
          8587 => x"1a",
          8588 => x"9b",
          8589 => x"57",
          8590 => x"39",
          8591 => x"fe",
          8592 => x"53",
          8593 => x"51",
          8594 => x"84",
          8595 => x"84",
          8596 => x"30",
          8597 => x"84",
          8598 => x"25",
          8599 => x"7a",
          8600 => x"74",
          8601 => x"75",
          8602 => x"9c",
          8603 => x"05",
          8604 => x"56",
          8605 => x"26",
          8606 => x"15",
          8607 => x"84",
          8608 => x"07",
          8609 => x"1a",
          8610 => x"74",
          8611 => x"0c",
          8612 => x"04",
          8613 => x"bb",
          8614 => x"3d",
          8615 => x"bb",
          8616 => x"fe",
          8617 => x"80",
          8618 => x"38",
          8619 => x"52",
          8620 => x"8b",
          8621 => x"84",
          8622 => x"a7",
          8623 => x"84",
          8624 => x"84",
          8625 => x"0d",
          8626 => x"74",
          8627 => x"b9",
          8628 => x"ff",
          8629 => x"3d",
          8630 => x"71",
          8631 => x"58",
          8632 => x"0a",
          8633 => x"38",
          8634 => x"53",
          8635 => x"38",
          8636 => x"0c",
          8637 => x"55",
          8638 => x"38",
          8639 => x"75",
          8640 => x"cc",
          8641 => x"2a",
          8642 => x"88",
          8643 => x"56",
          8644 => x"a9",
          8645 => x"08",
          8646 => x"74",
          8647 => x"98",
          8648 => x"82",
          8649 => x"2e",
          8650 => x"89",
          8651 => x"19",
          8652 => x"ff",
          8653 => x"05",
          8654 => x"80",
          8655 => x"bb",
          8656 => x"3d",
          8657 => x"0b",
          8658 => x"0c",
          8659 => x"04",
          8660 => x"55",
          8661 => x"ff",
          8662 => x"17",
          8663 => x"2b",
          8664 => x"76",
          8665 => x"9c",
          8666 => x"fe",
          8667 => x"54",
          8668 => x"75",
          8669 => x"38",
          8670 => x"76",
          8671 => x"19",
          8672 => x"53",
          8673 => x"0c",
          8674 => x"74",
          8675 => x"ec",
          8676 => x"bb",
          8677 => x"84",
          8678 => x"ff",
          8679 => x"81",
          8680 => x"84",
          8681 => x"9e",
          8682 => x"08",
          8683 => x"84",
          8684 => x"ff",
          8685 => x"76",
          8686 => x"76",
          8687 => x"ff",
          8688 => x"0b",
          8689 => x"0c",
          8690 => x"04",
          8691 => x"7f",
          8692 => x"12",
          8693 => x"5c",
          8694 => x"80",
          8695 => x"86",
          8696 => x"98",
          8697 => x"17",
          8698 => x"56",
          8699 => x"b2",
          8700 => x"ff",
          8701 => x"9d",
          8702 => x"94",
          8703 => x"58",
          8704 => x"79",
          8705 => x"1a",
          8706 => x"74",
          8707 => x"f5",
          8708 => x"18",
          8709 => x"18",
          8710 => x"b8",
          8711 => x"0c",
          8712 => x"84",
          8713 => x"8f",
          8714 => x"77",
          8715 => x"8a",
          8716 => x"05",
          8717 => x"06",
          8718 => x"38",
          8719 => x"51",
          8720 => x"84",
          8721 => x"5d",
          8722 => x"0b",
          8723 => x"08",
          8724 => x"81",
          8725 => x"84",
          8726 => x"c6",
          8727 => x"08",
          8728 => x"08",
          8729 => x"38",
          8730 => x"81",
          8731 => x"17",
          8732 => x"51",
          8733 => x"84",
          8734 => x"5d",
          8735 => x"bb",
          8736 => x"2e",
          8737 => x"82",
          8738 => x"84",
          8739 => x"ff",
          8740 => x"56",
          8741 => x"08",
          8742 => x"86",
          8743 => x"84",
          8744 => x"33",
          8745 => x"80",
          8746 => x"18",
          8747 => x"fe",
          8748 => x"80",
          8749 => x"27",
          8750 => x"19",
          8751 => x"29",
          8752 => x"05",
          8753 => x"b4",
          8754 => x"19",
          8755 => x"78",
          8756 => x"76",
          8757 => x"58",
          8758 => x"55",
          8759 => x"74",
          8760 => x"22",
          8761 => x"27",
          8762 => x"81",
          8763 => x"53",
          8764 => x"19",
          8765 => x"b2",
          8766 => x"84",
          8767 => x"38",
          8768 => x"dd",
          8769 => x"18",
          8770 => x"84",
          8771 => x"8f",
          8772 => x"75",
          8773 => x"08",
          8774 => x"70",
          8775 => x"33",
          8776 => x"86",
          8777 => x"84",
          8778 => x"38",
          8779 => x"08",
          8780 => x"b4",
          8781 => x"1a",
          8782 => x"74",
          8783 => x"27",
          8784 => x"82",
          8785 => x"7b",
          8786 => x"81",
          8787 => x"38",
          8788 => x"19",
          8789 => x"08",
          8790 => x"52",
          8791 => x"51",
          8792 => x"fe",
          8793 => x"19",
          8794 => x"83",
          8795 => x"55",
          8796 => x"09",
          8797 => x"38",
          8798 => x"0c",
          8799 => x"1a",
          8800 => x"5e",
          8801 => x"75",
          8802 => x"85",
          8803 => x"22",
          8804 => x"b0",
          8805 => x"98",
          8806 => x"fc",
          8807 => x"0b",
          8808 => x"0c",
          8809 => x"04",
          8810 => x"64",
          8811 => x"84",
          8812 => x"5b",
          8813 => x"98",
          8814 => x"5e",
          8815 => x"2e",
          8816 => x"b8",
          8817 => x"5a",
          8818 => x"19",
          8819 => x"82",
          8820 => x"19",
          8821 => x"55",
          8822 => x"09",
          8823 => x"94",
          8824 => x"75",
          8825 => x"52",
          8826 => x"51",
          8827 => x"84",
          8828 => x"80",
          8829 => x"ff",
          8830 => x"79",
          8831 => x"76",
          8832 => x"90",
          8833 => x"08",
          8834 => x"58",
          8835 => x"82",
          8836 => x"18",
          8837 => x"70",
          8838 => x"5b",
          8839 => x"1d",
          8840 => x"e5",
          8841 => x"78",
          8842 => x"30",
          8843 => x"71",
          8844 => x"54",
          8845 => x"55",
          8846 => x"74",
          8847 => x"43",
          8848 => x"2e",
          8849 => x"75",
          8850 => x"86",
          8851 => x"5d",
          8852 => x"51",
          8853 => x"84",
          8854 => x"5b",
          8855 => x"08",
          8856 => x"98",
          8857 => x"75",
          8858 => x"7a",
          8859 => x"0c",
          8860 => x"04",
          8861 => x"19",
          8862 => x"52",
          8863 => x"51",
          8864 => x"81",
          8865 => x"84",
          8866 => x"09",
          8867 => x"ef",
          8868 => x"84",
          8869 => x"34",
          8870 => x"a8",
          8871 => x"84",
          8872 => x"58",
          8873 => x"1a",
          8874 => x"b5",
          8875 => x"33",
          8876 => x"2e",
          8877 => x"fe",
          8878 => x"54",
          8879 => x"a0",
          8880 => x"53",
          8881 => x"19",
          8882 => x"de",
          8883 => x"fe",
          8884 => x"8f",
          8885 => x"06",
          8886 => x"76",
          8887 => x"06",
          8888 => x"2e",
          8889 => x"18",
          8890 => x"bf",
          8891 => x"1f",
          8892 => x"05",
          8893 => x"5e",
          8894 => x"ab",
          8895 => x"55",
          8896 => x"cc",
          8897 => x"75",
          8898 => x"81",
          8899 => x"38",
          8900 => x"5b",
          8901 => x"1d",
          8902 => x"bb",
          8903 => x"3d",
          8904 => x"5b",
          8905 => x"8d",
          8906 => x"7d",
          8907 => x"81",
          8908 => x"8c",
          8909 => x"19",
          8910 => x"33",
          8911 => x"07",
          8912 => x"75",
          8913 => x"77",
          8914 => x"bf",
          8915 => x"f3",
          8916 => x"81",
          8917 => x"83",
          8918 => x"33",
          8919 => x"11",
          8920 => x"71",
          8921 => x"52",
          8922 => x"80",
          8923 => x"38",
          8924 => x"26",
          8925 => x"79",
          8926 => x"76",
          8927 => x"62",
          8928 => x"5a",
          8929 => x"8c",
          8930 => x"38",
          8931 => x"86",
          8932 => x"59",
          8933 => x"2e",
          8934 => x"81",
          8935 => x"dd",
          8936 => x"61",
          8937 => x"63",
          8938 => x"70",
          8939 => x"5e",
          8940 => x"39",
          8941 => x"ff",
          8942 => x"81",
          8943 => x"c0",
          8944 => x"38",
          8945 => x"57",
          8946 => x"75",
          8947 => x"05",
          8948 => x"05",
          8949 => x"7f",
          8950 => x"ff",
          8951 => x"59",
          8952 => x"e4",
          8953 => x"2e",
          8954 => x"ff",
          8955 => x"0c",
          8956 => x"84",
          8957 => x"0d",
          8958 => x"0d",
          8959 => x"5c",
          8960 => x"7b",
          8961 => x"3f",
          8962 => x"08",
          8963 => x"84",
          8964 => x"38",
          8965 => x"40",
          8966 => x"ac",
          8967 => x"1b",
          8968 => x"08",
          8969 => x"b4",
          8970 => x"2e",
          8971 => x"83",
          8972 => x"58",
          8973 => x"2e",
          8974 => x"81",
          8975 => x"54",
          8976 => x"1b",
          8977 => x"33",
          8978 => x"3f",
          8979 => x"08",
          8980 => x"38",
          8981 => x"57",
          8982 => x"0c",
          8983 => x"81",
          8984 => x"1c",
          8985 => x"58",
          8986 => x"2e",
          8987 => x"8b",
          8988 => x"06",
          8989 => x"06",
          8990 => x"86",
          8991 => x"81",
          8992 => x"f2",
          8993 => x"2a",
          8994 => x"75",
          8995 => x"ef",
          8996 => x"e2",
          8997 => x"2e",
          8998 => x"7c",
          8999 => x"7d",
          9000 => x"57",
          9001 => x"75",
          9002 => x"05",
          9003 => x"05",
          9004 => x"76",
          9005 => x"ff",
          9006 => x"59",
          9007 => x"e4",
          9008 => x"2e",
          9009 => x"ab",
          9010 => x"06",
          9011 => x"38",
          9012 => x"1d",
          9013 => x"70",
          9014 => x"33",
          9015 => x"05",
          9016 => x"71",
          9017 => x"5a",
          9018 => x"76",
          9019 => x"dc",
          9020 => x"2e",
          9021 => x"ff",
          9022 => x"ac",
          9023 => x"52",
          9024 => x"c8",
          9025 => x"84",
          9026 => x"bb",
          9027 => x"2e",
          9028 => x"79",
          9029 => x"0c",
          9030 => x"04",
          9031 => x"1b",
          9032 => x"52",
          9033 => x"51",
          9034 => x"81",
          9035 => x"84",
          9036 => x"09",
          9037 => x"a4",
          9038 => x"84",
          9039 => x"34",
          9040 => x"a8",
          9041 => x"84",
          9042 => x"58",
          9043 => x"1c",
          9044 => x"ea",
          9045 => x"33",
          9046 => x"2e",
          9047 => x"fd",
          9048 => x"54",
          9049 => x"a0",
          9050 => x"53",
          9051 => x"1b",
          9052 => x"b6",
          9053 => x"fd",
          9054 => x"5a",
          9055 => x"ab",
          9056 => x"86",
          9057 => x"42",
          9058 => x"f2",
          9059 => x"2a",
          9060 => x"79",
          9061 => x"38",
          9062 => x"77",
          9063 => x"70",
          9064 => x"7f",
          9065 => x"59",
          9066 => x"7d",
          9067 => x"81",
          9068 => x"5d",
          9069 => x"51",
          9070 => x"84",
          9071 => x"5a",
          9072 => x"08",
          9073 => x"d9",
          9074 => x"39",
          9075 => x"fe",
          9076 => x"ff",
          9077 => x"ac",
          9078 => x"a2",
          9079 => x"33",
          9080 => x"2e",
          9081 => x"c7",
          9082 => x"08",
          9083 => x"9a",
          9084 => x"88",
          9085 => x"42",
          9086 => x"b3",
          9087 => x"70",
          9088 => x"29",
          9089 => x"55",
          9090 => x"56",
          9091 => x"18",
          9092 => x"81",
          9093 => x"33",
          9094 => x"07",
          9095 => x"75",
          9096 => x"ed",
          9097 => x"fe",
          9098 => x"38",
          9099 => x"a0",
          9100 => x"bb",
          9101 => x"10",
          9102 => x"22",
          9103 => x"1b",
          9104 => x"a0",
          9105 => x"84",
          9106 => x"2e",
          9107 => x"fe",
          9108 => x"56",
          9109 => x"8c",
          9110 => x"b0",
          9111 => x"70",
          9112 => x"06",
          9113 => x"80",
          9114 => x"74",
          9115 => x"38",
          9116 => x"05",
          9117 => x"41",
          9118 => x"38",
          9119 => x"81",
          9120 => x"5a",
          9121 => x"84",
          9122 => x"84",
          9123 => x"0d",
          9124 => x"ff",
          9125 => x"bc",
          9126 => x"55",
          9127 => x"ea",
          9128 => x"70",
          9129 => x"13",
          9130 => x"06",
          9131 => x"5e",
          9132 => x"85",
          9133 => x"8c",
          9134 => x"22",
          9135 => x"74",
          9136 => x"38",
          9137 => x"10",
          9138 => x"51",
          9139 => x"f4",
          9140 => x"a0",
          9141 => x"8c",
          9142 => x"58",
          9143 => x"81",
          9144 => x"77",
          9145 => x"59",
          9146 => x"55",
          9147 => x"02",
          9148 => x"33",
          9149 => x"58",
          9150 => x"2e",
          9151 => x"80",
          9152 => x"1f",
          9153 => x"94",
          9154 => x"8c",
          9155 => x"58",
          9156 => x"61",
          9157 => x"77",
          9158 => x"59",
          9159 => x"81",
          9160 => x"ff",
          9161 => x"ef",
          9162 => x"27",
          9163 => x"7a",
          9164 => x"57",
          9165 => x"b8",
          9166 => x"1a",
          9167 => x"58",
          9168 => x"77",
          9169 => x"81",
          9170 => x"ff",
          9171 => x"90",
          9172 => x"44",
          9173 => x"60",
          9174 => x"38",
          9175 => x"a1",
          9176 => x"18",
          9177 => x"25",
          9178 => x"22",
          9179 => x"38",
          9180 => x"05",
          9181 => x"57",
          9182 => x"07",
          9183 => x"b9",
          9184 => x"38",
          9185 => x"74",
          9186 => x"16",
          9187 => x"84",
          9188 => x"56",
          9189 => x"77",
          9190 => x"fe",
          9191 => x"7a",
          9192 => x"78",
          9193 => x"79",
          9194 => x"a0",
          9195 => x"81",
          9196 => x"78",
          9197 => x"38",
          9198 => x"33",
          9199 => x"a0",
          9200 => x"06",
          9201 => x"16",
          9202 => x"77",
          9203 => x"38",
          9204 => x"05",
          9205 => x"19",
          9206 => x"59",
          9207 => x"34",
          9208 => x"87",
          9209 => x"51",
          9210 => x"84",
          9211 => x"8b",
          9212 => x"5b",
          9213 => x"27",
          9214 => x"87",
          9215 => x"e4",
          9216 => x"38",
          9217 => x"08",
          9218 => x"84",
          9219 => x"09",
          9220 => x"d6",
          9221 => x"db",
          9222 => x"1f",
          9223 => x"02",
          9224 => x"db",
          9225 => x"58",
          9226 => x"81",
          9227 => x"5b",
          9228 => x"90",
          9229 => x"8c",
          9230 => x"88",
          9231 => x"bb",
          9232 => x"5b",
          9233 => x"51",
          9234 => x"84",
          9235 => x"56",
          9236 => x"08",
          9237 => x"84",
          9238 => x"b8",
          9239 => x"98",
          9240 => x"80",
          9241 => x"08",
          9242 => x"f3",
          9243 => x"33",
          9244 => x"2e",
          9245 => x"82",
          9246 => x"54",
          9247 => x"18",
          9248 => x"33",
          9249 => x"3f",
          9250 => x"08",
          9251 => x"38",
          9252 => x"57",
          9253 => x"0c",
          9254 => x"bc",
          9255 => x"08",
          9256 => x"42",
          9257 => x"2e",
          9258 => x"74",
          9259 => x"25",
          9260 => x"5f",
          9261 => x"81",
          9262 => x"19",
          9263 => x"2e",
          9264 => x"81",
          9265 => x"ee",
          9266 => x"bb",
          9267 => x"84",
          9268 => x"80",
          9269 => x"38",
          9270 => x"84",
          9271 => x"38",
          9272 => x"81",
          9273 => x"1b",
          9274 => x"f3",
          9275 => x"08",
          9276 => x"08",
          9277 => x"38",
          9278 => x"78",
          9279 => x"84",
          9280 => x"54",
          9281 => x"1c",
          9282 => x"33",
          9283 => x"3f",
          9284 => x"08",
          9285 => x"38",
          9286 => x"56",
          9287 => x"0c",
          9288 => x"80",
          9289 => x"0b",
          9290 => x"57",
          9291 => x"70",
          9292 => x"34",
          9293 => x"74",
          9294 => x"0b",
          9295 => x"7b",
          9296 => x"75",
          9297 => x"57",
          9298 => x"81",
          9299 => x"ff",
          9300 => x"ef",
          9301 => x"08",
          9302 => x"98",
          9303 => x"7c",
          9304 => x"81",
          9305 => x"34",
          9306 => x"84",
          9307 => x"98",
          9308 => x"81",
          9309 => x"80",
          9310 => x"57",
          9311 => x"fe",
          9312 => x"59",
          9313 => x"51",
          9314 => x"84",
          9315 => x"56",
          9316 => x"08",
          9317 => x"c7",
          9318 => x"39",
          9319 => x"18",
          9320 => x"52",
          9321 => x"51",
          9322 => x"84",
          9323 => x"77",
          9324 => x"06",
          9325 => x"84",
          9326 => x"83",
          9327 => x"18",
          9328 => x"08",
          9329 => x"a0",
          9330 => x"8b",
          9331 => x"33",
          9332 => x"2e",
          9333 => x"84",
          9334 => x"57",
          9335 => x"7f",
          9336 => x"1f",
          9337 => x"53",
          9338 => x"e9",
          9339 => x"bb",
          9340 => x"84",
          9341 => x"fe",
          9342 => x"84",
          9343 => x"56",
          9344 => x"74",
          9345 => x"81",
          9346 => x"78",
          9347 => x"5a",
          9348 => x"05",
          9349 => x"06",
          9350 => x"56",
          9351 => x"38",
          9352 => x"06",
          9353 => x"41",
          9354 => x"57",
          9355 => x"1c",
          9356 => x"b2",
          9357 => x"33",
          9358 => x"2e",
          9359 => x"82",
          9360 => x"54",
          9361 => x"1c",
          9362 => x"33",
          9363 => x"3f",
          9364 => x"08",
          9365 => x"38",
          9366 => x"56",
          9367 => x"0c",
          9368 => x"fe",
          9369 => x"1c",
          9370 => x"08",
          9371 => x"06",
          9372 => x"60",
          9373 => x"8f",
          9374 => x"34",
          9375 => x"34",
          9376 => x"34",
          9377 => x"34",
          9378 => x"f3",
          9379 => x"5a",
          9380 => x"83",
          9381 => x"8b",
          9382 => x"1f",
          9383 => x"1b",
          9384 => x"83",
          9385 => x"33",
          9386 => x"76",
          9387 => x"05",
          9388 => x"88",
          9389 => x"75",
          9390 => x"38",
          9391 => x"57",
          9392 => x"8c",
          9393 => x"38",
          9394 => x"ff",
          9395 => x"38",
          9396 => x"70",
          9397 => x"76",
          9398 => x"a6",
          9399 => x"34",
          9400 => x"1d",
          9401 => x"7d",
          9402 => x"3f",
          9403 => x"08",
          9404 => x"84",
          9405 => x"38",
          9406 => x"40",
          9407 => x"38",
          9408 => x"81",
          9409 => x"08",
          9410 => x"70",
          9411 => x"33",
          9412 => x"96",
          9413 => x"84",
          9414 => x"fc",
          9415 => x"bb",
          9416 => x"1d",
          9417 => x"08",
          9418 => x"31",
          9419 => x"08",
          9420 => x"a0",
          9421 => x"fb",
          9422 => x"1c",
          9423 => x"82",
          9424 => x"06",
          9425 => x"81",
          9426 => x"08",
          9427 => x"05",
          9428 => x"81",
          9429 => x"cf",
          9430 => x"56",
          9431 => x"76",
          9432 => x"70",
          9433 => x"56",
          9434 => x"2e",
          9435 => x"fa",
          9436 => x"ff",
          9437 => x"57",
          9438 => x"2e",
          9439 => x"fa",
          9440 => x"80",
          9441 => x"fe",
          9442 => x"54",
          9443 => x"53",
          9444 => x"1c",
          9445 => x"92",
          9446 => x"84",
          9447 => x"09",
          9448 => x"38",
          9449 => x"08",
          9450 => x"b4",
          9451 => x"1d",
          9452 => x"74",
          9453 => x"27",
          9454 => x"1c",
          9455 => x"82",
          9456 => x"84",
          9457 => x"56",
          9458 => x"75",
          9459 => x"58",
          9460 => x"fa",
          9461 => x"87",
          9462 => x"57",
          9463 => x"81",
          9464 => x"75",
          9465 => x"fe",
          9466 => x"39",
          9467 => x"1c",
          9468 => x"08",
          9469 => x"52",
          9470 => x"51",
          9471 => x"fc",
          9472 => x"54",
          9473 => x"a0",
          9474 => x"53",
          9475 => x"18",
          9476 => x"96",
          9477 => x"39",
          9478 => x"7f",
          9479 => x"40",
          9480 => x"0b",
          9481 => x"98",
          9482 => x"2e",
          9483 => x"ac",
          9484 => x"2e",
          9485 => x"80",
          9486 => x"8c",
          9487 => x"22",
          9488 => x"5c",
          9489 => x"2e",
          9490 => x"54",
          9491 => x"22",
          9492 => x"55",
          9493 => x"95",
          9494 => x"80",
          9495 => x"ff",
          9496 => x"5a",
          9497 => x"26",
          9498 => x"73",
          9499 => x"11",
          9500 => x"58",
          9501 => x"d4",
          9502 => x"70",
          9503 => x"30",
          9504 => x"5c",
          9505 => x"94",
          9506 => x"0b",
          9507 => x"80",
          9508 => x"59",
          9509 => x"1c",
          9510 => x"33",
          9511 => x"56",
          9512 => x"2e",
          9513 => x"85",
          9514 => x"38",
          9515 => x"70",
          9516 => x"07",
          9517 => x"5b",
          9518 => x"26",
          9519 => x"80",
          9520 => x"ae",
          9521 => x"05",
          9522 => x"18",
          9523 => x"70",
          9524 => x"34",
          9525 => x"8a",
          9526 => x"ba",
          9527 => x"88",
          9528 => x"0b",
          9529 => x"96",
          9530 => x"72",
          9531 => x"81",
          9532 => x"0b",
          9533 => x"81",
          9534 => x"94",
          9535 => x"0b",
          9536 => x"9c",
          9537 => x"11",
          9538 => x"73",
          9539 => x"89",
          9540 => x"1c",
          9541 => x"13",
          9542 => x"34",
          9543 => x"9c",
          9544 => x"33",
          9545 => x"71",
          9546 => x"88",
          9547 => x"14",
          9548 => x"07",
          9549 => x"33",
          9550 => x"0c",
          9551 => x"33",
          9552 => x"71",
          9553 => x"5f",
          9554 => x"5a",
          9555 => x"77",
          9556 => x"99",
          9557 => x"16",
          9558 => x"2b",
          9559 => x"7b",
          9560 => x"8f",
          9561 => x"81",
          9562 => x"c0",
          9563 => x"96",
          9564 => x"7a",
          9565 => x"57",
          9566 => x"7a",
          9567 => x"07",
          9568 => x"d0",
          9569 => x"84",
          9570 => x"ff",
          9571 => x"ff",
          9572 => x"38",
          9573 => x"81",
          9574 => x"88",
          9575 => x"7a",
          9576 => x"18",
          9577 => x"05",
          9578 => x"8c",
          9579 => x"5b",
          9580 => x"11",
          9581 => x"57",
          9582 => x"90",
          9583 => x"39",
          9584 => x"30",
          9585 => x"80",
          9586 => x"25",
          9587 => x"57",
          9588 => x"38",
          9589 => x"81",
          9590 => x"80",
          9591 => x"08",
          9592 => x"39",
          9593 => x"1f",
          9594 => x"57",
          9595 => x"fe",
          9596 => x"96",
          9597 => x"59",
          9598 => x"33",
          9599 => x"5a",
          9600 => x"26",
          9601 => x"1c",
          9602 => x"33",
          9603 => x"76",
          9604 => x"72",
          9605 => x"72",
          9606 => x"7d",
          9607 => x"38",
          9608 => x"83",
          9609 => x"55",
          9610 => x"70",
          9611 => x"34",
          9612 => x"16",
          9613 => x"89",
          9614 => x"57",
          9615 => x"79",
          9616 => x"fd",
          9617 => x"83",
          9618 => x"39",
          9619 => x"70",
          9620 => x"30",
          9621 => x"5d",
          9622 => x"a9",
          9623 => x"0d",
          9624 => x"70",
          9625 => x"80",
          9626 => x"57",
          9627 => x"af",
          9628 => x"81",
          9629 => x"dc",
          9630 => x"38",
          9631 => x"81",
          9632 => x"16",
          9633 => x"0c",
          9634 => x"3d",
          9635 => x"42",
          9636 => x"27",
          9637 => x"73",
          9638 => x"08",
          9639 => x"61",
          9640 => x"05",
          9641 => x"53",
          9642 => x"38",
          9643 => x"73",
          9644 => x"ec",
          9645 => x"ff",
          9646 => x"38",
          9647 => x"56",
          9648 => x"81",
          9649 => x"83",
          9650 => x"70",
          9651 => x"30",
          9652 => x"71",
          9653 => x"57",
          9654 => x"73",
          9655 => x"74",
          9656 => x"82",
          9657 => x"80",
          9658 => x"38",
          9659 => x"0b",
          9660 => x"33",
          9661 => x"06",
          9662 => x"73",
          9663 => x"ab",
          9664 => x"2e",
          9665 => x"16",
          9666 => x"81",
          9667 => x"54",
          9668 => x"38",
          9669 => x"06",
          9670 => x"84",
          9671 => x"fe",
          9672 => x"38",
          9673 => x"5d",
          9674 => x"81",
          9675 => x"70",
          9676 => x"33",
          9677 => x"73",
          9678 => x"f0",
          9679 => x"39",
          9680 => x"dc",
          9681 => x"70",
          9682 => x"07",
          9683 => x"55",
          9684 => x"a1",
          9685 => x"70",
          9686 => x"74",
          9687 => x"72",
          9688 => x"38",
          9689 => x"32",
          9690 => x"80",
          9691 => x"51",
          9692 => x"e1",
          9693 => x"1d",
          9694 => x"96",
          9695 => x"41",
          9696 => x"9f",
          9697 => x"38",
          9698 => x"b5",
          9699 => x"81",
          9700 => x"84",
          9701 => x"83",
          9702 => x"54",
          9703 => x"38",
          9704 => x"84",
          9705 => x"93",
          9706 => x"83",
          9707 => x"70",
          9708 => x"5c",
          9709 => x"2e",
          9710 => x"e4",
          9711 => x"0b",
          9712 => x"80",
          9713 => x"de",
          9714 => x"bb",
          9715 => x"bb",
          9716 => x"3d",
          9717 => x"73",
          9718 => x"70",
          9719 => x"25",
          9720 => x"55",
          9721 => x"80",
          9722 => x"81",
          9723 => x"62",
          9724 => x"55",
          9725 => x"2e",
          9726 => x"80",
          9727 => x"30",
          9728 => x"78",
          9729 => x"59",
          9730 => x"73",
          9731 => x"75",
          9732 => x"5a",
          9733 => x"84",
          9734 => x"82",
          9735 => x"38",
          9736 => x"76",
          9737 => x"38",
          9738 => x"11",
          9739 => x"22",
          9740 => x"70",
          9741 => x"2a",
          9742 => x"5f",
          9743 => x"ae",
          9744 => x"72",
          9745 => x"17",
          9746 => x"38",
          9747 => x"19",
          9748 => x"23",
          9749 => x"fe",
          9750 => x"78",
          9751 => x"ff",
          9752 => x"58",
          9753 => x"7a",
          9754 => x"e6",
          9755 => x"ff",
          9756 => x"72",
          9757 => x"f1",
          9758 => x"2e",
          9759 => x"19",
          9760 => x"22",
          9761 => x"ae",
          9762 => x"76",
          9763 => x"05",
          9764 => x"57",
          9765 => x"8f",
          9766 => x"70",
          9767 => x"7c",
          9768 => x"81",
          9769 => x"8b",
          9770 => x"55",
          9771 => x"70",
          9772 => x"34",
          9773 => x"72",
          9774 => x"73",
          9775 => x"78",
          9776 => x"81",
          9777 => x"54",
          9778 => x"2e",
          9779 => x"74",
          9780 => x"d0",
          9781 => x"32",
          9782 => x"80",
          9783 => x"54",
          9784 => x"85",
          9785 => x"83",
          9786 => x"59",
          9787 => x"83",
          9788 => x"75",
          9789 => x"30",
          9790 => x"80",
          9791 => x"07",
          9792 => x"54",
          9793 => x"83",
          9794 => x"8b",
          9795 => x"38",
          9796 => x"8a",
          9797 => x"07",
          9798 => x"26",
          9799 => x"56",
          9800 => x"7e",
          9801 => x"fc",
          9802 => x"57",
          9803 => x"15",
          9804 => x"18",
          9805 => x"74",
          9806 => x"a0",
          9807 => x"76",
          9808 => x"83",
          9809 => x"88",
          9810 => x"38",
          9811 => x"58",
          9812 => x"82",
          9813 => x"83",
          9814 => x"83",
          9815 => x"38",
          9816 => x"81",
          9817 => x"9d",
          9818 => x"06",
          9819 => x"2e",
          9820 => x"90",
          9821 => x"82",
          9822 => x"5e",
          9823 => x"85",
          9824 => x"07",
          9825 => x"1d",
          9826 => x"e4",
          9827 => x"bb",
          9828 => x"1d",
          9829 => x"84",
          9830 => x"80",
          9831 => x"38",
          9832 => x"08",
          9833 => x"81",
          9834 => x"38",
          9835 => x"81",
          9836 => x"80",
          9837 => x"38",
          9838 => x"81",
          9839 => x"82",
          9840 => x"08",
          9841 => x"73",
          9842 => x"08",
          9843 => x"f9",
          9844 => x"16",
          9845 => x"11",
          9846 => x"40",
          9847 => x"a0",
          9848 => x"75",
          9849 => x"85",
          9850 => x"07",
          9851 => x"39",
          9852 => x"56",
          9853 => x"09",
          9854 => x"ac",
          9855 => x"54",
          9856 => x"09",
          9857 => x"a0",
          9858 => x"18",
          9859 => x"23",
          9860 => x"1d",
          9861 => x"54",
          9862 => x"83",
          9863 => x"73",
          9864 => x"05",
          9865 => x"13",
          9866 => x"27",
          9867 => x"a0",
          9868 => x"ab",
          9869 => x"51",
          9870 => x"84",
          9871 => x"ab",
          9872 => x"54",
          9873 => x"08",
          9874 => x"74",
          9875 => x"06",
          9876 => x"ce",
          9877 => x"33",
          9878 => x"81",
          9879 => x"74",
          9880 => x"cd",
          9881 => x"08",
          9882 => x"60",
          9883 => x"11",
          9884 => x"12",
          9885 => x"2b",
          9886 => x"41",
          9887 => x"7d",
          9888 => x"d8",
          9889 => x"1d",
          9890 => x"65",
          9891 => x"b7",
          9892 => x"55",
          9893 => x"fe",
          9894 => x"17",
          9895 => x"88",
          9896 => x"39",
          9897 => x"76",
          9898 => x"fd",
          9899 => x"82",
          9900 => x"06",
          9901 => x"59",
          9902 => x"2e",
          9903 => x"fd",
          9904 => x"82",
          9905 => x"98",
          9906 => x"a0",
          9907 => x"88",
          9908 => x"06",
          9909 => x"d6",
          9910 => x"0b",
          9911 => x"80",
          9912 => x"84",
          9913 => x"0d",
          9914 => x"ff",
          9915 => x"81",
          9916 => x"80",
          9917 => x"1d",
          9918 => x"26",
          9919 => x"79",
          9920 => x"77",
          9921 => x"5a",
          9922 => x"79",
          9923 => x"83",
          9924 => x"51",
          9925 => x"3f",
          9926 => x"08",
          9927 => x"06",
          9928 => x"81",
          9929 => x"78",
          9930 => x"38",
          9931 => x"06",
          9932 => x"11",
          9933 => x"74",
          9934 => x"ff",
          9935 => x"80",
          9936 => x"38",
          9937 => x"0b",
          9938 => x"33",
          9939 => x"06",
          9940 => x"73",
          9941 => x"e0",
          9942 => x"2e",
          9943 => x"19",
          9944 => x"81",
          9945 => x"54",
          9946 => x"38",
          9947 => x"06",
          9948 => x"d4",
          9949 => x"15",
          9950 => x"26",
          9951 => x"82",
          9952 => x"ff",
          9953 => x"ff",
          9954 => x"78",
          9955 => x"38",
          9956 => x"70",
          9957 => x"e0",
          9958 => x"ff",
          9959 => x"56",
          9960 => x"1b",
          9961 => x"74",
          9962 => x"1b",
          9963 => x"55",
          9964 => x"80",
          9965 => x"39",
          9966 => x"33",
          9967 => x"06",
          9968 => x"80",
          9969 => x"38",
          9970 => x"83",
          9971 => x"a0",
          9972 => x"55",
          9973 => x"81",
          9974 => x"39",
          9975 => x"33",
          9976 => x"33",
          9977 => x"71",
          9978 => x"77",
          9979 => x"0c",
          9980 => x"95",
          9981 => x"a0",
          9982 => x"2a",
          9983 => x"74",
          9984 => x"7c",
          9985 => x"5a",
          9986 => x"34",
          9987 => x"ff",
          9988 => x"83",
          9989 => x"33",
          9990 => x"81",
          9991 => x"81",
          9992 => x"38",
          9993 => x"74",
          9994 => x"06",
          9995 => x"f2",
          9996 => x"84",
          9997 => x"93",
          9998 => x"eb",
          9999 => x"69",
         10000 => x"80",
         10001 => x"42",
         10002 => x"61",
         10003 => x"08",
         10004 => x"42",
         10005 => x"85",
         10006 => x"70",
         10007 => x"33",
         10008 => x"56",
         10009 => x"2e",
         10010 => x"74",
         10011 => x"ba",
         10012 => x"38",
         10013 => x"33",
         10014 => x"24",
         10015 => x"75",
         10016 => x"e2",
         10017 => x"08",
         10018 => x"58",
         10019 => x"85",
         10020 => x"61",
         10021 => x"fe",
         10022 => x"5d",
         10023 => x"2e",
         10024 => x"17",
         10025 => x"bb",
         10026 => x"bb",
         10027 => x"ff",
         10028 => x"06",
         10029 => x"80",
         10030 => x"38",
         10031 => x"75",
         10032 => x"ba",
         10033 => x"81",
         10034 => x"52",
         10035 => x"51",
         10036 => x"3f",
         10037 => x"08",
         10038 => x"70",
         10039 => x"56",
         10040 => x"84",
         10041 => x"80",
         10042 => x"75",
         10043 => x"06",
         10044 => x"60",
         10045 => x"80",
         10046 => x"18",
         10047 => x"b4",
         10048 => x"7b",
         10049 => x"54",
         10050 => x"17",
         10051 => x"18",
         10052 => x"ff",
         10053 => x"84",
         10054 => x"7b",
         10055 => x"ff",
         10056 => x"74",
         10057 => x"84",
         10058 => x"38",
         10059 => x"33",
         10060 => x"33",
         10061 => x"07",
         10062 => x"56",
         10063 => x"d5",
         10064 => x"38",
         10065 => x"8b",
         10066 => x"f9",
         10067 => x"61",
         10068 => x"81",
         10069 => x"2e",
         10070 => x"8d",
         10071 => x"26",
         10072 => x"80",
         10073 => x"80",
         10074 => x"71",
         10075 => x"5e",
         10076 => x"80",
         10077 => x"06",
         10078 => x"80",
         10079 => x"80",
         10080 => x"71",
         10081 => x"57",
         10082 => x"38",
         10083 => x"83",
         10084 => x"12",
         10085 => x"2b",
         10086 => x"07",
         10087 => x"70",
         10088 => x"2b",
         10089 => x"07",
         10090 => x"43",
         10091 => x"75",
         10092 => x"80",
         10093 => x"82",
         10094 => x"c8",
         10095 => x"11",
         10096 => x"06",
         10097 => x"8d",
         10098 => x"26",
         10099 => x"78",
         10100 => x"76",
         10101 => x"c5",
         10102 => x"5f",
         10103 => x"18",
         10104 => x"77",
         10105 => x"c4",
         10106 => x"78",
         10107 => x"87",
         10108 => x"ca",
         10109 => x"c9",
         10110 => x"88",
         10111 => x"40",
         10112 => x"23",
         10113 => x"06",
         10114 => x"58",
         10115 => x"38",
         10116 => x"33",
         10117 => x"33",
         10118 => x"07",
         10119 => x"a4",
         10120 => x"17",
         10121 => x"82",
         10122 => x"90",
         10123 => x"2b",
         10124 => x"33",
         10125 => x"88",
         10126 => x"71",
         10127 => x"5a",
         10128 => x"42",
         10129 => x"33",
         10130 => x"33",
         10131 => x"07",
         10132 => x"58",
         10133 => x"81",
         10134 => x"1c",
         10135 => x"05",
         10136 => x"26",
         10137 => x"78",
         10138 => x"31",
         10139 => x"b5",
         10140 => x"84",
         10141 => x"bb",
         10142 => x"2e",
         10143 => x"84",
         10144 => x"80",
         10145 => x"f5",
         10146 => x"83",
         10147 => x"ff",
         10148 => x"38",
         10149 => x"9f",
         10150 => x"eb",
         10151 => x"82",
         10152 => x"19",
         10153 => x"19",
         10154 => x"70",
         10155 => x"7b",
         10156 => x"0c",
         10157 => x"83",
         10158 => x"38",
         10159 => x"5c",
         10160 => x"80",
         10161 => x"38",
         10162 => x"18",
         10163 => x"55",
         10164 => x"8d",
         10165 => x"19",
         10166 => x"7a",
         10167 => x"56",
         10168 => x"15",
         10169 => x"8d",
         10170 => x"18",
         10171 => x"38",
         10172 => x"18",
         10173 => x"90",
         10174 => x"80",
         10175 => x"34",
         10176 => x"86",
         10177 => x"77",
         10178 => x"dc",
         10179 => x"5d",
         10180 => x"dc",
         10181 => x"18",
         10182 => x"e4",
         10183 => x"0c",
         10184 => x"18",
         10185 => x"77",
         10186 => x"0c",
         10187 => x"04",
         10188 => x"bb",
         10189 => x"3d",
         10190 => x"33",
         10191 => x"81",
         10192 => x"57",
         10193 => x"26",
         10194 => x"17",
         10195 => x"06",
         10196 => x"59",
         10197 => x"87",
         10198 => x"7e",
         10199 => x"f4",
         10200 => x"7c",
         10201 => x"5b",
         10202 => x"05",
         10203 => x"70",
         10204 => x"33",
         10205 => x"5a",
         10206 => x"99",
         10207 => x"e0",
         10208 => x"ff",
         10209 => x"ff",
         10210 => x"77",
         10211 => x"38",
         10212 => x"81",
         10213 => x"55",
         10214 => x"9f",
         10215 => x"75",
         10216 => x"81",
         10217 => x"77",
         10218 => x"78",
         10219 => x"30",
         10220 => x"9f",
         10221 => x"5d",
         10222 => x"80",
         10223 => x"38",
         10224 => x"1e",
         10225 => x"7c",
         10226 => x"38",
         10227 => x"a9",
         10228 => x"2e",
         10229 => x"77",
         10230 => x"06",
         10231 => x"7d",
         10232 => x"80",
         10233 => x"39",
         10234 => x"57",
         10235 => x"e9",
         10236 => x"06",
         10237 => x"59",
         10238 => x"32",
         10239 => x"80",
         10240 => x"5a",
         10241 => x"83",
         10242 => x"81",
         10243 => x"a6",
         10244 => x"77",
         10245 => x"59",
         10246 => x"33",
         10247 => x"7a",
         10248 => x"38",
         10249 => x"33",
         10250 => x"33",
         10251 => x"71",
         10252 => x"83",
         10253 => x"70",
         10254 => x"2b",
         10255 => x"33",
         10256 => x"59",
         10257 => x"40",
         10258 => x"84",
         10259 => x"ff",
         10260 => x"57",
         10261 => x"25",
         10262 => x"84",
         10263 => x"33",
         10264 => x"9f",
         10265 => x"31",
         10266 => x"10",
         10267 => x"05",
         10268 => x"44",
         10269 => x"5b",
         10270 => x"5b",
         10271 => x"80",
         10272 => x"38",
         10273 => x"18",
         10274 => x"b4",
         10275 => x"55",
         10276 => x"ff",
         10277 => x"81",
         10278 => x"b8",
         10279 => x"17",
         10280 => x"b4",
         10281 => x"bb",
         10282 => x"2e",
         10283 => x"55",
         10284 => x"b4",
         10285 => x"58",
         10286 => x"81",
         10287 => x"33",
         10288 => x"07",
         10289 => x"58",
         10290 => x"d5",
         10291 => x"06",
         10292 => x"0b",
         10293 => x"57",
         10294 => x"e9",
         10295 => x"38",
         10296 => x"32",
         10297 => x"80",
         10298 => x"42",
         10299 => x"bc",
         10300 => x"e8",
         10301 => x"82",
         10302 => x"ff",
         10303 => x"0b",
         10304 => x"1e",
         10305 => x"7b",
         10306 => x"81",
         10307 => x"81",
         10308 => x"27",
         10309 => x"77",
         10310 => x"b7",
         10311 => x"84",
         10312 => x"83",
         10313 => x"d1",
         10314 => x"39",
         10315 => x"ee",
         10316 => x"b4",
         10317 => x"7b",
         10318 => x"5d",
         10319 => x"81",
         10320 => x"71",
         10321 => x"1b",
         10322 => x"56",
         10323 => x"80",
         10324 => x"80",
         10325 => x"85",
         10326 => x"18",
         10327 => x"40",
         10328 => x"70",
         10329 => x"33",
         10330 => x"05",
         10331 => x"71",
         10332 => x"5b",
         10333 => x"77",
         10334 => x"8e",
         10335 => x"2e",
         10336 => x"58",
         10337 => x"8d",
         10338 => x"93",
         10339 => x"bb",
         10340 => x"3d",
         10341 => x"58",
         10342 => x"fe",
         10343 => x"0b",
         10344 => x"83",
         10345 => x"5d",
         10346 => x"39",
         10347 => x"bb",
         10348 => x"3d",
         10349 => x"0b",
         10350 => x"83",
         10351 => x"5a",
         10352 => x"81",
         10353 => x"7a",
         10354 => x"5c",
         10355 => x"31",
         10356 => x"57",
         10357 => x"80",
         10358 => x"38",
         10359 => x"e1",
         10360 => x"81",
         10361 => x"e6",
         10362 => x"58",
         10363 => x"05",
         10364 => x"70",
         10365 => x"33",
         10366 => x"ff",
         10367 => x"42",
         10368 => x"2e",
         10369 => x"75",
         10370 => x"38",
         10371 => x"57",
         10372 => x"fc",
         10373 => x"58",
         10374 => x"80",
         10375 => x"80",
         10376 => x"71",
         10377 => x"57",
         10378 => x"2e",
         10379 => x"f9",
         10380 => x"1b",
         10381 => x"b4",
         10382 => x"2e",
         10383 => x"17",
         10384 => x"7a",
         10385 => x"06",
         10386 => x"81",
         10387 => x"b8",
         10388 => x"17",
         10389 => x"b0",
         10390 => x"bb",
         10391 => x"2e",
         10392 => x"58",
         10393 => x"b4",
         10394 => x"f9",
         10395 => x"84",
         10396 => x"b7",
         10397 => x"b6",
         10398 => x"88",
         10399 => x"5e",
         10400 => x"d5",
         10401 => x"06",
         10402 => x"b8",
         10403 => x"33",
         10404 => x"71",
         10405 => x"88",
         10406 => x"14",
         10407 => x"07",
         10408 => x"33",
         10409 => x"41",
         10410 => x"5c",
         10411 => x"8b",
         10412 => x"2e",
         10413 => x"f8",
         10414 => x"9c",
         10415 => x"33",
         10416 => x"71",
         10417 => x"88",
         10418 => x"14",
         10419 => x"07",
         10420 => x"33",
         10421 => x"44",
         10422 => x"5a",
         10423 => x"8a",
         10424 => x"2e",
         10425 => x"f8",
         10426 => x"a0",
         10427 => x"33",
         10428 => x"71",
         10429 => x"88",
         10430 => x"14",
         10431 => x"07",
         10432 => x"33",
         10433 => x"1e",
         10434 => x"a4",
         10435 => x"33",
         10436 => x"71",
         10437 => x"88",
         10438 => x"14",
         10439 => x"07",
         10440 => x"33",
         10441 => x"90",
         10442 => x"44",
         10443 => x"45",
         10444 => x"56",
         10445 => x"34",
         10446 => x"22",
         10447 => x"7c",
         10448 => x"23",
         10449 => x"23",
         10450 => x"0b",
         10451 => x"80",
         10452 => x"0c",
         10453 => x"7b",
         10454 => x"f0",
         10455 => x"7f",
         10456 => x"95",
         10457 => x"b4",
         10458 => x"b8",
         10459 => x"81",
         10460 => x"59",
         10461 => x"3f",
         10462 => x"08",
         10463 => x"81",
         10464 => x"38",
         10465 => x"08",
         10466 => x"b4",
         10467 => x"18",
         10468 => x"7f",
         10469 => x"27",
         10470 => x"17",
         10471 => x"82",
         10472 => x"38",
         10473 => x"08",
         10474 => x"39",
         10475 => x"80",
         10476 => x"38",
         10477 => x"8a",
         10478 => x"b8",
         10479 => x"fc",
         10480 => x"e3",
         10481 => x"e2",
         10482 => x"88",
         10483 => x"5a",
         10484 => x"f6",
         10485 => x"17",
         10486 => x"f6",
         10487 => x"e4",
         10488 => x"33",
         10489 => x"71",
         10490 => x"88",
         10491 => x"14",
         10492 => x"07",
         10493 => x"33",
         10494 => x"1e",
         10495 => x"82",
         10496 => x"44",
         10497 => x"f5",
         10498 => x"58",
         10499 => x"f9",
         10500 => x"58",
         10501 => x"75",
         10502 => x"a8",
         10503 => x"77",
         10504 => x"59",
         10505 => x"75",
         10506 => x"da",
         10507 => x"39",
         10508 => x"17",
         10509 => x"08",
         10510 => x"52",
         10511 => x"51",
         10512 => x"3f",
         10513 => x"f0",
         10514 => x"80",
         10515 => x"64",
         10516 => x"3d",
         10517 => x"ff",
         10518 => x"75",
         10519 => x"e9",
         10520 => x"81",
         10521 => x"70",
         10522 => x"55",
         10523 => x"80",
         10524 => x"ed",
         10525 => x"2e",
         10526 => x"84",
         10527 => x"54",
         10528 => x"80",
         10529 => x"10",
         10530 => x"cc",
         10531 => x"55",
         10532 => x"2e",
         10533 => x"74",
         10534 => x"73",
         10535 => x"38",
         10536 => x"62",
         10537 => x"0c",
         10538 => x"80",
         10539 => x"80",
         10540 => x"70",
         10541 => x"51",
         10542 => x"84",
         10543 => x"54",
         10544 => x"84",
         10545 => x"0d",
         10546 => x"84",
         10547 => x"92",
         10548 => x"75",
         10549 => x"70",
         10550 => x"56",
         10551 => x"89",
         10552 => x"82",
         10553 => x"ff",
         10554 => x"5c",
         10555 => x"2e",
         10556 => x"80",
         10557 => x"e6",
         10558 => x"5b",
         10559 => x"59",
         10560 => x"81",
         10561 => x"78",
         10562 => x"5a",
         10563 => x"12",
         10564 => x"76",
         10565 => x"38",
         10566 => x"81",
         10567 => x"54",
         10568 => x"57",
         10569 => x"89",
         10570 => x"70",
         10571 => x"57",
         10572 => x"70",
         10573 => x"54",
         10574 => x"09",
         10575 => x"38",
         10576 => x"38",
         10577 => x"70",
         10578 => x"07",
         10579 => x"07",
         10580 => x"79",
         10581 => x"38",
         10582 => x"1d",
         10583 => x"7b",
         10584 => x"38",
         10585 => x"98",
         10586 => x"24",
         10587 => x"79",
         10588 => x"fe",
         10589 => x"3d",
         10590 => x"84",
         10591 => x"05",
         10592 => x"89",
         10593 => x"2e",
         10594 => x"bf",
         10595 => x"9d",
         10596 => x"53",
         10597 => x"05",
         10598 => x"9f",
         10599 => x"84",
         10600 => x"bb",
         10601 => x"2e",
         10602 => x"7a",
         10603 => x"75",
         10604 => x"0c",
         10605 => x"04",
         10606 => x"52",
         10607 => x"52",
         10608 => x"3f",
         10609 => x"08",
         10610 => x"84",
         10611 => x"81",
         10612 => x"9c",
         10613 => x"80",
         10614 => x"38",
         10615 => x"83",
         10616 => x"84",
         10617 => x"38",
         10618 => x"59",
         10619 => x"38",
         10620 => x"81",
         10621 => x"80",
         10622 => x"38",
         10623 => x"33",
         10624 => x"71",
         10625 => x"61",
         10626 => x"58",
         10627 => x"7d",
         10628 => x"97",
         10629 => x"8e",
         10630 => x"0b",
         10631 => x"a1",
         10632 => x"34",
         10633 => x"91",
         10634 => x"56",
         10635 => x"17",
         10636 => x"57",
         10637 => x"9a",
         10638 => x"0b",
         10639 => x"7d",
         10640 => x"83",
         10641 => x"38",
         10642 => x"0b",
         10643 => x"80",
         10644 => x"34",
         10645 => x"19",
         10646 => x"9f",
         10647 => x"55",
         10648 => x"16",
         10649 => x"2e",
         10650 => x"7e",
         10651 => x"7c",
         10652 => x"57",
         10653 => x"7b",
         10654 => x"9c",
         10655 => x"26",
         10656 => x"82",
         10657 => x"0c",
         10658 => x"02",
         10659 => x"33",
         10660 => x"5c",
         10661 => x"25",
         10662 => x"86",
         10663 => x"5e",
         10664 => x"b8",
         10665 => x"82",
         10666 => x"c2",
         10667 => x"84",
         10668 => x"5d",
         10669 => x"b0",
         10670 => x"2a",
         10671 => x"7c",
         10672 => x"38",
         10673 => x"58",
         10674 => x"38",
         10675 => x"81",
         10676 => x"80",
         10677 => x"78",
         10678 => x"59",
         10679 => x"08",
         10680 => x"67",
         10681 => x"67",
         10682 => x"9a",
         10683 => x"88",
         10684 => x"33",
         10685 => x"57",
         10686 => x"2e",
         10687 => x"77",
         10688 => x"9c",
         10689 => x"33",
         10690 => x"71",
         10691 => x"88",
         10692 => x"14",
         10693 => x"07",
         10694 => x"33",
         10695 => x"8c",
         10696 => x"7f",
         10697 => x"58",
         10698 => x"86",
         10699 => x"1b",
         10700 => x"1b",
         10701 => x"91",
         10702 => x"0b",
         10703 => x"80",
         10704 => x"0c",
         10705 => x"84",
         10706 => x"55",
         10707 => x"81",
         10708 => x"ff",
         10709 => x"f4",
         10710 => x"2a",
         10711 => x"78",
         10712 => x"c9",
         10713 => x"08",
         10714 => x"2e",
         10715 => x"74",
         10716 => x"8a",
         10717 => x"89",
         10718 => x"08",
         10719 => x"5a",
         10720 => x"70",
         10721 => x"25",
         10722 => x"76",
         10723 => x"38",
         10724 => x"06",
         10725 => x"80",
         10726 => x"38",
         10727 => x"51",
         10728 => x"3f",
         10729 => x"08",
         10730 => x"84",
         10731 => x"83",
         10732 => x"84",
         10733 => x"ff",
         10734 => x"75",
         10735 => x"c1",
         10736 => x"c2",
         10737 => x"06",
         10738 => x"38",
         10739 => x"81",
         10740 => x"80",
         10741 => x"38",
         10742 => x"7a",
         10743 => x"39",
         10744 => x"7a",
         10745 => x"39",
         10746 => x"7a",
         10747 => x"39",
         10748 => x"31",
         10749 => x"89",
         10750 => x"33",
         10751 => x"71",
         10752 => x"90",
         10753 => x"07",
         10754 => x"9c",
         10755 => x"33",
         10756 => x"71",
         10757 => x"88",
         10758 => x"14",
         10759 => x"07",
         10760 => x"33",
         10761 => x"8c",
         10762 => x"61",
         10763 => x"5a",
         10764 => x"5e",
         10765 => x"22",
         10766 => x"78",
         10767 => x"80",
         10768 => x"34",
         10769 => x"1b",
         10770 => x"94",
         10771 => x"1a",
         10772 => x"7c",
         10773 => x"f4",
         10774 => x"cc",
         10775 => x"bb",
         10776 => x"88",
         10777 => x"76",
         10778 => x"fb",
         10779 => x"52",
         10780 => x"aa",
         10781 => x"bb",
         10782 => x"84",
         10783 => x"80",
         10784 => x"38",
         10785 => x"08",
         10786 => x"f7",
         10787 => x"84",
         10788 => x"82",
         10789 => x"53",
         10790 => x"51",
         10791 => x"3f",
         10792 => x"08",
         10793 => x"9c",
         10794 => x"11",
         10795 => x"59",
         10796 => x"75",
         10797 => x"81",
         10798 => x"0c",
         10799 => x"81",
         10800 => x"84",
         10801 => x"55",
         10802 => x"ff",
         10803 => x"7f",
         10804 => x"59",
         10805 => x"16",
         10806 => x"af",
         10807 => x"33",
         10808 => x"2e",
         10809 => x"81",
         10810 => x"54",
         10811 => x"16",
         10812 => x"33",
         10813 => x"b3",
         10814 => x"84",
         10815 => x"85",
         10816 => x"81",
         10817 => x"17",
         10818 => x"7b",
         10819 => x"18",
         10820 => x"80",
         10821 => x"38",
         10822 => x"f9",
         10823 => x"0b",
         10824 => x"80",
         10825 => x"34",
         10826 => x"95",
         10827 => x"17",
         10828 => x"2b",
         10829 => x"07",
         10830 => x"56",
         10831 => x"8e",
         10832 => x"0b",
         10833 => x"a1",
         10834 => x"34",
         10835 => x"91",
         10836 => x"56",
         10837 => x"17",
         10838 => x"57",
         10839 => x"9a",
         10840 => x"0b",
         10841 => x"7d",
         10842 => x"83",
         10843 => x"06",
         10844 => x"ff",
         10845 => x"98",
         10846 => x"f8",
         10847 => x"83",
         10848 => x"78",
         10849 => x"a5",
         10850 => x"19",
         10851 => x"fe",
         10852 => x"59",
         10853 => x"f9",
         10854 => x"19",
         10855 => x"29",
         10856 => x"05",
         10857 => x"80",
         10858 => x"38",
         10859 => x"15",
         10860 => x"0c",
         10861 => x"77",
         10862 => x"81",
         10863 => x"ff",
         10864 => x"84",
         10865 => x"80",
         10866 => x"38",
         10867 => x"7a",
         10868 => x"39",
         10869 => x"16",
         10870 => x"16",
         10871 => x"17",
         10872 => x"ff",
         10873 => x"84",
         10874 => x"7d",
         10875 => x"06",
         10876 => x"84",
         10877 => x"83",
         10878 => x"16",
         10879 => x"08",
         10880 => x"84",
         10881 => x"74",
         10882 => x"27",
         10883 => x"82",
         10884 => x"74",
         10885 => x"81",
         10886 => x"38",
         10887 => x"16",
         10888 => x"08",
         10889 => x"52",
         10890 => x"51",
         10891 => x"3f",
         10892 => x"b6",
         10893 => x"84",
         10894 => x"7a",
         10895 => x"39",
         10896 => x"c5",
         10897 => x"0d",
         10898 => x"64",
         10899 => x"59",
         10900 => x"89",
         10901 => x"2e",
         10902 => x"08",
         10903 => x"2e",
         10904 => x"33",
         10905 => x"2e",
         10906 => x"16",
         10907 => x"22",
         10908 => x"78",
         10909 => x"38",
         10910 => x"5f",
         10911 => x"81",
         10912 => x"19",
         10913 => x"81",
         10914 => x"19",
         10915 => x"57",
         10916 => x"80",
         10917 => x"38",
         10918 => x"8c",
         10919 => x"31",
         10920 => x"75",
         10921 => x"38",
         10922 => x"81",
         10923 => x"83",
         10924 => x"7b",
         10925 => x"7e",
         10926 => x"ff",
         10927 => x"2a",
         10928 => x"7b",
         10929 => x"82",
         10930 => x"19",
         10931 => x"75",
         10932 => x"38",
         10933 => x"83",
         10934 => x"98",
         10935 => x"58",
         10936 => x"fe",
         10937 => x"08",
         10938 => x"57",
         10939 => x"83",
         10940 => x"18",
         10941 => x"29",
         10942 => x"05",
         10943 => x"80",
         10944 => x"38",
         10945 => x"89",
         10946 => x"7a",
         10947 => x"e6",
         10948 => x"55",
         10949 => x"85",
         10950 => x"31",
         10951 => x"76",
         10952 => x"81",
         10953 => x"ff",
         10954 => x"84",
         10955 => x"82",
         10956 => x"19",
         10957 => x"2b",
         10958 => x"78",
         10959 => x"38",
         10960 => x"57",
         10961 => x"7e",
         10962 => x"0c",
         10963 => x"1b",
         10964 => x"59",
         10965 => x"5e",
         10966 => x"d2",
         10967 => x"75",
         10968 => x"0c",
         10969 => x"04",
         10970 => x"84",
         10971 => x"0d",
         10972 => x"fe",
         10973 => x"19",
         10974 => x"77",
         10975 => x"38",
         10976 => x"70",
         10977 => x"1b",
         10978 => x"7b",
         10979 => x"38",
         10980 => x"53",
         10981 => x"18",
         10982 => x"9f",
         10983 => x"bb",
         10984 => x"e3",
         10985 => x"33",
         10986 => x"55",
         10987 => x"34",
         10988 => x"54",
         10989 => x"52",
         10990 => x"51",
         10991 => x"3f",
         10992 => x"08",
         10993 => x"76",
         10994 => x"94",
         10995 => x"75",
         10996 => x"84",
         10997 => x"58",
         10998 => x"27",
         10999 => x"57",
         11000 => x"17",
         11001 => x"59",
         11002 => x"2e",
         11003 => x"74",
         11004 => x"56",
         11005 => x"81",
         11006 => x"ff",
         11007 => x"80",
         11008 => x"38",
         11009 => x"05",
         11010 => x"70",
         11011 => x"34",
         11012 => x"75",
         11013 => x"ac",
         11014 => x"08",
         11015 => x"ff",
         11016 => x"84",
         11017 => x"55",
         11018 => x"81",
         11019 => x"ff",
         11020 => x"84",
         11021 => x"81",
         11022 => x"fc",
         11023 => x"79",
         11024 => x"fc",
         11025 => x"19",
         11026 => x"56",
         11027 => x"fd",
         11028 => x"80",
         11029 => x"1e",
         11030 => x"58",
         11031 => x"81",
         11032 => x"77",
         11033 => x"59",
         11034 => x"55",
         11035 => x"fd",
         11036 => x"70",
         11037 => x"33",
         11038 => x"05",
         11039 => x"15",
         11040 => x"38",
         11041 => x"81",
         11042 => x"34",
         11043 => x"bb",
         11044 => x"3d",
         11045 => x"0b",
         11046 => x"82",
         11047 => x"84",
         11048 => x"0d",
         11049 => x"0d",
         11050 => x"65",
         11051 => x"59",
         11052 => x"89",
         11053 => x"2e",
         11054 => x"08",
         11055 => x"2e",
         11056 => x"33",
         11057 => x"2e",
         11058 => x"16",
         11059 => x"22",
         11060 => x"78",
         11061 => x"38",
         11062 => x"40",
         11063 => x"82",
         11064 => x"19",
         11065 => x"82",
         11066 => x"19",
         11067 => x"2a",
         11068 => x"58",
         11069 => x"80",
         11070 => x"38",
         11071 => x"7b",
         11072 => x"7b",
         11073 => x"38",
         11074 => x"7a",
         11075 => x"89",
         11076 => x"ff",
         11077 => x"82",
         11078 => x"8a",
         11079 => x"05",
         11080 => x"06",
         11081 => x"aa",
         11082 => x"f9",
         11083 => x"08",
         11084 => x"2e",
         11085 => x"74",
         11086 => x"ed",
         11087 => x"2e",
         11088 => x"74",
         11089 => x"88",
         11090 => x"38",
         11091 => x"0c",
         11092 => x"19",
         11093 => x"2b",
         11094 => x"7a",
         11095 => x"38",
         11096 => x"fe",
         11097 => x"08",
         11098 => x"57",
         11099 => x"83",
         11100 => x"18",
         11101 => x"29",
         11102 => x"05",
         11103 => x"80",
         11104 => x"38",
         11105 => x"89",
         11106 => x"79",
         11107 => x"a6",
         11108 => x"55",
         11109 => x"85",
         11110 => x"31",
         11111 => x"7b",
         11112 => x"81",
         11113 => x"ff",
         11114 => x"84",
         11115 => x"82",
         11116 => x"19",
         11117 => x"56",
         11118 => x"ab",
         11119 => x"0b",
         11120 => x"72",
         11121 => x"58",
         11122 => x"70",
         11123 => x"33",
         11124 => x"05",
         11125 => x"15",
         11126 => x"38",
         11127 => x"80",
         11128 => x"7c",
         11129 => x"79",
         11130 => x"7a",
         11131 => x"08",
         11132 => x"78",
         11133 => x"08",
         11134 => x"94",
         11135 => x"1d",
         11136 => x"58",
         11137 => x"76",
         11138 => x"75",
         11139 => x"1a",
         11140 => x"fd",
         11141 => x"33",
         11142 => x"c0",
         11143 => x"90",
         11144 => x"56",
         11145 => x"84",
         11146 => x"0d",
         11147 => x"bb",
         11148 => x"3d",
         11149 => x"19",
         11150 => x"a2",
         11151 => x"08",
         11152 => x"1a",
         11153 => x"38",
         11154 => x"53",
         11155 => x"81",
         11156 => x"ff",
         11157 => x"84",
         11158 => x"81",
         11159 => x"19",
         11160 => x"9c",
         11161 => x"83",
         11162 => x"80",
         11163 => x"55",
         11164 => x"83",
         11165 => x"77",
         11166 => x"05",
         11167 => x"56",
         11168 => x"93",
         11169 => x"81",
         11170 => x"75",
         11171 => x"57",
         11172 => x"56",
         11173 => x"90",
         11174 => x"80",
         11175 => x"90",
         11176 => x"c7",
         11177 => x"08",
         11178 => x"ff",
         11179 => x"84",
         11180 => x"55",
         11181 => x"08",
         11182 => x"90",
         11183 => x"fe",
         11184 => x"52",
         11185 => x"ac",
         11186 => x"bb",
         11187 => x"84",
         11188 => x"fc",
         11189 => x"39",
         11190 => x"19",
         11191 => x"19",
         11192 => x"33",
         11193 => x"c2",
         11194 => x"84",
         11195 => x"90",
         11196 => x"ff",
         11197 => x"90",
         11198 => x"58",
         11199 => x"81",
         11200 => x"ff",
         11201 => x"84",
         11202 => x"81",
         11203 => x"fb",
         11204 => x"79",
         11205 => x"fb",
         11206 => x"0b",
         11207 => x"81",
         11208 => x"84",
         11209 => x"0d",
         11210 => x"91",
         11211 => x"0b",
         11212 => x"0c",
         11213 => x"04",
         11214 => x"7d",
         11215 => x"77",
         11216 => x"38",
         11217 => x"75",
         11218 => x"38",
         11219 => x"74",
         11220 => x"38",
         11221 => x"84",
         11222 => x"5a",
         11223 => x"83",
         11224 => x"55",
         11225 => x"56",
         11226 => x"38",
         11227 => x"70",
         11228 => x"06",
         11229 => x"80",
         11230 => x"38",
         11231 => x"56",
         11232 => x"83",
         11233 => x"a0",
         11234 => x"56",
         11235 => x"77",
         11236 => x"80",
         11237 => x"33",
         11238 => x"5a",
         11239 => x"09",
         11240 => x"c0",
         11241 => x"76",
         11242 => x"52",
         11243 => x"51",
         11244 => x"3f",
         11245 => x"08",
         11246 => x"38",
         11247 => x"59",
         11248 => x"0c",
         11249 => x"81",
         11250 => x"18",
         11251 => x"33",
         11252 => x"57",
         11253 => x"34",
         11254 => x"19",
         11255 => x"ff",
         11256 => x"5a",
         11257 => x"18",
         11258 => x"2a",
         11259 => x"18",
         11260 => x"76",
         11261 => x"5c",
         11262 => x"83",
         11263 => x"38",
         11264 => x"55",
         11265 => x"74",
         11266 => x"7a",
         11267 => x"74",
         11268 => x"75",
         11269 => x"74",
         11270 => x"78",
         11271 => x"80",
         11272 => x"0b",
         11273 => x"a1",
         11274 => x"34",
         11275 => x"99",
         11276 => x"0b",
         11277 => x"80",
         11278 => x"34",
         11279 => x"0b",
         11280 => x"7b",
         11281 => x"95",
         11282 => x"84",
         11283 => x"33",
         11284 => x"5b",
         11285 => x"19",
         11286 => x"74",
         11287 => x"0c",
         11288 => x"04",
         11289 => x"16",
         11290 => x"16",
         11291 => x"17",
         11292 => x"ff",
         11293 => x"81",
         11294 => x"84",
         11295 => x"09",
         11296 => x"c0",
         11297 => x"84",
         11298 => x"34",
         11299 => x"a8",
         11300 => x"84",
         11301 => x"5a",
         11302 => x"17",
         11303 => x"85",
         11304 => x"33",
         11305 => x"2e",
         11306 => x"fd",
         11307 => x"54",
         11308 => x"a0",
         11309 => x"53",
         11310 => x"16",
         11311 => x"94",
         11312 => x"59",
         11313 => x"78",
         11314 => x"74",
         11315 => x"74",
         11316 => x"75",
         11317 => x"8c",
         11318 => x"74",
         11319 => x"88",
         11320 => x"9d",
         11321 => x"90",
         11322 => x"9e",
         11323 => x"98",
         11324 => x"9f",
         11325 => x"7a",
         11326 => x"97",
         11327 => x"0b",
         11328 => x"80",
         11329 => x"18",
         11330 => x"92",
         11331 => x"0b",
         11332 => x"7b",
         11333 => x"83",
         11334 => x"51",
         11335 => x"3f",
         11336 => x"08",
         11337 => x"81",
         11338 => x"56",
         11339 => x"34",
         11340 => x"81",
         11341 => x"ff",
         11342 => x"84",
         11343 => x"81",
         11344 => x"fc",
         11345 => x"78",
         11346 => x"fc",
         11347 => x"54",
         11348 => x"53",
         11349 => x"7b",
         11350 => x"52",
         11351 => x"ca",
         11352 => x"84",
         11353 => x"fd",
         11354 => x"18",
         11355 => x"06",
         11356 => x"19",
         11357 => x"19",
         11358 => x"b4",
         11359 => x"2e",
         11360 => x"fc",
         11361 => x"c2",
         11362 => x"0d",
         11363 => x"55",
         11364 => x"84",
         11365 => x"54",
         11366 => x"08",
         11367 => x"56",
         11368 => x"9e",
         11369 => x"53",
         11370 => x"96",
         11371 => x"52",
         11372 => x"8e",
         11373 => x"22",
         11374 => x"58",
         11375 => x"2e",
         11376 => x"52",
         11377 => x"54",
         11378 => x"75",
         11379 => x"84",
         11380 => x"89",
         11381 => x"81",
         11382 => x"ff",
         11383 => x"84",
         11384 => x"81",
         11385 => x"da",
         11386 => x"08",
         11387 => x"39",
         11388 => x"ff",
         11389 => x"57",
         11390 => x"2e",
         11391 => x"70",
         11392 => x"33",
         11393 => x"52",
         11394 => x"2e",
         11395 => x"ee",
         11396 => x"2e",
         11397 => x"e2",
         11398 => x"80",
         11399 => x"38",
         11400 => x"e0",
         11401 => x"84",
         11402 => x"8c",
         11403 => x"8b",
         11404 => x"84",
         11405 => x"0d",
         11406 => x"d0",
         11407 => x"ff",
         11408 => x"53",
         11409 => x"91",
         11410 => x"73",
         11411 => x"d0",
         11412 => x"73",
         11413 => x"f5",
         11414 => x"83",
         11415 => x"58",
         11416 => x"56",
         11417 => x"81",
         11418 => x"75",
         11419 => x"57",
         11420 => x"12",
         11421 => x"70",
         11422 => x"38",
         11423 => x"81",
         11424 => x"54",
         11425 => x"51",
         11426 => x"89",
         11427 => x"70",
         11428 => x"54",
         11429 => x"70",
         11430 => x"51",
         11431 => x"09",
         11432 => x"38",
         11433 => x"38",
         11434 => x"70",
         11435 => x"07",
         11436 => x"07",
         11437 => x"76",
         11438 => x"38",
         11439 => x"1b",
         11440 => x"78",
         11441 => x"38",
         11442 => x"cf",
         11443 => x"24",
         11444 => x"76",
         11445 => x"c3",
         11446 => x"0d",
         11447 => x"3d",
         11448 => x"99",
         11449 => x"d3",
         11450 => x"84",
         11451 => x"bb",
         11452 => x"2e",
         11453 => x"84",
         11454 => x"98",
         11455 => x"7a",
         11456 => x"98",
         11457 => x"51",
         11458 => x"84",
         11459 => x"55",
         11460 => x"08",
         11461 => x"02",
         11462 => x"33",
         11463 => x"58",
         11464 => x"24",
         11465 => x"02",
         11466 => x"70",
         11467 => x"06",
         11468 => x"80",
         11469 => x"7a",
         11470 => x"33",
         11471 => x"71",
         11472 => x"73",
         11473 => x"5b",
         11474 => x"83",
         11475 => x"76",
         11476 => x"74",
         11477 => x"0c",
         11478 => x"04",
         11479 => x"08",
         11480 => x"81",
         11481 => x"38",
         11482 => x"bb",
         11483 => x"3d",
         11484 => x"16",
         11485 => x"33",
         11486 => x"71",
         11487 => x"79",
         11488 => x"0c",
         11489 => x"39",
         11490 => x"12",
         11491 => x"84",
         11492 => x"98",
         11493 => x"ff",
         11494 => x"80",
         11495 => x"80",
         11496 => x"5d",
         11497 => x"34",
         11498 => x"e4",
         11499 => x"05",
         11500 => x"3d",
         11501 => x"3f",
         11502 => x"08",
         11503 => x"84",
         11504 => x"38",
         11505 => x"3d",
         11506 => x"98",
         11507 => x"dd",
         11508 => x"80",
         11509 => x"5b",
         11510 => x"2e",
         11511 => x"80",
         11512 => x"3d",
         11513 => x"52",
         11514 => x"a5",
         11515 => x"bb",
         11516 => x"84",
         11517 => x"83",
         11518 => x"80",
         11519 => x"58",
         11520 => x"08",
         11521 => x"38",
         11522 => x"08",
         11523 => x"5f",
         11524 => x"c7",
         11525 => x"76",
         11526 => x"52",
         11527 => x"51",
         11528 => x"3f",
         11529 => x"08",
         11530 => x"38",
         11531 => x"59",
         11532 => x"0c",
         11533 => x"38",
         11534 => x"08",
         11535 => x"9a",
         11536 => x"88",
         11537 => x"70",
         11538 => x"59",
         11539 => x"83",
         11540 => x"38",
         11541 => x"3d",
         11542 => x"7a",
         11543 => x"f6",
         11544 => x"84",
         11545 => x"bb",
         11546 => x"9f",
         11547 => x"7a",
         11548 => x"b4",
         11549 => x"84",
         11550 => x"bb",
         11551 => x"38",
         11552 => x"08",
         11553 => x"9a",
         11554 => x"88",
         11555 => x"70",
         11556 => x"59",
         11557 => x"83",
         11558 => x"38",
         11559 => x"a4",
         11560 => x"84",
         11561 => x"51",
         11562 => x"3f",
         11563 => x"08",
         11564 => x"84",
         11565 => x"ff",
         11566 => x"84",
         11567 => x"38",
         11568 => x"38",
         11569 => x"fd",
         11570 => x"7a",
         11571 => x"c8",
         11572 => x"82",
         11573 => x"57",
         11574 => x"90",
         11575 => x"56",
         11576 => x"17",
         11577 => x"57",
         11578 => x"38",
         11579 => x"75",
         11580 => x"95",
         11581 => x"2e",
         11582 => x"17",
         11583 => x"ff",
         11584 => x"3d",
         11585 => x"19",
         11586 => x"59",
         11587 => x"33",
         11588 => x"eb",
         11589 => x"80",
         11590 => x"11",
         11591 => x"7e",
         11592 => x"3d",
         11593 => x"fd",
         11594 => x"60",
         11595 => x"38",
         11596 => x"e2",
         11597 => x"10",
         11598 => x"f4",
         11599 => x"70",
         11600 => x"59",
         11601 => x"7a",
         11602 => x"81",
         11603 => x"70",
         11604 => x"5a",
         11605 => x"82",
         11606 => x"78",
         11607 => x"80",
         11608 => x"27",
         11609 => x"16",
         11610 => x"7c",
         11611 => x"5e",
         11612 => x"57",
         11613 => x"ee",
         11614 => x"70",
         11615 => x"34",
         11616 => x"09",
         11617 => x"df",
         11618 => x"80",
         11619 => x"84",
         11620 => x"80",
         11621 => x"04",
         11622 => x"94",
         11623 => x"98",
         11624 => x"2b",
         11625 => x"59",
         11626 => x"f0",
         11627 => x"33",
         11628 => x"71",
         11629 => x"90",
         11630 => x"07",
         11631 => x"0c",
         11632 => x"52",
         11633 => x"a2",
         11634 => x"bb",
         11635 => x"84",
         11636 => x"80",
         11637 => x"38",
         11638 => x"81",
         11639 => x"08",
         11640 => x"70",
         11641 => x"33",
         11642 => x"8a",
         11643 => x"59",
         11644 => x"08",
         11645 => x"84",
         11646 => x"83",
         11647 => x"16",
         11648 => x"08",
         11649 => x"84",
         11650 => x"74",
         11651 => x"27",
         11652 => x"82",
         11653 => x"74",
         11654 => x"81",
         11655 => x"38",
         11656 => x"16",
         11657 => x"08",
         11658 => x"52",
         11659 => x"51",
         11660 => x"3f",
         11661 => x"dd",
         11662 => x"80",
         11663 => x"11",
         11664 => x"7b",
         11665 => x"84",
         11666 => x"70",
         11667 => x"e6",
         11668 => x"08",
         11669 => x"59",
         11670 => x"7e",
         11671 => x"81",
         11672 => x"38",
         11673 => x"80",
         11674 => x"18",
         11675 => x"5a",
         11676 => x"70",
         11677 => x"34",
         11678 => x"fe",
         11679 => x"e5",
         11680 => x"81",
         11681 => x"79",
         11682 => x"81",
         11683 => x"7f",
         11684 => x"38",
         11685 => x"82",
         11686 => x"34",
         11687 => x"84",
         11688 => x"3d",
         11689 => x"3d",
         11690 => x"5a",
         11691 => x"76",
         11692 => x"38",
         11693 => x"75",
         11694 => x"38",
         11695 => x"74",
         11696 => x"38",
         11697 => x"84",
         11698 => x"5b",
         11699 => x"83",
         11700 => x"55",
         11701 => x"55",
         11702 => x"38",
         11703 => x"55",
         11704 => x"38",
         11705 => x"58",
         11706 => x"82",
         11707 => x"17",
         11708 => x"5a",
         11709 => x"83",
         11710 => x"8a",
         11711 => x"89",
         11712 => x"58",
         11713 => x"82",
         11714 => x"52",
         11715 => x"fd",
         11716 => x"84",
         11717 => x"ff",
         11718 => x"70",
         11719 => x"fd",
         11720 => x"84",
         11721 => x"75",
         11722 => x"38",
         11723 => x"06",
         11724 => x"0c",
         11725 => x"98",
         11726 => x"5a",
         11727 => x"2e",
         11728 => x"77",
         11729 => x"d3",
         11730 => x"31",
         11731 => x"19",
         11732 => x"90",
         11733 => x"81",
         11734 => x"51",
         11735 => x"80",
         11736 => x"38",
         11737 => x"51",
         11738 => x"3f",
         11739 => x"08",
         11740 => x"84",
         11741 => x"9e",
         11742 => x"2e",
         11743 => x"81",
         11744 => x"82",
         11745 => x"75",
         11746 => x"27",
         11747 => x"75",
         11748 => x"ff",
         11749 => x"bb",
         11750 => x"94",
         11751 => x"94",
         11752 => x"83",
         11753 => x"77",
         11754 => x"38",
         11755 => x"9c",
         11756 => x"05",
         11757 => x"75",
         11758 => x"ca",
         11759 => x"22",
         11760 => x"b0",
         11761 => x"7a",
         11762 => x"5c",
         11763 => x"80",
         11764 => x"38",
         11765 => x"58",
         11766 => x"56",
         11767 => x"90",
         11768 => x"18",
         11769 => x"33",
         11770 => x"59",
         11771 => x"34",
         11772 => x"06",
         11773 => x"2e",
         11774 => x"9c",
         11775 => x"75",
         11776 => x"a1",
         11777 => x"33",
         11778 => x"a8",
         11779 => x"59",
         11780 => x"a2",
         11781 => x"75",
         11782 => x"7b",
         11783 => x"52",
         11784 => x"86",
         11785 => x"84",
         11786 => x"90",
         11787 => x"ff",
         11788 => x"90",
         11789 => x"54",
         11790 => x"52",
         11791 => x"33",
         11792 => x"84",
         11793 => x"bb",
         11794 => x"2e",
         11795 => x"81",
         11796 => x"34",
         11797 => x"84",
         11798 => x"8d",
         11799 => x"90",
         11800 => x"81",
         11801 => x"57",
         11802 => x"82",
         11803 => x"18",
         11804 => x"80",
         11805 => x"2e",
         11806 => x"fc",
         11807 => x"94",
         11808 => x"d4",
         11809 => x"94",
         11810 => x"17",
         11811 => x"80",
         11812 => x"38",
         11813 => x"0c",
         11814 => x"fe",
         11815 => x"a3",
         11816 => x"18",
         11817 => x"84",
         11818 => x"8d",
         11819 => x"75",
         11820 => x"ff",
         11821 => x"84",
         11822 => x"56",
         11823 => x"81",
         11824 => x"ff",
         11825 => x"84",
         11826 => x"81",
         11827 => x"fc",
         11828 => x"77",
         11829 => x"fb",
         11830 => x"52",
         11831 => x"98",
         11832 => x"bb",
         11833 => x"84",
         11834 => x"81",
         11835 => x"84",
         11836 => x"ff",
         11837 => x"38",
         11838 => x"08",
         11839 => x"75",
         11840 => x"ff",
         11841 => x"0b",
         11842 => x"82",
         11843 => x"84",
         11844 => x"0d",
         11845 => x"0d",
         11846 => x"54",
         11847 => x"a2",
         11848 => x"8c",
         11849 => x"52",
         11850 => x"05",
         11851 => x"3f",
         11852 => x"08",
         11853 => x"84",
         11854 => x"8f",
         11855 => x"0c",
         11856 => x"84",
         11857 => x"8c",
         11858 => x"7a",
         11859 => x"52",
         11860 => x"ba",
         11861 => x"bb",
         11862 => x"84",
         11863 => x"80",
         11864 => x"16",
         11865 => x"2b",
         11866 => x"78",
         11867 => x"86",
         11868 => x"84",
         11869 => x"5b",
         11870 => x"2e",
         11871 => x"9c",
         11872 => x"11",
         11873 => x"33",
         11874 => x"07",
         11875 => x"5d",
         11876 => x"57",
         11877 => x"b3",
         11878 => x"17",
         11879 => x"86",
         11880 => x"17",
         11881 => x"75",
         11882 => x"aa",
         11883 => x"84",
         11884 => x"84",
         11885 => x"74",
         11886 => x"84",
         11887 => x"0c",
         11888 => x"85",
         11889 => x"0c",
         11890 => x"95",
         11891 => x"18",
         11892 => x"2b",
         11893 => x"07",
         11894 => x"19",
         11895 => x"ff",
         11896 => x"3d",
         11897 => x"89",
         11898 => x"2e",
         11899 => x"08",
         11900 => x"2e",
         11901 => x"33",
         11902 => x"2e",
         11903 => x"13",
         11904 => x"22",
         11905 => x"76",
         11906 => x"80",
         11907 => x"73",
         11908 => x"75",
         11909 => x"bb",
         11910 => x"3d",
         11911 => x"13",
         11912 => x"80",
         11913 => x"bb",
         11914 => x"06",
         11915 => x"38",
         11916 => x"53",
         11917 => x"f8",
         11918 => x"7c",
         11919 => x"56",
         11920 => x"9f",
         11921 => x"54",
         11922 => x"97",
         11923 => x"53",
         11924 => x"8f",
         11925 => x"22",
         11926 => x"59",
         11927 => x"2e",
         11928 => x"80",
         11929 => x"75",
         11930 => x"c7",
         11931 => x"2e",
         11932 => x"75",
         11933 => x"ff",
         11934 => x"84",
         11935 => x"53",
         11936 => x"08",
         11937 => x"38",
         11938 => x"08",
         11939 => x"52",
         11940 => x"b3",
         11941 => x"52",
         11942 => x"9a",
         11943 => x"bb",
         11944 => x"32",
         11945 => x"72",
         11946 => x"84",
         11947 => x"06",
         11948 => x"72",
         11949 => x"0c",
         11950 => x"04",
         11951 => x"75",
         11952 => x"b2",
         11953 => x"52",
         11954 => x"99",
         11955 => x"bb",
         11956 => x"32",
         11957 => x"72",
         11958 => x"84",
         11959 => x"06",
         11960 => x"cf",
         11961 => x"74",
         11962 => x"ea",
         11963 => x"84",
         11964 => x"84",
         11965 => x"0d",
         11966 => x"33",
         11967 => x"d9",
         11968 => x"84",
         11969 => x"53",
         11970 => x"38",
         11971 => x"54",
         11972 => x"39",
         11973 => x"66",
         11974 => x"89",
         11975 => x"97",
         11976 => x"c2",
         11977 => x"bb",
         11978 => x"84",
         11979 => x"80",
         11980 => x"74",
         11981 => x"0c",
         11982 => x"04",
         11983 => x"51",
         11984 => x"3f",
         11985 => x"08",
         11986 => x"84",
         11987 => x"02",
         11988 => x"33",
         11989 => x"55",
         11990 => x"24",
         11991 => x"80",
         11992 => x"76",
         11993 => x"ff",
         11994 => x"74",
         11995 => x"0c",
         11996 => x"04",
         11997 => x"bb",
         11998 => x"3d",
         11999 => x"3d",
         12000 => x"56",
         12001 => x"95",
         12002 => x"52",
         12003 => x"c1",
         12004 => x"bb",
         12005 => x"84",
         12006 => x"9a",
         12007 => x"0c",
         12008 => x"11",
         12009 => x"94",
         12010 => x"57",
         12011 => x"75",
         12012 => x"75",
         12013 => x"84",
         12014 => x"95",
         12015 => x"84",
         12016 => x"77",
         12017 => x"78",
         12018 => x"93",
         12019 => x"18",
         12020 => x"84",
         12021 => x"59",
         12022 => x"38",
         12023 => x"71",
         12024 => x"b4",
         12025 => x"2e",
         12026 => x"83",
         12027 => x"5f",
         12028 => x"8d",
         12029 => x"75",
         12030 => x"52",
         12031 => x"51",
         12032 => x"3f",
         12033 => x"08",
         12034 => x"38",
         12035 => x"5e",
         12036 => x"0c",
         12037 => x"57",
         12038 => x"38",
         12039 => x"7d",
         12040 => x"8d",
         12041 => x"b8",
         12042 => x"33",
         12043 => x"71",
         12044 => x"88",
         12045 => x"14",
         12046 => x"07",
         12047 => x"33",
         12048 => x"ff",
         12049 => x"07",
         12050 => x"80",
         12051 => x"60",
         12052 => x"ff",
         12053 => x"05",
         12054 => x"53",
         12055 => x"58",
         12056 => x"78",
         12057 => x"7a",
         12058 => x"94",
         12059 => x"17",
         12060 => x"58",
         12061 => x"34",
         12062 => x"84",
         12063 => x"0d",
         12064 => x"b4",
         12065 => x"b8",
         12066 => x"81",
         12067 => x"5d",
         12068 => x"3f",
         12069 => x"bb",
         12070 => x"f8",
         12071 => x"84",
         12072 => x"34",
         12073 => x"a8",
         12074 => x"84",
         12075 => x"5f",
         12076 => x"18",
         12077 => x"bd",
         12078 => x"33",
         12079 => x"2e",
         12080 => x"fe",
         12081 => x"54",
         12082 => x"a0",
         12083 => x"53",
         12084 => x"17",
         12085 => x"fc",
         12086 => x"5e",
         12087 => x"82",
         12088 => x"3d",
         12089 => x"52",
         12090 => x"81",
         12091 => x"bb",
         12092 => x"2e",
         12093 => x"84",
         12094 => x"81",
         12095 => x"38",
         12096 => x"08",
         12097 => x"bb",
         12098 => x"80",
         12099 => x"81",
         12100 => x"58",
         12101 => x"17",
         12102 => x"ca",
         12103 => x"0c",
         12104 => x"0c",
         12105 => x"81",
         12106 => x"84",
         12107 => x"c8",
         12108 => x"b8",
         12109 => x"33",
         12110 => x"88",
         12111 => x"30",
         12112 => x"1f",
         12113 => x"ff",
         12114 => x"5f",
         12115 => x"5f",
         12116 => x"fd",
         12117 => x"8f",
         12118 => x"fd",
         12119 => x"60",
         12120 => x"7f",
         12121 => x"18",
         12122 => x"33",
         12123 => x"77",
         12124 => x"fe",
         12125 => x"60",
         12126 => x"39",
         12127 => x"7c",
         12128 => x"77",
         12129 => x"38",
         12130 => x"75",
         12131 => x"38",
         12132 => x"74",
         12133 => x"38",
         12134 => x"84",
         12135 => x"5a",
         12136 => x"82",
         12137 => x"55",
         12138 => x"81",
         12139 => x"18",
         12140 => x"80",
         12141 => x"18",
         12142 => x"2a",
         12143 => x"59",
         12144 => x"80",
         12145 => x"38",
         12146 => x"55",
         12147 => x"08",
         12148 => x"38",
         12149 => x"38",
         12150 => x"78",
         12151 => x"81",
         12152 => x"38",
         12153 => x"75",
         12154 => x"38",
         12155 => x"0b",
         12156 => x"94",
         12157 => x"19",
         12158 => x"c0",
         12159 => x"90",
         12160 => x"a8",
         12161 => x"2b",
         12162 => x"25",
         12163 => x"54",
         12164 => x"53",
         12165 => x"7a",
         12166 => x"52",
         12167 => x"8a",
         12168 => x"84",
         12169 => x"83",
         12170 => x"57",
         12171 => x"34",
         12172 => x"84",
         12173 => x"8c",
         12174 => x"79",
         12175 => x"27",
         12176 => x"74",
         12177 => x"fe",
         12178 => x"84",
         12179 => x"5a",
         12180 => x"08",
         12181 => x"e9",
         12182 => x"84",
         12183 => x"82",
         12184 => x"bb",
         12185 => x"2e",
         12186 => x"80",
         12187 => x"76",
         12188 => x"cb",
         12189 => x"84",
         12190 => x"38",
         12191 => x"fe",
         12192 => x"08",
         12193 => x"75",
         12194 => x"af",
         12195 => x"94",
         12196 => x"17",
         12197 => x"55",
         12198 => x"34",
         12199 => x"7a",
         12200 => x"38",
         12201 => x"16",
         12202 => x"f7",
         12203 => x"bb",
         12204 => x"06",
         12205 => x"ee",
         12206 => x"08",
         12207 => x"e8",
         12208 => x"90",
         12209 => x"55",
         12210 => x"0b",
         12211 => x"fe",
         12212 => x"18",
         12213 => x"51",
         12214 => x"3f",
         12215 => x"08",
         12216 => x"c2",
         12217 => x"84",
         12218 => x"81",
         12219 => x"81",
         12220 => x"59",
         12221 => x"08",
         12222 => x"27",
         12223 => x"84",
         12224 => x"98",
         12225 => x"08",
         12226 => x"81",
         12227 => x"84",
         12228 => x"a1",
         12229 => x"84",
         12230 => x"08",
         12231 => x"38",
         12232 => x"97",
         12233 => x"75",
         12234 => x"ff",
         12235 => x"84",
         12236 => x"56",
         12237 => x"08",
         12238 => x"74",
         12239 => x"fe",
         12240 => x"84",
         12241 => x"5a",
         12242 => x"08",
         12243 => x"cb",
         12244 => x"84",
         12245 => x"80",
         12246 => x"bb",
         12247 => x"2e",
         12248 => x"80",
         12249 => x"76",
         12250 => x"d3",
         12251 => x"84",
         12252 => x"38",
         12253 => x"fe",
         12254 => x"08",
         12255 => x"75",
         12256 => x"38",
         12257 => x"18",
         12258 => x"33",
         12259 => x"74",
         12260 => x"79",
         12261 => x"26",
         12262 => x"80",
         12263 => x"90",
         12264 => x"fc",
         12265 => x"57",
         12266 => x"82",
         12267 => x"33",
         12268 => x"bf",
         12269 => x"e7",
         12270 => x"33",
         12271 => x"55",
         12272 => x"34",
         12273 => x"ea",
         12274 => x"90",
         12275 => x"55",
         12276 => x"84",
         12277 => x"90",
         12278 => x"55",
         12279 => x"81",
         12280 => x"33",
         12281 => x"e0",
         12282 => x"84",
         12283 => x"af",
         12284 => x"ff",
         12285 => x"3d",
         12286 => x"a7",
         12287 => x"05",
         12288 => x"51",
         12289 => x"3f",
         12290 => x"08",
         12291 => x"84",
         12292 => x"8a",
         12293 => x"bb",
         12294 => x"3d",
         12295 => x"4b",
         12296 => x"52",
         12297 => x"52",
         12298 => x"b1",
         12299 => x"84",
         12300 => x"bb",
         12301 => x"38",
         12302 => x"05",
         12303 => x"2a",
         12304 => x"57",
         12305 => x"cd",
         12306 => x"2b",
         12307 => x"24",
         12308 => x"80",
         12309 => x"70",
         12310 => x"57",
         12311 => x"ff",
         12312 => x"a3",
         12313 => x"11",
         12314 => x"33",
         12315 => x"07",
         12316 => x"5e",
         12317 => x"7c",
         12318 => x"d5",
         12319 => x"2a",
         12320 => x"76",
         12321 => x"ed",
         12322 => x"98",
         12323 => x"2e",
         12324 => x"77",
         12325 => x"84",
         12326 => x"52",
         12327 => x"52",
         12328 => x"b2",
         12329 => x"84",
         12330 => x"bb",
         12331 => x"e5",
         12332 => x"84",
         12333 => x"51",
         12334 => x"3f",
         12335 => x"08",
         12336 => x"84",
         12337 => x"87",
         12338 => x"84",
         12339 => x"0d",
         12340 => x"33",
         12341 => x"71",
         12342 => x"90",
         12343 => x"07",
         12344 => x"ff",
         12345 => x"bb",
         12346 => x"2e",
         12347 => x"bb",
         12348 => x"a1",
         12349 => x"6f",
         12350 => x"57",
         12351 => x"ff",
         12352 => x"38",
         12353 => x"51",
         12354 => x"3f",
         12355 => x"08",
         12356 => x"84",
         12357 => x"be",
         12358 => x"70",
         12359 => x"25",
         12360 => x"80",
         12361 => x"74",
         12362 => x"38",
         12363 => x"58",
         12364 => x"27",
         12365 => x"17",
         12366 => x"81",
         12367 => x"56",
         12368 => x"38",
         12369 => x"f6",
         12370 => x"bb",
         12371 => x"bb",
         12372 => x"3d",
         12373 => x"17",
         12374 => x"08",
         12375 => x"b4",
         12376 => x"2e",
         12377 => x"83",
         12378 => x"59",
         12379 => x"2e",
         12380 => x"80",
         12381 => x"54",
         12382 => x"17",
         12383 => x"33",
         12384 => x"a7",
         12385 => x"84",
         12386 => x"85",
         12387 => x"81",
         12388 => x"18",
         12389 => x"77",
         12390 => x"19",
         12391 => x"78",
         12392 => x"83",
         12393 => x"19",
         12394 => x"fe",
         12395 => x"52",
         12396 => x"8c",
         12397 => x"bb",
         12398 => x"84",
         12399 => x"80",
         12400 => x"38",
         12401 => x"09",
         12402 => x"cd",
         12403 => x"fe",
         12404 => x"54",
         12405 => x"53",
         12406 => x"17",
         12407 => x"f2",
         12408 => x"58",
         12409 => x"08",
         12410 => x"81",
         12411 => x"38",
         12412 => x"08",
         12413 => x"b4",
         12414 => x"18",
         12415 => x"bb",
         12416 => x"55",
         12417 => x"08",
         12418 => x"38",
         12419 => x"55",
         12420 => x"09",
         12421 => x"de",
         12422 => x"b4",
         12423 => x"18",
         12424 => x"7c",
         12425 => x"33",
         12426 => x"fe",
         12427 => x"fe",
         12428 => x"55",
         12429 => x"80",
         12430 => x"52",
         12431 => x"f7",
         12432 => x"bb",
         12433 => x"84",
         12434 => x"80",
         12435 => x"38",
         12436 => x"08",
         12437 => x"e6",
         12438 => x"84",
         12439 => x"80",
         12440 => x"53",
         12441 => x"51",
         12442 => x"3f",
         12443 => x"08",
         12444 => x"17",
         12445 => x"94",
         12446 => x"5c",
         12447 => x"27",
         12448 => x"81",
         12449 => x"0c",
         12450 => x"81",
         12451 => x"84",
         12452 => x"55",
         12453 => x"ff",
         12454 => x"56",
         12455 => x"79",
         12456 => x"39",
         12457 => x"08",
         12458 => x"39",
         12459 => x"90",
         12460 => x"0d",
         12461 => x"3d",
         12462 => x"52",
         12463 => x"ff",
         12464 => x"84",
         12465 => x"56",
         12466 => x"08",
         12467 => x"38",
         12468 => x"84",
         12469 => x"0d",
         12470 => x"6f",
         12471 => x"70",
         12472 => x"a6",
         12473 => x"bb",
         12474 => x"84",
         12475 => x"8b",
         12476 => x"84",
         12477 => x"9f",
         12478 => x"84",
         12479 => x"84",
         12480 => x"06",
         12481 => x"80",
         12482 => x"70",
         12483 => x"06",
         12484 => x"56",
         12485 => x"38",
         12486 => x"52",
         12487 => x"52",
         12488 => x"f9",
         12489 => x"84",
         12490 => x"5c",
         12491 => x"08",
         12492 => x"56",
         12493 => x"08",
         12494 => x"f9",
         12495 => x"84",
         12496 => x"81",
         12497 => x"81",
         12498 => x"84",
         12499 => x"83",
         12500 => x"5a",
         12501 => x"e2",
         12502 => x"9c",
         12503 => x"05",
         12504 => x"5b",
         12505 => x"8d",
         12506 => x"22",
         12507 => x"b0",
         12508 => x"5c",
         12509 => x"18",
         12510 => x"59",
         12511 => x"57",
         12512 => x"70",
         12513 => x"34",
         12514 => x"74",
         12515 => x"58",
         12516 => x"55",
         12517 => x"81",
         12518 => x"54",
         12519 => x"78",
         12520 => x"33",
         12521 => x"82",
         12522 => x"84",
         12523 => x"38",
         12524 => x"dc",
         12525 => x"ff",
         12526 => x"54",
         12527 => x"53",
         12528 => x"53",
         12529 => x"52",
         12530 => x"de",
         12531 => x"84",
         12532 => x"be",
         12533 => x"84",
         12534 => x"34",
         12535 => x"a8",
         12536 => x"55",
         12537 => x"08",
         12538 => x"38",
         12539 => x"5b",
         12540 => x"09",
         12541 => x"e1",
         12542 => x"b4",
         12543 => x"18",
         12544 => x"77",
         12545 => x"33",
         12546 => x"9e",
         12547 => x"39",
         12548 => x"7d",
         12549 => x"81",
         12550 => x"b4",
         12551 => x"18",
         12552 => x"ac",
         12553 => x"7c",
         12554 => x"b2",
         12555 => x"84",
         12556 => x"bb",
         12557 => x"2e",
         12558 => x"84",
         12559 => x"81",
         12560 => x"38",
         12561 => x"08",
         12562 => x"84",
         12563 => x"74",
         12564 => x"fe",
         12565 => x"84",
         12566 => x"fc",
         12567 => x"17",
         12568 => x"94",
         12569 => x"5c",
         12570 => x"27",
         12571 => x"18",
         12572 => x"84",
         12573 => x"07",
         12574 => x"18",
         12575 => x"78",
         12576 => x"a1",
         12577 => x"bb",
         12578 => x"3d",
         12579 => x"17",
         12580 => x"83",
         12581 => x"57",
         12582 => x"78",
         12583 => x"06",
         12584 => x"8b",
         12585 => x"56",
         12586 => x"70",
         12587 => x"34",
         12588 => x"75",
         12589 => x"57",
         12590 => x"18",
         12591 => x"90",
         12592 => x"19",
         12593 => x"75",
         12594 => x"34",
         12595 => x"1a",
         12596 => x"80",
         12597 => x"80",
         12598 => x"d1",
         12599 => x"7c",
         12600 => x"06",
         12601 => x"80",
         12602 => x"77",
         12603 => x"7a",
         12604 => x"34",
         12605 => x"74",
         12606 => x"cc",
         12607 => x"a0",
         12608 => x"1a",
         12609 => x"58",
         12610 => x"81",
         12611 => x"77",
         12612 => x"59",
         12613 => x"56",
         12614 => x"7d",
         12615 => x"80",
         12616 => x"64",
         12617 => x"ff",
         12618 => x"57",
         12619 => x"f2",
         12620 => x"88",
         12621 => x"80",
         12622 => x"75",
         12623 => x"83",
         12624 => x"38",
         12625 => x"0b",
         12626 => x"79",
         12627 => x"cf",
         12628 => x"84",
         12629 => x"bb",
         12630 => x"b6",
         12631 => x"84",
         12632 => x"96",
         12633 => x"bb",
         12634 => x"17",
         12635 => x"98",
         12636 => x"cc",
         12637 => x"34",
         12638 => x"5d",
         12639 => x"34",
         12640 => x"59",
         12641 => x"34",
         12642 => x"79",
         12643 => x"d9",
         12644 => x"90",
         12645 => x"34",
         12646 => x"0b",
         12647 => x"7d",
         12648 => x"b9",
         12649 => x"84",
         12650 => x"84",
         12651 => x"9f",
         12652 => x"76",
         12653 => x"74",
         12654 => x"34",
         12655 => x"57",
         12656 => x"17",
         12657 => x"39",
         12658 => x"5b",
         12659 => x"17",
         12660 => x"2a",
         12661 => x"cd",
         12662 => x"59",
         12663 => x"d8",
         12664 => x"57",
         12665 => x"a1",
         12666 => x"2a",
         12667 => x"18",
         12668 => x"2a",
         12669 => x"18",
         12670 => x"90",
         12671 => x"34",
         12672 => x"0b",
         12673 => x"7d",
         12674 => x"d1",
         12675 => x"84",
         12676 => x"96",
         12677 => x"0d",
         12678 => x"3d",
         12679 => x"5b",
         12680 => x"2e",
         12681 => x"70",
         12682 => x"33",
         12683 => x"56",
         12684 => x"2e",
         12685 => x"74",
         12686 => x"ba",
         12687 => x"38",
         12688 => x"3d",
         12689 => x"52",
         12690 => x"ff",
         12691 => x"84",
         12692 => x"56",
         12693 => x"08",
         12694 => x"38",
         12695 => x"84",
         12696 => x"0d",
         12697 => x"3d",
         12698 => x"08",
         12699 => x"70",
         12700 => x"9f",
         12701 => x"bb",
         12702 => x"84",
         12703 => x"dc",
         12704 => x"bb",
         12705 => x"a0",
         12706 => x"56",
         12707 => x"a0",
         12708 => x"ae",
         12709 => x"58",
         12710 => x"81",
         12711 => x"77",
         12712 => x"59",
         12713 => x"55",
         12714 => x"99",
         12715 => x"78",
         12716 => x"55",
         12717 => x"05",
         12718 => x"70",
         12719 => x"34",
         12720 => x"74",
         12721 => x"3d",
         12722 => x"51",
         12723 => x"3f",
         12724 => x"08",
         12725 => x"84",
         12726 => x"38",
         12727 => x"08",
         12728 => x"38",
         12729 => x"bb",
         12730 => x"3d",
         12731 => x"33",
         12732 => x"81",
         12733 => x"57",
         12734 => x"26",
         12735 => x"17",
         12736 => x"06",
         12737 => x"59",
         12738 => x"80",
         12739 => x"7f",
         12740 => x"f4",
         12741 => x"5d",
         12742 => x"5c",
         12743 => x"05",
         12744 => x"70",
         12745 => x"33",
         12746 => x"5a",
         12747 => x"99",
         12748 => x"e0",
         12749 => x"ff",
         12750 => x"ff",
         12751 => x"77",
         12752 => x"38",
         12753 => x"81",
         12754 => x"55",
         12755 => x"9f",
         12756 => x"75",
         12757 => x"81",
         12758 => x"77",
         12759 => x"78",
         12760 => x"30",
         12761 => x"9f",
         12762 => x"5d",
         12763 => x"80",
         12764 => x"81",
         12765 => x"5e",
         12766 => x"24",
         12767 => x"7c",
         12768 => x"5b",
         12769 => x"7b",
         12770 => x"b4",
         12771 => x"0c",
         12772 => x"3d",
         12773 => x"52",
         12774 => x"ff",
         12775 => x"84",
         12776 => x"56",
         12777 => x"08",
         12778 => x"fd",
         12779 => x"aa",
         12780 => x"09",
         12781 => x"ac",
         12782 => x"ff",
         12783 => x"84",
         12784 => x"56",
         12785 => x"08",
         12786 => x"6f",
         12787 => x"8d",
         12788 => x"05",
         12789 => x"58",
         12790 => x"70",
         12791 => x"33",
         12792 => x"05",
         12793 => x"1a",
         12794 => x"38",
         12795 => x"05",
         12796 => x"34",
         12797 => x"70",
         12798 => x"06",
         12799 => x"89",
         12800 => x"07",
         12801 => x"19",
         12802 => x"81",
         12803 => x"34",
         12804 => x"70",
         12805 => x"06",
         12806 => x"80",
         12807 => x"38",
         12808 => x"6b",
         12809 => x"38",
         12810 => x"33",
         12811 => x"71",
         12812 => x"72",
         12813 => x"5c",
         12814 => x"2e",
         12815 => x"fe",
         12816 => x"08",
         12817 => x"56",
         12818 => x"82",
         12819 => x"17",
         12820 => x"29",
         12821 => x"05",
         12822 => x"80",
         12823 => x"38",
         12824 => x"58",
         12825 => x"76",
         12826 => x"83",
         12827 => x"7e",
         12828 => x"81",
         12829 => x"b8",
         12830 => x"17",
         12831 => x"e4",
         12832 => x"bb",
         12833 => x"2e",
         12834 => x"58",
         12835 => x"b4",
         12836 => x"57",
         12837 => x"18",
         12838 => x"fb",
         12839 => x"15",
         12840 => x"ae",
         12841 => x"06",
         12842 => x"70",
         12843 => x"06",
         12844 => x"80",
         12845 => x"7b",
         12846 => x"77",
         12847 => x"34",
         12848 => x"7a",
         12849 => x"81",
         12850 => x"75",
         12851 => x"7d",
         12852 => x"34",
         12853 => x"56",
         12854 => x"18",
         12855 => x"81",
         12856 => x"34",
         12857 => x"3d",
         12858 => x"08",
         12859 => x"74",
         12860 => x"38",
         12861 => x"51",
         12862 => x"3f",
         12863 => x"08",
         12864 => x"84",
         12865 => x"38",
         12866 => x"98",
         12867 => x"80",
         12868 => x"08",
         12869 => x"38",
         12870 => x"7a",
         12871 => x"7a",
         12872 => x"06",
         12873 => x"81",
         12874 => x"b8",
         12875 => x"16",
         12876 => x"e2",
         12877 => x"bb",
         12878 => x"2e",
         12879 => x"57",
         12880 => x"b4",
         12881 => x"55",
         12882 => x"9c",
         12883 => x"e5",
         12884 => x"0b",
         12885 => x"90",
         12886 => x"27",
         12887 => x"52",
         12888 => x"fc",
         12889 => x"bb",
         12890 => x"84",
         12891 => x"80",
         12892 => x"38",
         12893 => x"84",
         12894 => x"38",
         12895 => x"f9",
         12896 => x"51",
         12897 => x"3f",
         12898 => x"08",
         12899 => x"0c",
         12900 => x"04",
         12901 => x"bb",
         12902 => x"3d",
         12903 => x"18",
         12904 => x"33",
         12905 => x"71",
         12906 => x"78",
         12907 => x"5c",
         12908 => x"84",
         12909 => x"84",
         12910 => x"38",
         12911 => x"08",
         12912 => x"a0",
         12913 => x"bb",
         12914 => x"3d",
         12915 => x"54",
         12916 => x"53",
         12917 => x"16",
         12918 => x"e2",
         12919 => x"58",
         12920 => x"08",
         12921 => x"81",
         12922 => x"38",
         12923 => x"08",
         12924 => x"b4",
         12925 => x"17",
         12926 => x"bb",
         12927 => x"55",
         12928 => x"08",
         12929 => x"38",
         12930 => x"5d",
         12931 => x"09",
         12932 => x"93",
         12933 => x"b4",
         12934 => x"17",
         12935 => x"7b",
         12936 => x"33",
         12937 => x"82",
         12938 => x"fd",
         12939 => x"54",
         12940 => x"53",
         12941 => x"53",
         12942 => x"52",
         12943 => x"ea",
         12944 => x"84",
         12945 => x"fc",
         12946 => x"bb",
         12947 => x"18",
         12948 => x"08",
         12949 => x"31",
         12950 => x"08",
         12951 => x"a0",
         12952 => x"fc",
         12953 => x"17",
         12954 => x"82",
         12955 => x"06",
         12956 => x"81",
         12957 => x"08",
         12958 => x"05",
         12959 => x"81",
         12960 => x"fe",
         12961 => x"79",
         12962 => x"39",
         12963 => x"02",
         12964 => x"33",
         12965 => x"80",
         12966 => x"56",
         12967 => x"96",
         12968 => x"52",
         12969 => x"ff",
         12970 => x"84",
         12971 => x"56",
         12972 => x"08",
         12973 => x"38",
         12974 => x"84",
         12975 => x"0d",
         12976 => x"66",
         12977 => x"d0",
         12978 => x"97",
         12979 => x"bb",
         12980 => x"84",
         12981 => x"e0",
         12982 => x"cf",
         12983 => x"a0",
         12984 => x"56",
         12985 => x"74",
         12986 => x"71",
         12987 => x"33",
         12988 => x"74",
         12989 => x"56",
         12990 => x"8b",
         12991 => x"55",
         12992 => x"16",
         12993 => x"fe",
         12994 => x"84",
         12995 => x"84",
         12996 => x"96",
         12997 => x"ec",
         12998 => x"57",
         12999 => x"3d",
         13000 => x"97",
         13001 => x"a2",
         13002 => x"bb",
         13003 => x"84",
         13004 => x"80",
         13005 => x"74",
         13006 => x"0c",
         13007 => x"04",
         13008 => x"52",
         13009 => x"05",
         13010 => x"91",
         13011 => x"84",
         13012 => x"bb",
         13013 => x"38",
         13014 => x"05",
         13015 => x"06",
         13016 => x"75",
         13017 => x"84",
         13018 => x"19",
         13019 => x"2b",
         13020 => x"56",
         13021 => x"34",
         13022 => x"55",
         13023 => x"34",
         13024 => x"58",
         13025 => x"34",
         13026 => x"54",
         13027 => x"34",
         13028 => x"0b",
         13029 => x"78",
         13030 => x"c1",
         13031 => x"84",
         13032 => x"84",
         13033 => x"0d",
         13034 => x"0d",
         13035 => x"5b",
         13036 => x"3d",
         13037 => x"9b",
         13038 => x"a0",
         13039 => x"bb",
         13040 => x"bb",
         13041 => x"70",
         13042 => x"08",
         13043 => x"51",
         13044 => x"80",
         13045 => x"81",
         13046 => x"5a",
         13047 => x"a4",
         13048 => x"70",
         13049 => x"25",
         13050 => x"80",
         13051 => x"38",
         13052 => x"06",
         13053 => x"80",
         13054 => x"38",
         13055 => x"08",
         13056 => x"5a",
         13057 => x"77",
         13058 => x"38",
         13059 => x"7a",
         13060 => x"7a",
         13061 => x"06",
         13062 => x"81",
         13063 => x"b8",
         13064 => x"16",
         13065 => x"dd",
         13066 => x"bb",
         13067 => x"2e",
         13068 => x"57",
         13069 => x"b4",
         13070 => x"57",
         13071 => x"7c",
         13072 => x"58",
         13073 => x"74",
         13074 => x"38",
         13075 => x"74",
         13076 => x"38",
         13077 => x"18",
         13078 => x"11",
         13079 => x"33",
         13080 => x"71",
         13081 => x"81",
         13082 => x"72",
         13083 => x"75",
         13084 => x"62",
         13085 => x"5e",
         13086 => x"76",
         13087 => x"0c",
         13088 => x"04",
         13089 => x"40",
         13090 => x"3d",
         13091 => x"fe",
         13092 => x"84",
         13093 => x"57",
         13094 => x"08",
         13095 => x"8d",
         13096 => x"2e",
         13097 => x"fe",
         13098 => x"7b",
         13099 => x"fe",
         13100 => x"54",
         13101 => x"53",
         13102 => x"53",
         13103 => x"52",
         13104 => x"e6",
         13105 => x"84",
         13106 => x"7a",
         13107 => x"06",
         13108 => x"84",
         13109 => x"83",
         13110 => x"16",
         13111 => x"08",
         13112 => x"84",
         13113 => x"74",
         13114 => x"27",
         13115 => x"82",
         13116 => x"74",
         13117 => x"81",
         13118 => x"38",
         13119 => x"16",
         13120 => x"08",
         13121 => x"52",
         13122 => x"51",
         13123 => x"3f",
         13124 => x"54",
         13125 => x"16",
         13126 => x"33",
         13127 => x"8b",
         13128 => x"84",
         13129 => x"fe",
         13130 => x"86",
         13131 => x"74",
         13132 => x"f4",
         13133 => x"84",
         13134 => x"bb",
         13135 => x"e1",
         13136 => x"84",
         13137 => x"84",
         13138 => x"59",
         13139 => x"81",
         13140 => x"57",
         13141 => x"33",
         13142 => x"19",
         13143 => x"27",
         13144 => x"70",
         13145 => x"80",
         13146 => x"80",
         13147 => x"38",
         13148 => x"11",
         13149 => x"57",
         13150 => x"2e",
         13151 => x"e1",
         13152 => x"fd",
         13153 => x"3d",
         13154 => x"a1",
         13155 => x"05",
         13156 => x"51",
         13157 => x"3f",
         13158 => x"08",
         13159 => x"84",
         13160 => x"38",
         13161 => x"8b",
         13162 => x"a0",
         13163 => x"05",
         13164 => x"15",
         13165 => x"38",
         13166 => x"08",
         13167 => x"81",
         13168 => x"58",
         13169 => x"78",
         13170 => x"38",
         13171 => x"3d",
         13172 => x"81",
         13173 => x"18",
         13174 => x"81",
         13175 => x"7c",
         13176 => x"ff",
         13177 => x"ff",
         13178 => x"a1",
         13179 => x"b5",
         13180 => x"84",
         13181 => x"dc",
         13182 => x"84",
         13183 => x"ff",
         13184 => x"80",
         13185 => x"38",
         13186 => x"0b",
         13187 => x"33",
         13188 => x"06",
         13189 => x"78",
         13190 => x"d6",
         13191 => x"78",
         13192 => x"38",
         13193 => x"33",
         13194 => x"06",
         13195 => x"74",
         13196 => x"38",
         13197 => x"09",
         13198 => x"38",
         13199 => x"06",
         13200 => x"a3",
         13201 => x"77",
         13202 => x"38",
         13203 => x"81",
         13204 => x"ff",
         13205 => x"38",
         13206 => x"55",
         13207 => x"81",
         13208 => x"81",
         13209 => x"7b",
         13210 => x"5d",
         13211 => x"a3",
         13212 => x"33",
         13213 => x"06",
         13214 => x"5a",
         13215 => x"fe",
         13216 => x"3d",
         13217 => x"56",
         13218 => x"2e",
         13219 => x"80",
         13220 => x"02",
         13221 => x"79",
         13222 => x"5c",
         13223 => x"2e",
         13224 => x"87",
         13225 => x"5a",
         13226 => x"7d",
         13227 => x"80",
         13228 => x"70",
         13229 => x"f0",
         13230 => x"bb",
         13231 => x"84",
         13232 => x"80",
         13233 => x"74",
         13234 => x"bb",
         13235 => x"3d",
         13236 => x"b5",
         13237 => x"9e",
         13238 => x"bb",
         13239 => x"ff",
         13240 => x"74",
         13241 => x"86",
         13242 => x"bb",
         13243 => x"3d",
         13244 => x"e8",
         13245 => x"fe",
         13246 => x"52",
         13247 => x"f5",
         13248 => x"bb",
         13249 => x"84",
         13250 => x"80",
         13251 => x"80",
         13252 => x"38",
         13253 => x"59",
         13254 => x"70",
         13255 => x"33",
         13256 => x"05",
         13257 => x"15",
         13258 => x"38",
         13259 => x"0b",
         13260 => x"7d",
         13261 => x"a5",
         13262 => x"84",
         13263 => x"56",
         13264 => x"8a",
         13265 => x"8a",
         13266 => x"ff",
         13267 => x"bb",
         13268 => x"2e",
         13269 => x"fe",
         13270 => x"55",
         13271 => x"fe",
         13272 => x"08",
         13273 => x"52",
         13274 => x"ea",
         13275 => x"84",
         13276 => x"bb",
         13277 => x"2e",
         13278 => x"81",
         13279 => x"bb",
         13280 => x"19",
         13281 => x"16",
         13282 => x"59",
         13283 => x"77",
         13284 => x"83",
         13285 => x"74",
         13286 => x"81",
         13287 => x"38",
         13288 => x"53",
         13289 => x"81",
         13290 => x"fe",
         13291 => x"84",
         13292 => x"80",
         13293 => x"ff",
         13294 => x"76",
         13295 => x"78",
         13296 => x"38",
         13297 => x"08",
         13298 => x"5a",
         13299 => x"e5",
         13300 => x"38",
         13301 => x"80",
         13302 => x"56",
         13303 => x"2e",
         13304 => x"81",
         13305 => x"81",
         13306 => x"81",
         13307 => x"fe",
         13308 => x"84",
         13309 => x"57",
         13310 => x"08",
         13311 => x"86",
         13312 => x"76",
         13313 => x"bf",
         13314 => x"76",
         13315 => x"a0",
         13316 => x"80",
         13317 => x"05",
         13318 => x"15",
         13319 => x"38",
         13320 => x"0b",
         13321 => x"8b",
         13322 => x"57",
         13323 => x"81",
         13324 => x"76",
         13325 => x"58",
         13326 => x"55",
         13327 => x"fd",
         13328 => x"70",
         13329 => x"33",
         13330 => x"05",
         13331 => x"15",
         13332 => x"38",
         13333 => x"6b",
         13334 => x"34",
         13335 => x"0b",
         13336 => x"7d",
         13337 => x"f5",
         13338 => x"84",
         13339 => x"ce",
         13340 => x"fe",
         13341 => x"54",
         13342 => x"53",
         13343 => x"18",
         13344 => x"d5",
         13345 => x"bb",
         13346 => x"2e",
         13347 => x"80",
         13348 => x"bb",
         13349 => x"19",
         13350 => x"08",
         13351 => x"31",
         13352 => x"19",
         13353 => x"38",
         13354 => x"55",
         13355 => x"b1",
         13356 => x"84",
         13357 => x"e8",
         13358 => x"81",
         13359 => x"fe",
         13360 => x"84",
         13361 => x"57",
         13362 => x"08",
         13363 => x"b6",
         13364 => x"39",
         13365 => x"59",
         13366 => x"fd",
         13367 => x"a1",
         13368 => x"b4",
         13369 => x"19",
         13370 => x"7a",
         13371 => x"33",
         13372 => x"b6",
         13373 => x"39",
         13374 => x"60",
         13375 => x"05",
         13376 => x"33",
         13377 => x"89",
         13378 => x"2e",
         13379 => x"08",
         13380 => x"2e",
         13381 => x"33",
         13382 => x"2e",
         13383 => x"15",
         13384 => x"22",
         13385 => x"78",
         13386 => x"38",
         13387 => x"5f",
         13388 => x"38",
         13389 => x"56",
         13390 => x"38",
         13391 => x"81",
         13392 => x"17",
         13393 => x"38",
         13394 => x"70",
         13395 => x"06",
         13396 => x"80",
         13397 => x"38",
         13398 => x"22",
         13399 => x"70",
         13400 => x"57",
         13401 => x"86",
         13402 => x"15",
         13403 => x"30",
         13404 => x"9f",
         13405 => x"84",
         13406 => x"1c",
         13407 => x"53",
         13408 => x"81",
         13409 => x"38",
         13410 => x"78",
         13411 => x"82",
         13412 => x"56",
         13413 => x"74",
         13414 => x"fe",
         13415 => x"81",
         13416 => x"55",
         13417 => x"75",
         13418 => x"82",
         13419 => x"84",
         13420 => x"81",
         13421 => x"bb",
         13422 => x"2e",
         13423 => x"84",
         13424 => x"81",
         13425 => x"19",
         13426 => x"2e",
         13427 => x"78",
         13428 => x"06",
         13429 => x"56",
         13430 => x"84",
         13431 => x"90",
         13432 => x"87",
         13433 => x"84",
         13434 => x"0d",
         13435 => x"33",
         13436 => x"e5",
         13437 => x"84",
         13438 => x"54",
         13439 => x"38",
         13440 => x"55",
         13441 => x"39",
         13442 => x"81",
         13443 => x"7d",
         13444 => x"80",
         13445 => x"81",
         13446 => x"81",
         13447 => x"38",
         13448 => x"52",
         13449 => x"de",
         13450 => x"bb",
         13451 => x"84",
         13452 => x"ff",
         13453 => x"81",
         13454 => x"57",
         13455 => x"d7",
         13456 => x"90",
         13457 => x"7b",
         13458 => x"8c",
         13459 => x"18",
         13460 => x"18",
         13461 => x"33",
         13462 => x"5c",
         13463 => x"34",
         13464 => x"fe",
         13465 => x"08",
         13466 => x"7a",
         13467 => x"38",
         13468 => x"94",
         13469 => x"15",
         13470 => x"5d",
         13471 => x"34",
         13472 => x"d6",
         13473 => x"ff",
         13474 => x"5b",
         13475 => x"be",
         13476 => x"fe",
         13477 => x"54",
         13478 => x"ff",
         13479 => x"a1",
         13480 => x"90",
         13481 => x"0d",
         13482 => x"a5",
         13483 => x"88",
         13484 => x"05",
         13485 => x"5f",
         13486 => x"3d",
         13487 => x"5b",
         13488 => x"2e",
         13489 => x"79",
         13490 => x"5b",
         13491 => x"26",
         13492 => x"ba",
         13493 => x"38",
         13494 => x"75",
         13495 => x"92",
         13496 => x"e0",
         13497 => x"76",
         13498 => x"38",
         13499 => x"84",
         13500 => x"70",
         13501 => x"74",
         13502 => x"38",
         13503 => x"75",
         13504 => x"f8",
         13505 => x"ba",
         13506 => x"40",
         13507 => x"52",
         13508 => x"ce",
         13509 => x"bb",
         13510 => x"ff",
         13511 => x"06",
         13512 => x"57",
         13513 => x"38",
         13514 => x"81",
         13515 => x"57",
         13516 => x"38",
         13517 => x"05",
         13518 => x"79",
         13519 => x"e9",
         13520 => x"84",
         13521 => x"38",
         13522 => x"80",
         13523 => x"38",
         13524 => x"80",
         13525 => x"38",
         13526 => x"06",
         13527 => x"ff",
         13528 => x"2e",
         13529 => x"80",
         13530 => x"f8",
         13531 => x"80",
         13532 => x"f0",
         13533 => x"7f",
         13534 => x"83",
         13535 => x"89",
         13536 => x"08",
         13537 => x"89",
         13538 => x"4c",
         13539 => x"80",
         13540 => x"38",
         13541 => x"80",
         13542 => x"56",
         13543 => x"74",
         13544 => x"7d",
         13545 => x"df",
         13546 => x"74",
         13547 => x"79",
         13548 => x"f7",
         13549 => x"84",
         13550 => x"83",
         13551 => x"83",
         13552 => x"61",
         13553 => x"33",
         13554 => x"07",
         13555 => x"57",
         13556 => x"d5",
         13557 => x"06",
         13558 => x"7d",
         13559 => x"05",
         13560 => x"33",
         13561 => x"80",
         13562 => x"38",
         13563 => x"83",
         13564 => x"12",
         13565 => x"2b",
         13566 => x"07",
         13567 => x"70",
         13568 => x"2b",
         13569 => x"07",
         13570 => x"83",
         13571 => x"12",
         13572 => x"2b",
         13573 => x"07",
         13574 => x"70",
         13575 => x"2b",
         13576 => x"07",
         13577 => x"0c",
         13578 => x"0c",
         13579 => x"44",
         13580 => x"59",
         13581 => x"4b",
         13582 => x"57",
         13583 => x"27",
         13584 => x"93",
         13585 => x"80",
         13586 => x"38",
         13587 => x"70",
         13588 => x"49",
         13589 => x"83",
         13590 => x"87",
         13591 => x"82",
         13592 => x"61",
         13593 => x"66",
         13594 => x"83",
         13595 => x"4a",
         13596 => x"58",
         13597 => x"8a",
         13598 => x"ae",
         13599 => x"2a",
         13600 => x"83",
         13601 => x"56",
         13602 => x"2e",
         13603 => x"77",
         13604 => x"83",
         13605 => x"77",
         13606 => x"70",
         13607 => x"58",
         13608 => x"86",
         13609 => x"27",
         13610 => x"52",
         13611 => x"ff",
         13612 => x"bb",
         13613 => x"84",
         13614 => x"bb",
         13615 => x"f5",
         13616 => x"81",
         13617 => x"84",
         13618 => x"bb",
         13619 => x"71",
         13620 => x"83",
         13621 => x"43",
         13622 => x"89",
         13623 => x"5c",
         13624 => x"1f",
         13625 => x"05",
         13626 => x"05",
         13627 => x"72",
         13628 => x"57",
         13629 => x"2e",
         13630 => x"74",
         13631 => x"90",
         13632 => x"60",
         13633 => x"74",
         13634 => x"f2",
         13635 => x"31",
         13636 => x"53",
         13637 => x"52",
         13638 => x"89",
         13639 => x"84",
         13640 => x"83",
         13641 => x"38",
         13642 => x"09",
         13643 => x"dd",
         13644 => x"f5",
         13645 => x"84",
         13646 => x"ac",
         13647 => x"f9",
         13648 => x"55",
         13649 => x"26",
         13650 => x"74",
         13651 => x"39",
         13652 => x"84",
         13653 => x"9f",
         13654 => x"bb",
         13655 => x"81",
         13656 => x"39",
         13657 => x"bb",
         13658 => x"3d",
         13659 => x"90",
         13660 => x"33",
         13661 => x"81",
         13662 => x"57",
         13663 => x"26",
         13664 => x"1d",
         13665 => x"06",
         13666 => x"58",
         13667 => x"81",
         13668 => x"0b",
         13669 => x"5f",
         13670 => x"7d",
         13671 => x"70",
         13672 => x"33",
         13673 => x"05",
         13674 => x"9f",
         13675 => x"57",
         13676 => x"89",
         13677 => x"70",
         13678 => x"58",
         13679 => x"18",
         13680 => x"26",
         13681 => x"18",
         13682 => x"06",
         13683 => x"30",
         13684 => x"5a",
         13685 => x"2e",
         13686 => x"85",
         13687 => x"be",
         13688 => x"32",
         13689 => x"72",
         13690 => x"7b",
         13691 => x"4a",
         13692 => x"80",
         13693 => x"1c",
         13694 => x"5c",
         13695 => x"ff",
         13696 => x"56",
         13697 => x"9f",
         13698 => x"53",
         13699 => x"51",
         13700 => x"3f",
         13701 => x"bb",
         13702 => x"b6",
         13703 => x"2a",
         13704 => x"bb",
         13705 => x"56",
         13706 => x"bf",
         13707 => x"8e",
         13708 => x"26",
         13709 => x"74",
         13710 => x"fb",
         13711 => x"56",
         13712 => x"7b",
         13713 => x"ba",
         13714 => x"a3",
         13715 => x"f9",
         13716 => x"81",
         13717 => x"57",
         13718 => x"fd",
         13719 => x"6e",
         13720 => x"46",
         13721 => x"39",
         13722 => x"08",
         13723 => x"9d",
         13724 => x"38",
         13725 => x"81",
         13726 => x"fb",
         13727 => x"57",
         13728 => x"84",
         13729 => x"0d",
         13730 => x"0c",
         13731 => x"62",
         13732 => x"99",
         13733 => x"60",
         13734 => x"74",
         13735 => x"8e",
         13736 => x"ae",
         13737 => x"61",
         13738 => x"76",
         13739 => x"58",
         13740 => x"55",
         13741 => x"8b",
         13742 => x"c0",
         13743 => x"76",
         13744 => x"58",
         13745 => x"81",
         13746 => x"ff",
         13747 => x"ef",
         13748 => x"05",
         13749 => x"34",
         13750 => x"05",
         13751 => x"8d",
         13752 => x"83",
         13753 => x"4b",
         13754 => x"05",
         13755 => x"2a",
         13756 => x"8f",
         13757 => x"61",
         13758 => x"62",
         13759 => x"30",
         13760 => x"61",
         13761 => x"78",
         13762 => x"06",
         13763 => x"92",
         13764 => x"56",
         13765 => x"ff",
         13766 => x"38",
         13767 => x"ff",
         13768 => x"61",
         13769 => x"74",
         13770 => x"6b",
         13771 => x"34",
         13772 => x"05",
         13773 => x"98",
         13774 => x"61",
         13775 => x"ff",
         13776 => x"34",
         13777 => x"05",
         13778 => x"9c",
         13779 => x"88",
         13780 => x"61",
         13781 => x"7e",
         13782 => x"6b",
         13783 => x"34",
         13784 => x"84",
         13785 => x"84",
         13786 => x"61",
         13787 => x"62",
         13788 => x"f7",
         13789 => x"a7",
         13790 => x"61",
         13791 => x"a1",
         13792 => x"34",
         13793 => x"aa",
         13794 => x"83",
         13795 => x"55",
         13796 => x"05",
         13797 => x"2a",
         13798 => x"97",
         13799 => x"80",
         13800 => x"34",
         13801 => x"05",
         13802 => x"ab",
         13803 => x"cc",
         13804 => x"76",
         13805 => x"58",
         13806 => x"81",
         13807 => x"ff",
         13808 => x"ef",
         13809 => x"fe",
         13810 => x"d5",
         13811 => x"83",
         13812 => x"ff",
         13813 => x"81",
         13814 => x"60",
         13815 => x"fe",
         13816 => x"81",
         13817 => x"84",
         13818 => x"38",
         13819 => x"62",
         13820 => x"9c",
         13821 => x"57",
         13822 => x"70",
         13823 => x"34",
         13824 => x"74",
         13825 => x"75",
         13826 => x"83",
         13827 => x"38",
         13828 => x"f8",
         13829 => x"2e",
         13830 => x"57",
         13831 => x"76",
         13832 => x"45",
         13833 => x"70",
         13834 => x"34",
         13835 => x"59",
         13836 => x"81",
         13837 => x"76",
         13838 => x"75",
         13839 => x"57",
         13840 => x"66",
         13841 => x"76",
         13842 => x"7a",
         13843 => x"79",
         13844 => x"d6",
         13845 => x"84",
         13846 => x"38",
         13847 => x"57",
         13848 => x"70",
         13849 => x"34",
         13850 => x"74",
         13851 => x"1b",
         13852 => x"58",
         13853 => x"38",
         13854 => x"40",
         13855 => x"ff",
         13856 => x"56",
         13857 => x"83",
         13858 => x"65",
         13859 => x"26",
         13860 => x"55",
         13861 => x"53",
         13862 => x"51",
         13863 => x"3f",
         13864 => x"08",
         13865 => x"74",
         13866 => x"31",
         13867 => x"db",
         13868 => x"62",
         13869 => x"38",
         13870 => x"83",
         13871 => x"8a",
         13872 => x"62",
         13873 => x"38",
         13874 => x"84",
         13875 => x"83",
         13876 => x"5e",
         13877 => x"38",
         13878 => x"56",
         13879 => x"70",
         13880 => x"34",
         13881 => x"78",
         13882 => x"d5",
         13883 => x"aa",
         13884 => x"83",
         13885 => x"78",
         13886 => x"67",
         13887 => x"81",
         13888 => x"34",
         13889 => x"05",
         13890 => x"84",
         13891 => x"43",
         13892 => x"52",
         13893 => x"fc",
         13894 => x"fe",
         13895 => x"34",
         13896 => x"08",
         13897 => x"07",
         13898 => x"86",
         13899 => x"bb",
         13900 => x"87",
         13901 => x"61",
         13902 => x"34",
         13903 => x"c7",
         13904 => x"61",
         13905 => x"34",
         13906 => x"08",
         13907 => x"05",
         13908 => x"83",
         13909 => x"62",
         13910 => x"64",
         13911 => x"05",
         13912 => x"2a",
         13913 => x"83",
         13914 => x"62",
         13915 => x"7e",
         13916 => x"05",
         13917 => x"78",
         13918 => x"79",
         13919 => x"aa",
         13920 => x"84",
         13921 => x"f7",
         13922 => x"53",
         13923 => x"51",
         13924 => x"3f",
         13925 => x"bb",
         13926 => x"b6",
         13927 => x"84",
         13928 => x"84",
         13929 => x"0d",
         13930 => x"0c",
         13931 => x"f9",
         13932 => x"1c",
         13933 => x"5c",
         13934 => x"7a",
         13935 => x"91",
         13936 => x"0b",
         13937 => x"22",
         13938 => x"80",
         13939 => x"74",
         13940 => x"38",
         13941 => x"56",
         13942 => x"17",
         13943 => x"57",
         13944 => x"2e",
         13945 => x"75",
         13946 => x"77",
         13947 => x"fc",
         13948 => x"84",
         13949 => x"10",
         13950 => x"05",
         13951 => x"5e",
         13952 => x"80",
         13953 => x"84",
         13954 => x"8a",
         13955 => x"fd",
         13956 => x"77",
         13957 => x"38",
         13958 => x"e4",
         13959 => x"84",
         13960 => x"f5",
         13961 => x"38",
         13962 => x"38",
         13963 => x"5b",
         13964 => x"38",
         13965 => x"c8",
         13966 => x"06",
         13967 => x"2e",
         13968 => x"83",
         13969 => x"39",
         13970 => x"05",
         13971 => x"2a",
         13972 => x"a1",
         13973 => x"90",
         13974 => x"61",
         13975 => x"75",
         13976 => x"76",
         13977 => x"34",
         13978 => x"80",
         13979 => x"05",
         13980 => x"80",
         13981 => x"a1",
         13982 => x"05",
         13983 => x"61",
         13984 => x"34",
         13985 => x"05",
         13986 => x"2a",
         13987 => x"a5",
         13988 => x"90",
         13989 => x"61",
         13990 => x"7c",
         13991 => x"75",
         13992 => x"34",
         13993 => x"05",
         13994 => x"ad",
         13995 => x"61",
         13996 => x"80",
         13997 => x"34",
         13998 => x"05",
         13999 => x"b1",
         14000 => x"61",
         14001 => x"80",
         14002 => x"34",
         14003 => x"80",
         14004 => x"a9",
         14005 => x"05",
         14006 => x"80",
         14007 => x"e6",
         14008 => x"55",
         14009 => x"05",
         14010 => x"70",
         14011 => x"34",
         14012 => x"74",
         14013 => x"cd",
         14014 => x"81",
         14015 => x"76",
         14016 => x"58",
         14017 => x"55",
         14018 => x"f9",
         14019 => x"54",
         14020 => x"52",
         14021 => x"bf",
         14022 => x"57",
         14023 => x"08",
         14024 => x"7d",
         14025 => x"05",
         14026 => x"83",
         14027 => x"76",
         14028 => x"84",
         14029 => x"52",
         14030 => x"bf",
         14031 => x"c3",
         14032 => x"84",
         14033 => x"9f",
         14034 => x"bb",
         14035 => x"f8",
         14036 => x"4a",
         14037 => x"81",
         14038 => x"ff",
         14039 => x"05",
         14040 => x"6a",
         14041 => x"84",
         14042 => x"61",
         14043 => x"ff",
         14044 => x"34",
         14045 => x"05",
         14046 => x"88",
         14047 => x"61",
         14048 => x"ff",
         14049 => x"34",
         14050 => x"7c",
         14051 => x"39",
         14052 => x"1f",
         14053 => x"79",
         14054 => x"8e",
         14055 => x"61",
         14056 => x"75",
         14057 => x"57",
         14058 => x"57",
         14059 => x"60",
         14060 => x"7c",
         14061 => x"5e",
         14062 => x"80",
         14063 => x"81",
         14064 => x"80",
         14065 => x"81",
         14066 => x"80",
         14067 => x"80",
         14068 => x"e4",
         14069 => x"f2",
         14070 => x"05",
         14071 => x"61",
         14072 => x"34",
         14073 => x"83",
         14074 => x"7f",
         14075 => x"7a",
         14076 => x"05",
         14077 => x"2a",
         14078 => x"83",
         14079 => x"7a",
         14080 => x"75",
         14081 => x"05",
         14082 => x"2a",
         14083 => x"83",
         14084 => x"82",
         14085 => x"05",
         14086 => x"83",
         14087 => x"76",
         14088 => x"05",
         14089 => x"83",
         14090 => x"80",
         14091 => x"ff",
         14092 => x"81",
         14093 => x"53",
         14094 => x"51",
         14095 => x"3f",
         14096 => x"1f",
         14097 => x"79",
         14098 => x"de",
         14099 => x"57",
         14100 => x"39",
         14101 => x"7e",
         14102 => x"80",
         14103 => x"05",
         14104 => x"76",
         14105 => x"38",
         14106 => x"8e",
         14107 => x"54",
         14108 => x"52",
         14109 => x"9b",
         14110 => x"81",
         14111 => x"06",
         14112 => x"3d",
         14113 => x"8d",
         14114 => x"74",
         14115 => x"05",
         14116 => x"17",
         14117 => x"2e",
         14118 => x"77",
         14119 => x"80",
         14120 => x"55",
         14121 => x"76",
         14122 => x"bb",
         14123 => x"3d",
         14124 => x"3d",
         14125 => x"84",
         14126 => x"33",
         14127 => x"8a",
         14128 => x"38",
         14129 => x"56",
         14130 => x"9e",
         14131 => x"08",
         14132 => x"05",
         14133 => x"75",
         14134 => x"55",
         14135 => x"8e",
         14136 => x"18",
         14137 => x"88",
         14138 => x"3d",
         14139 => x"3d",
         14140 => x"74",
         14141 => x"52",
         14142 => x"ff",
         14143 => x"74",
         14144 => x"30",
         14145 => x"9f",
         14146 => x"84",
         14147 => x"1c",
         14148 => x"5a",
         14149 => x"39",
         14150 => x"51",
         14151 => x"ff",
         14152 => x"3d",
         14153 => x"ff",
         14154 => x"3d",
         14155 => x"cc",
         14156 => x"80",
         14157 => x"05",
         14158 => x"15",
         14159 => x"38",
         14160 => x"77",
         14161 => x"2e",
         14162 => x"7c",
         14163 => x"24",
         14164 => x"7d",
         14165 => x"05",
         14166 => x"75",
         14167 => x"55",
         14168 => x"b8",
         14169 => x"18",
         14170 => x"88",
         14171 => x"55",
         14172 => x"9e",
         14173 => x"ff",
         14174 => x"75",
         14175 => x"52",
         14176 => x"ff",
         14177 => x"84",
         14178 => x"86",
         14179 => x"2e",
         14180 => x"0b",
         14181 => x"0c",
         14182 => x"04",
         14183 => x"b0",
         14184 => x"54",
         14185 => x"76",
         14186 => x"9d",
         14187 => x"7b",
         14188 => x"70",
         14189 => x"2a",
         14190 => x"5a",
         14191 => x"a5",
         14192 => x"76",
         14193 => x"3f",
         14194 => x"7d",
         14195 => x"0c",
         14196 => x"04",
         14197 => x"75",
         14198 => x"9a",
         14199 => x"53",
         14200 => x"80",
         14201 => x"38",
         14202 => x"ff",
         14203 => x"84",
         14204 => x"85",
         14205 => x"83",
         14206 => x"27",
         14207 => x"b5",
         14208 => x"06",
         14209 => x"80",
         14210 => x"83",
         14211 => x"51",
         14212 => x"9c",
         14213 => x"70",
         14214 => x"06",
         14215 => x"80",
         14216 => x"38",
         14217 => x"e8",
         14218 => x"22",
         14219 => x"39",
         14220 => x"70",
         14221 => x"84",
         14222 => x"53",
         14223 => x"04",
         14224 => x"02",
         14225 => x"02",
         14226 => x"05",
         14227 => x"80",
         14228 => x"ff",
         14229 => x"70",
         14230 => x"bb",
         14231 => x"3d",
         14232 => x"83",
         14233 => x"81",
         14234 => x"70",
         14235 => x"e9",
         14236 => x"83",
         14237 => x"70",
         14238 => x"84",
         14239 => x"3d",
         14240 => x"3d",
         14241 => x"70",
         14242 => x"26",
         14243 => x"70",
         14244 => x"06",
         14245 => x"56",
         14246 => x"ff",
         14247 => x"38",
         14248 => x"05",
         14249 => x"71",
         14250 => x"25",
         14251 => x"07",
         14252 => x"53",
         14253 => x"71",
         14254 => x"53",
         14255 => x"88",
         14256 => x"81",
         14257 => x"14",
         14258 => x"76",
         14259 => x"71",
         14260 => x"10",
         14261 => x"82",
         14262 => x"54",
         14263 => x"80",
         14264 => x"26",
         14265 => x"52",
         14266 => x"cb",
         14267 => x"70",
         14268 => x"0c",
         14269 => x"04",
         14270 => x"55",
         14271 => x"71",
         14272 => x"38",
         14273 => x"83",
         14274 => x"54",
         14275 => x"c7",
         14276 => x"83",
         14277 => x"57",
         14278 => x"d3",
         14279 => x"16",
         14280 => x"ff",
         14281 => x"f1",
         14282 => x"70",
         14283 => x"06",
         14284 => x"39",
         14285 => x"83",
         14286 => x"57",
         14287 => x"d0",
         14288 => x"ff",
         14289 => x"51",
         14290 => x"16",
         14291 => x"ff",
         14292 => x"c5",
         14293 => x"70",
         14294 => x"06",
         14295 => x"b9",
         14296 => x"31",
         14297 => x"71",
         14298 => x"ff",
         14299 => x"52",
         14300 => x"39",
         14301 => x"10",
         14302 => x"22",
         14303 => x"ef",
         14304 => x"00",
         14305 => x"ff",
         14306 => x"ff",
         14307 => x"ff",
         14308 => x"00",
         14309 => x"8b",
         14310 => x"80",
         14311 => x"75",
         14312 => x"6a",
         14313 => x"5f",
         14314 => x"54",
         14315 => x"49",
         14316 => x"3e",
         14317 => x"33",
         14318 => x"28",
         14319 => x"1d",
         14320 => x"12",
         14321 => x"07",
         14322 => x"fc",
         14323 => x"f1",
         14324 => x"e6",
         14325 => x"db",
         14326 => x"d0",
         14327 => x"c5",
         14328 => x"ba",
         14329 => x"ca",
         14330 => x"64",
         14331 => x"64",
         14332 => x"64",
         14333 => x"64",
         14334 => x"64",
         14335 => x"64",
         14336 => x"64",
         14337 => x"64",
         14338 => x"64",
         14339 => x"64",
         14340 => x"64",
         14341 => x"64",
         14342 => x"64",
         14343 => x"64",
         14344 => x"64",
         14345 => x"64",
         14346 => x"64",
         14347 => x"64",
         14348 => x"64",
         14349 => x"64",
         14350 => x"64",
         14351 => x"64",
         14352 => x"64",
         14353 => x"64",
         14354 => x"64",
         14355 => x"64",
         14356 => x"64",
         14357 => x"64",
         14358 => x"64",
         14359 => x"64",
         14360 => x"64",
         14361 => x"64",
         14362 => x"64",
         14363 => x"64",
         14364 => x"64",
         14365 => x"64",
         14366 => x"64",
         14367 => x"64",
         14368 => x"64",
         14369 => x"64",
         14370 => x"64",
         14371 => x"64",
         14372 => x"81",
         14373 => x"64",
         14374 => x"64",
         14375 => x"64",
         14376 => x"64",
         14377 => x"64",
         14378 => x"64",
         14379 => x"64",
         14380 => x"64",
         14381 => x"64",
         14382 => x"64",
         14383 => x"64",
         14384 => x"64",
         14385 => x"64",
         14386 => x"64",
         14387 => x"64",
         14388 => x"64",
         14389 => x"17",
         14390 => x"16",
         14391 => x"64",
         14392 => x"9a",
         14393 => x"b8",
         14394 => x"77",
         14395 => x"3c",
         14396 => x"de",
         14397 => x"64",
         14398 => x"64",
         14399 => x"64",
         14400 => x"64",
         14401 => x"64",
         14402 => x"64",
         14403 => x"64",
         14404 => x"64",
         14405 => x"64",
         14406 => x"64",
         14407 => x"64",
         14408 => x"64",
         14409 => x"64",
         14410 => x"64",
         14411 => x"64",
         14412 => x"64",
         14413 => x"64",
         14414 => x"64",
         14415 => x"64",
         14416 => x"64",
         14417 => x"64",
         14418 => x"64",
         14419 => x"64",
         14420 => x"64",
         14421 => x"64",
         14422 => x"64",
         14423 => x"64",
         14424 => x"64",
         14425 => x"64",
         14426 => x"64",
         14427 => x"64",
         14428 => x"64",
         14429 => x"64",
         14430 => x"64",
         14431 => x"64",
         14432 => x"64",
         14433 => x"64",
         14434 => x"64",
         14435 => x"64",
         14436 => x"64",
         14437 => x"64",
         14438 => x"64",
         14439 => x"64",
         14440 => x"64",
         14441 => x"64",
         14442 => x"64",
         14443 => x"64",
         14444 => x"64",
         14445 => x"64",
         14446 => x"64",
         14447 => x"64",
         14448 => x"64",
         14449 => x"bb",
         14450 => x"80",
         14451 => x"64",
         14452 => x"64",
         14453 => x"64",
         14454 => x"64",
         14455 => x"64",
         14456 => x"64",
         14457 => x"64",
         14458 => x"64",
         14459 => x"73",
         14460 => x"68",
         14461 => x"64",
         14462 => x"50",
         14463 => x"64",
         14464 => x"61",
         14465 => x"56",
         14466 => x"49",
         14467 => x"33",
         14468 => x"4b",
         14469 => x"57",
         14470 => x"63",
         14471 => x"6f",
         14472 => x"3f",
         14473 => x"10",
         14474 => x"9a",
         14475 => x"62",
         14476 => x"90",
         14477 => x"ac",
         14478 => x"fd",
         14479 => x"fc",
         14480 => x"b5",
         14481 => x"44",
         14482 => x"e4",
         14483 => x"59",
         14484 => x"8b",
         14485 => x"fd",
         14486 => x"62",
         14487 => x"6c",
         14488 => x"fc",
         14489 => x"fd",
         14490 => x"fd",
         14491 => x"59",
         14492 => x"e4",
         14493 => x"b5",
         14494 => x"90",
         14495 => x"44",
         14496 => x"5d",
         14497 => x"82",
         14498 => x"a3",
         14499 => x"04",
         14500 => x"c8",
         14501 => x"1d",
         14502 => x"6d",
         14503 => x"2a",
         14504 => x"2a",
         14505 => x"2a",
         14506 => x"2a",
         14507 => x"2a",
         14508 => x"2a",
         14509 => x"03",
         14510 => x"2a",
         14511 => x"2a",
         14512 => x"2a",
         14513 => x"2a",
         14514 => x"2a",
         14515 => x"2a",
         14516 => x"2a",
         14517 => x"2a",
         14518 => x"2a",
         14519 => x"2a",
         14520 => x"2a",
         14521 => x"2a",
         14522 => x"2a",
         14523 => x"2a",
         14524 => x"2a",
         14525 => x"2a",
         14526 => x"2a",
         14527 => x"2a",
         14528 => x"2a",
         14529 => x"2a",
         14530 => x"2a",
         14531 => x"2a",
         14532 => x"42",
         14533 => x"30",
         14534 => x"1d",
         14535 => x"0a",
         14536 => x"34",
         14537 => x"f8",
         14538 => x"e5",
         14539 => x"4d",
         14540 => x"2a",
         14541 => x"4d",
         14542 => x"d5",
         14543 => x"52",
         14544 => x"7e",
         14545 => x"5c",
         14546 => x"c3",
         14547 => x"b1",
         14548 => x"9f",
         14549 => x"90",
         14550 => x"2a",
         14551 => x"34",
         14552 => x"d0",
         14553 => x"3f",
         14554 => x"11",
         14555 => x"68",
         14556 => x"45",
         14557 => x"24",
         14558 => x"fa",
         14559 => x"ca",
         14560 => x"51",
         14561 => x"a4",
         14562 => x"93",
         14563 => x"51",
         14564 => x"51",
         14565 => x"51",
         14566 => x"51",
         14567 => x"51",
         14568 => x"51",
         14569 => x"6d",
         14570 => x"7b",
         14571 => x"32",
         14572 => x"51",
         14573 => x"51",
         14574 => x"51",
         14575 => x"51",
         14576 => x"51",
         14577 => x"51",
         14578 => x"51",
         14579 => x"51",
         14580 => x"51",
         14581 => x"51",
         14582 => x"51",
         14583 => x"51",
         14584 => x"51",
         14585 => x"51",
         14586 => x"51",
         14587 => x"51",
         14588 => x"51",
         14589 => x"51",
         14590 => x"51",
         14591 => x"ef",
         14592 => x"51",
         14593 => x"51",
         14594 => x"51",
         14595 => x"92",
         14596 => x"a1",
         14597 => x"43",
         14598 => x"51",
         14599 => x"51",
         14600 => x"51",
         14601 => x"51",
         14602 => x"28",
         14603 => x"51",
         14604 => x"0b",
         14605 => x"74",
         14606 => x"e9",
         14607 => x"e9",
         14608 => x"e9",
         14609 => x"e9",
         14610 => x"e9",
         14611 => x"e9",
         14612 => x"c4",
         14613 => x"e9",
         14614 => x"e9",
         14615 => x"e9",
         14616 => x"e9",
         14617 => x"e9",
         14618 => x"e9",
         14619 => x"e9",
         14620 => x"e9",
         14621 => x"e9",
         14622 => x"e9",
         14623 => x"e9",
         14624 => x"e9",
         14625 => x"e9",
         14626 => x"e9",
         14627 => x"e9",
         14628 => x"e9",
         14629 => x"e9",
         14630 => x"e9",
         14631 => x"e9",
         14632 => x"e9",
         14633 => x"e9",
         14634 => x"e9",
         14635 => x"86",
         14636 => x"ce",
         14637 => x"bb",
         14638 => x"a8",
         14639 => x"96",
         14640 => x"59",
         14641 => x"46",
         14642 => x"36",
         14643 => x"e9",
         14644 => x"26",
         14645 => x"16",
         14646 => x"04",
         14647 => x"f2",
         14648 => x"e0",
         14649 => x"51",
         14650 => x"40",
         14651 => x"2f",
         14652 => x"18",
         14653 => x"e9",
         14654 => x"62",
         14655 => x"43",
         14656 => x"9f",
         14657 => x"9f",
         14658 => x"9f",
         14659 => x"9f",
         14660 => x"9f",
         14661 => x"9f",
         14662 => x"9f",
         14663 => x"9f",
         14664 => x"9f",
         14665 => x"9f",
         14666 => x"9f",
         14667 => x"9f",
         14668 => x"9f",
         14669 => x"c1",
         14670 => x"9f",
         14671 => x"9f",
         14672 => x"9f",
         14673 => x"9f",
         14674 => x"9f",
         14675 => x"9f",
         14676 => x"8d",
         14677 => x"9f",
         14678 => x"9f",
         14679 => x"18",
         14680 => x"9f",
         14681 => x"2f",
         14682 => x"a0",
         14683 => x"01",
         14684 => x"74",
         14685 => x"61",
         14686 => x"55",
         14687 => x"4a",
         14688 => x"3f",
         14689 => x"34",
         14690 => x"29",
         14691 => x"1d",
         14692 => x"0f",
         14693 => x"01",
         14694 => x"fd",
         14695 => x"fd",
         14696 => x"49",
         14697 => x"fd",
         14698 => x"fd",
         14699 => x"fd",
         14700 => x"fd",
         14701 => x"fd",
         14702 => x"fd",
         14703 => x"fd",
         14704 => x"fd",
         14705 => x"fd",
         14706 => x"7f",
         14707 => x"0d",
         14708 => x"fd",
         14709 => x"fd",
         14710 => x"fd",
         14711 => x"fd",
         14712 => x"fd",
         14713 => x"fd",
         14714 => x"fd",
         14715 => x"fd",
         14716 => x"fd",
         14717 => x"fd",
         14718 => x"fd",
         14719 => x"fd",
         14720 => x"fd",
         14721 => x"fd",
         14722 => x"fd",
         14723 => x"fd",
         14724 => x"fd",
         14725 => x"fd",
         14726 => x"fd",
         14727 => x"fd",
         14728 => x"fd",
         14729 => x"fd",
         14730 => x"fd",
         14731 => x"fd",
         14732 => x"fd",
         14733 => x"fd",
         14734 => x"fd",
         14735 => x"fd",
         14736 => x"fd",
         14737 => x"fd",
         14738 => x"fd",
         14739 => x"fd",
         14740 => x"fd",
         14741 => x"fd",
         14742 => x"fd",
         14743 => x"fd",
         14744 => x"1d",
         14745 => x"fd",
         14746 => x"fd",
         14747 => x"fd",
         14748 => x"fd",
         14749 => x"17",
         14750 => x"fd",
         14751 => x"fd",
         14752 => x"fd",
         14753 => x"fd",
         14754 => x"fd",
         14755 => x"fd",
         14756 => x"fd",
         14757 => x"fd",
         14758 => x"fd",
         14759 => x"fd",
         14760 => x"2b",
         14761 => x"e1",
         14762 => x"b8",
         14763 => x"b8",
         14764 => x"b8",
         14765 => x"fd",
         14766 => x"e1",
         14767 => x"fd",
         14768 => x"fd",
         14769 => x"ff",
         14770 => x"fd",
         14771 => x"fd",
         14772 => x"16",
         14773 => x"0f",
         14774 => x"fd",
         14775 => x"fd",
         14776 => x"58",
         14777 => x"fd",
         14778 => x"18",
         14779 => x"fd",
         14780 => x"fd",
         14781 => x"17",
         14782 => x"69",
         14783 => x"00",
         14784 => x"63",
         14785 => x"00",
         14786 => x"69",
         14787 => x"00",
         14788 => x"61",
         14789 => x"00",
         14790 => x"65",
         14791 => x"00",
         14792 => x"65",
         14793 => x"00",
         14794 => x"70",
         14795 => x"00",
         14796 => x"66",
         14797 => x"00",
         14798 => x"6d",
         14799 => x"00",
         14800 => x"00",
         14801 => x"00",
         14802 => x"00",
         14803 => x"00",
         14804 => x"00",
         14805 => x"00",
         14806 => x"00",
         14807 => x"6c",
         14808 => x"00",
         14809 => x"00",
         14810 => x"74",
         14811 => x"00",
         14812 => x"65",
         14813 => x"00",
         14814 => x"6f",
         14815 => x"00",
         14816 => x"74",
         14817 => x"00",
         14818 => x"00",
         14819 => x"00",
         14820 => x"73",
         14821 => x"00",
         14822 => x"73",
         14823 => x"00",
         14824 => x"6f",
         14825 => x"00",
         14826 => x"00",
         14827 => x"6e",
         14828 => x"20",
         14829 => x"6f",
         14830 => x"00",
         14831 => x"61",
         14832 => x"65",
         14833 => x"69",
         14834 => x"72",
         14835 => x"74",
         14836 => x"00",
         14837 => x"20",
         14838 => x"79",
         14839 => x"65",
         14840 => x"69",
         14841 => x"2e",
         14842 => x"00",
         14843 => x"75",
         14844 => x"63",
         14845 => x"74",
         14846 => x"6d",
         14847 => x"2e",
         14848 => x"00",
         14849 => x"65",
         14850 => x"20",
         14851 => x"6b",
         14852 => x"00",
         14853 => x"65",
         14854 => x"2c",
         14855 => x"65",
         14856 => x"69",
         14857 => x"63",
         14858 => x"65",
         14859 => x"64",
         14860 => x"00",
         14861 => x"6d",
         14862 => x"61",
         14863 => x"74",
         14864 => x"00",
         14865 => x"63",
         14866 => x"61",
         14867 => x"6c",
         14868 => x"69",
         14869 => x"79",
         14870 => x"6d",
         14871 => x"75",
         14872 => x"6f",
         14873 => x"69",
         14874 => x"00",
         14875 => x"6b",
         14876 => x"74",
         14877 => x"61",
         14878 => x"64",
         14879 => x"00",
         14880 => x"76",
         14881 => x"75",
         14882 => x"72",
         14883 => x"20",
         14884 => x"61",
         14885 => x"2e",
         14886 => x"00",
         14887 => x"69",
         14888 => x"72",
         14889 => x"20",
         14890 => x"74",
         14891 => x"65",
         14892 => x"00",
         14893 => x"65",
         14894 => x"6e",
         14895 => x"20",
         14896 => x"61",
         14897 => x"2e",
         14898 => x"00",
         14899 => x"65",
         14900 => x"72",
         14901 => x"79",
         14902 => x"69",
         14903 => x"2e",
         14904 => x"00",
         14905 => x"65",
         14906 => x"64",
         14907 => x"65",
         14908 => x"00",
         14909 => x"61",
         14910 => x"20",
         14911 => x"65",
         14912 => x"65",
         14913 => x"00",
         14914 => x"70",
         14915 => x"20",
         14916 => x"6e",
         14917 => x"00",
         14918 => x"66",
         14919 => x"20",
         14920 => x"6e",
         14921 => x"00",
         14922 => x"6b",
         14923 => x"74",
         14924 => x"61",
         14925 => x"00",
         14926 => x"65",
         14927 => x"6c",
         14928 => x"72",
         14929 => x"00",
         14930 => x"6b",
         14931 => x"72",
         14932 => x"00",
         14933 => x"63",
         14934 => x"2e",
         14935 => x"00",
         14936 => x"75",
         14937 => x"74",
         14938 => x"25",
         14939 => x"74",
         14940 => x"75",
         14941 => x"74",
         14942 => x"73",
         14943 => x"0a",
         14944 => x"00",
         14945 => x"64",
         14946 => x"00",
         14947 => x"6c",
         14948 => x"00",
         14949 => x"00",
         14950 => x"58",
         14951 => x"00",
         14952 => x"00",
         14953 => x"00",
         14954 => x"00",
         14955 => x"58",
         14956 => x"00",
         14957 => x"20",
         14958 => x"20",
         14959 => x"00",
         14960 => x"00",
         14961 => x"25",
         14962 => x"00",
         14963 => x"30",
         14964 => x"30",
         14965 => x"00",
         14966 => x"33",
         14967 => x"00",
         14968 => x"55",
         14969 => x"65",
         14970 => x"30",
         14971 => x"20",
         14972 => x"25",
         14973 => x"2a",
         14974 => x"00",
         14975 => x"00",
         14976 => x"20",
         14977 => x"65",
         14978 => x"64",
         14979 => x"73",
         14980 => x"20",
         14981 => x"20",
         14982 => x"20",
         14983 => x"25",
         14984 => x"78",
         14985 => x"00",
         14986 => x"20",
         14987 => x"20",
         14988 => x"72",
         14989 => x"20",
         14990 => x"20",
         14991 => x"20",
         14992 => x"20",
         14993 => x"25",
         14994 => x"78",
         14995 => x"00",
         14996 => x"20",
         14997 => x"65",
         14998 => x"70",
         14999 => x"61",
         15000 => x"65",
         15001 => x"00",
         15002 => x"54",
         15003 => x"58",
         15004 => x"74",
         15005 => x"75",
         15006 => x"00",
         15007 => x"54",
         15008 => x"58",
         15009 => x"74",
         15010 => x"75",
         15011 => x"00",
         15012 => x"54",
         15013 => x"58",
         15014 => x"74",
         15015 => x"75",
         15016 => x"00",
         15017 => x"54",
         15018 => x"58",
         15019 => x"74",
         15020 => x"75",
         15021 => x"00",
         15022 => x"54",
         15023 => x"52",
         15024 => x"74",
         15025 => x"75",
         15026 => x"00",
         15027 => x"54",
         15028 => x"44",
         15029 => x"74",
         15030 => x"75",
         15031 => x"00",
         15032 => x"20",
         15033 => x"65",
         15034 => x"70",
         15035 => x"00",
         15036 => x"65",
         15037 => x"6e",
         15038 => x"72",
         15039 => x"00",
         15040 => x"74",
         15041 => x"20",
         15042 => x"74",
         15043 => x"72",
         15044 => x"00",
         15045 => x"62",
         15046 => x"67",
         15047 => x"6d",
         15048 => x"2e",
         15049 => x"00",
         15050 => x"6f",
         15051 => x"63",
         15052 => x"74",
         15053 => x"00",
         15054 => x"5f",
         15055 => x"2e",
         15056 => x"00",
         15057 => x"6c",
         15058 => x"74",
         15059 => x"6e",
         15060 => x"61",
         15061 => x"65",
         15062 => x"20",
         15063 => x"64",
         15064 => x"20",
         15065 => x"61",
         15066 => x"69",
         15067 => x"20",
         15068 => x"75",
         15069 => x"79",
         15070 => x"00",
         15071 => x"00",
         15072 => x"5c",
         15073 => x"00",
         15074 => x"00",
         15075 => x"20",
         15076 => x"6d",
         15077 => x"2e",
         15078 => x"00",
         15079 => x"00",
         15080 => x"00",
         15081 => x"5c",
         15082 => x"25",
         15083 => x"73",
         15084 => x"00",
         15085 => x"64",
         15086 => x"62",
         15087 => x"69",
         15088 => x"2e",
         15089 => x"00",
         15090 => x"74",
         15091 => x"69",
         15092 => x"61",
         15093 => x"69",
         15094 => x"69",
         15095 => x"2e",
         15096 => x"00",
         15097 => x"6c",
         15098 => x"20",
         15099 => x"65",
         15100 => x"25",
         15101 => x"78",
         15102 => x"2e",
         15103 => x"00",
         15104 => x"6c",
         15105 => x"74",
         15106 => x"65",
         15107 => x"6f",
         15108 => x"28",
         15109 => x"2e",
         15110 => x"00",
         15111 => x"63",
         15112 => x"6e",
         15113 => x"6f",
         15114 => x"40",
         15115 => x"38",
         15116 => x"2e",
         15117 => x"00",
         15118 => x"6c",
         15119 => x"30",
         15120 => x"2d",
         15121 => x"00",
         15122 => x"6c",
         15123 => x"30",
         15124 => x"00",
         15125 => x"70",
         15126 => x"6e",
         15127 => x"2e",
         15128 => x"00",
         15129 => x"6c",
         15130 => x"30",
         15131 => x"2d",
         15132 => x"38",
         15133 => x"25",
         15134 => x"29",
         15135 => x"00",
         15136 => x"79",
         15137 => x"2e",
         15138 => x"00",
         15139 => x"6c",
         15140 => x"30",
         15141 => x"00",
         15142 => x"61",
         15143 => x"67",
         15144 => x"2e",
         15145 => x"00",
         15146 => x"70",
         15147 => x"6d",
         15148 => x"00",
         15149 => x"6d",
         15150 => x"74",
         15151 => x"00",
         15152 => x"5c",
         15153 => x"25",
         15154 => x"00",
         15155 => x"6f",
         15156 => x"65",
         15157 => x"75",
         15158 => x"64",
         15159 => x"61",
         15160 => x"74",
         15161 => x"6f",
         15162 => x"73",
         15163 => x"6d",
         15164 => x"64",
         15165 => x"00",
         15166 => x"00",
         15167 => x"25",
         15168 => x"64",
         15169 => x"3a",
         15170 => x"25",
         15171 => x"64",
         15172 => x"00",
         15173 => x"20",
         15174 => x"66",
         15175 => x"72",
         15176 => x"6f",
         15177 => x"00",
         15178 => x"65",
         15179 => x"65",
         15180 => x"6d",
         15181 => x"6d",
         15182 => x"65",
         15183 => x"00",
         15184 => x"72",
         15185 => x"65",
         15186 => x"00",
         15187 => x"20",
         15188 => x"20",
         15189 => x"65",
         15190 => x"65",
         15191 => x"72",
         15192 => x"64",
         15193 => x"73",
         15194 => x"25",
         15195 => x"0a",
         15196 => x"00",
         15197 => x"20",
         15198 => x"20",
         15199 => x"6f",
         15200 => x"53",
         15201 => x"74",
         15202 => x"64",
         15203 => x"73",
         15204 => x"25",
         15205 => x"0a",
         15206 => x"00",
         15207 => x"20",
         15208 => x"63",
         15209 => x"74",
         15210 => x"20",
         15211 => x"72",
         15212 => x"20",
         15213 => x"20",
         15214 => x"25",
         15215 => x"0a",
         15216 => x"00",
         15217 => x"63",
         15218 => x"00",
         15219 => x"20",
         15220 => x"20",
         15221 => x"20",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"20",
         15226 => x"25",
         15227 => x"0a",
         15228 => x"00",
         15229 => x"20",
         15230 => x"74",
         15231 => x"43",
         15232 => x"6b",
         15233 => x"65",
         15234 => x"20",
         15235 => x"20",
         15236 => x"25",
         15237 => x"30",
         15238 => x"48",
         15239 => x"00",
         15240 => x"20",
         15241 => x"68",
         15242 => x"65",
         15243 => x"52",
         15244 => x"43",
         15245 => x"6b",
         15246 => x"65",
         15247 => x"25",
         15248 => x"30",
         15249 => x"48",
         15250 => x"00",
         15251 => x"20",
         15252 => x"41",
         15253 => x"6c",
         15254 => x"20",
         15255 => x"71",
         15256 => x"20",
         15257 => x"20",
         15258 => x"25",
         15259 => x"30",
         15260 => x"48",
         15261 => x"00",
         15262 => x"20",
         15263 => x"00",
         15264 => x"20",
         15265 => x"00",
         15266 => x"20",
         15267 => x"54",
         15268 => x"00",
         15269 => x"20",
         15270 => x"49",
         15271 => x"00",
         15272 => x"20",
         15273 => x"48",
         15274 => x"45",
         15275 => x"53",
         15276 => x"00",
         15277 => x"20",
         15278 => x"52",
         15279 => x"52",
         15280 => x"43",
         15281 => x"6e",
         15282 => x"3d",
         15283 => x"64",
         15284 => x"00",
         15285 => x"20",
         15286 => x"45",
         15287 => x"20",
         15288 => x"54",
         15289 => x"72",
         15290 => x"3d",
         15291 => x"64",
         15292 => x"00",
         15293 => x"20",
         15294 => x"43",
         15295 => x"20",
         15296 => x"44",
         15297 => x"63",
         15298 => x"3d",
         15299 => x"64",
         15300 => x"00",
         15301 => x"20",
         15302 => x"20",
         15303 => x"20",
         15304 => x"25",
         15305 => x"3a",
         15306 => x"58",
         15307 => x"00",
         15308 => x"20",
         15309 => x"4d",
         15310 => x"20",
         15311 => x"25",
         15312 => x"3a",
         15313 => x"58",
         15314 => x"00",
         15315 => x"20",
         15316 => x"4e",
         15317 => x"41",
         15318 => x"25",
         15319 => x"3a",
         15320 => x"58",
         15321 => x"00",
         15322 => x"20",
         15323 => x"41",
         15324 => x"20",
         15325 => x"25",
         15326 => x"3a",
         15327 => x"58",
         15328 => x"00",
         15329 => x"20",
         15330 => x"53",
         15331 => x"4d",
         15332 => x"25",
         15333 => x"3a",
         15334 => x"58",
         15335 => x"00",
         15336 => x"72",
         15337 => x"53",
         15338 => x"63",
         15339 => x"69",
         15340 => x"00",
         15341 => x"6e",
         15342 => x"00",
         15343 => x"6d",
         15344 => x"00",
         15345 => x"6c",
         15346 => x"00",
         15347 => x"69",
         15348 => x"00",
         15349 => x"78",
         15350 => x"00",
         15351 => x"00",
         15352 => x"3c",
         15353 => x"00",
         15354 => x"02",
         15355 => x"38",
         15356 => x"00",
         15357 => x"03",
         15358 => x"34",
         15359 => x"00",
         15360 => x"04",
         15361 => x"30",
         15362 => x"00",
         15363 => x"05",
         15364 => x"2c",
         15365 => x"00",
         15366 => x"06",
         15367 => x"28",
         15368 => x"00",
         15369 => x"07",
         15370 => x"24",
         15371 => x"00",
         15372 => x"01",
         15373 => x"20",
         15374 => x"00",
         15375 => x"08",
         15376 => x"1c",
         15377 => x"00",
         15378 => x"0b",
         15379 => x"18",
         15380 => x"00",
         15381 => x"09",
         15382 => x"14",
         15383 => x"00",
         15384 => x"0a",
         15385 => x"10",
         15386 => x"00",
         15387 => x"0d",
         15388 => x"0c",
         15389 => x"00",
         15390 => x"0c",
         15391 => x"08",
         15392 => x"00",
         15393 => x"0e",
         15394 => x"04",
         15395 => x"00",
         15396 => x"0f",
         15397 => x"00",
         15398 => x"00",
         15399 => x"0f",
         15400 => x"fc",
         15401 => x"00",
         15402 => x"10",
         15403 => x"f8",
         15404 => x"00",
         15405 => x"11",
         15406 => x"f4",
         15407 => x"00",
         15408 => x"12",
         15409 => x"f0",
         15410 => x"00",
         15411 => x"13",
         15412 => x"ec",
         15413 => x"00",
         15414 => x"14",
         15415 => x"e8",
         15416 => x"00",
         15417 => x"15",
         15418 => x"00",
         15419 => x"00",
         15420 => x"00",
         15421 => x"00",
         15422 => x"7e",
         15423 => x"7e",
         15424 => x"7e",
         15425 => x"00",
         15426 => x"7e",
         15427 => x"7e",
         15428 => x"7e",
         15429 => x"00",
         15430 => x"00",
         15431 => x"00",
         15432 => x"00",
         15433 => x"00",
         15434 => x"00",
         15435 => x"00",
         15436 => x"00",
         15437 => x"00",
         15438 => x"00",
         15439 => x"00",
         15440 => x"74",
         15441 => x"20",
         15442 => x"70",
         15443 => x"38",
         15444 => x"00",
         15445 => x"6e",
         15446 => x"6f",
         15447 => x"2f",
         15448 => x"61",
         15449 => x"68",
         15450 => x"6f",
         15451 => x"66",
         15452 => x"2c",
         15453 => x"73",
         15454 => x"69",
         15455 => x"00",
         15456 => x"74",
         15457 => x"00",
         15458 => x"74",
         15459 => x"00",
         15460 => x"00",
         15461 => x"74",
         15462 => x"20",
         15463 => x"66",
         15464 => x"25",
         15465 => x"78",
         15466 => x"00",
         15467 => x"6c",
         15468 => x"25",
         15469 => x"00",
         15470 => x"6c",
         15471 => x"74",
         15472 => x"65",
         15473 => x"20",
         15474 => x"20",
         15475 => x"74",
         15476 => x"20",
         15477 => x"65",
         15478 => x"20",
         15479 => x"2e",
         15480 => x"00",
         15481 => x"0a",
         15482 => x"00",
         15483 => x"7e",
         15484 => x"00",
         15485 => x"00",
         15486 => x"00",
         15487 => x"00",
         15488 => x"00",
         15489 => x"30",
         15490 => x"00",
         15491 => x"31",
         15492 => x"00",
         15493 => x"32",
         15494 => x"00",
         15495 => x"33",
         15496 => x"00",
         15497 => x"34",
         15498 => x"00",
         15499 => x"35",
         15500 => x"00",
         15501 => x"37",
         15502 => x"00",
         15503 => x"38",
         15504 => x"00",
         15505 => x"39",
         15506 => x"00",
         15507 => x"30",
         15508 => x"00",
         15509 => x"7e",
         15510 => x"00",
         15511 => x"7e",
         15512 => x"00",
         15513 => x"00",
         15514 => x"7e",
         15515 => x"00",
         15516 => x"7e",
         15517 => x"00",
         15518 => x"64",
         15519 => x"2c",
         15520 => x"25",
         15521 => x"64",
         15522 => x"3a",
         15523 => x"78",
         15524 => x"00",
         15525 => x"64",
         15526 => x"2d",
         15527 => x"25",
         15528 => x"64",
         15529 => x"2c",
         15530 => x"00",
         15531 => x"00",
         15532 => x"64",
         15533 => x"00",
         15534 => x"78",
         15535 => x"00",
         15536 => x"25",
         15537 => x"64",
         15538 => x"00",
         15539 => x"6f",
         15540 => x"43",
         15541 => x"6f",
         15542 => x"00",
         15543 => x"25",
         15544 => x"20",
         15545 => x"78",
         15546 => x"00",
         15547 => x"25",
         15548 => x"20",
         15549 => x"78",
         15550 => x"00",
         15551 => x"25",
         15552 => x"20",
         15553 => x"00",
         15554 => x"74",
         15555 => x"20",
         15556 => x"69",
         15557 => x"2e",
         15558 => x"00",
         15559 => x"00",
         15560 => x"3c",
         15561 => x"7f",
         15562 => x"00",
         15563 => x"3d",
         15564 => x"00",
         15565 => x"00",
         15566 => x"33",
         15567 => x"00",
         15568 => x"4d",
         15569 => x"53",
         15570 => x"00",
         15571 => x"4e",
         15572 => x"20",
         15573 => x"46",
         15574 => x"20",
         15575 => x"00",
         15576 => x"4e",
         15577 => x"20",
         15578 => x"46",
         15579 => x"32",
         15580 => x"00",
         15581 => x"1c",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"07",
         15586 => x"12",
         15587 => x"1c",
         15588 => x"00",
         15589 => x"41",
         15590 => x"80",
         15591 => x"49",
         15592 => x"8f",
         15593 => x"4f",
         15594 => x"55",
         15595 => x"9b",
         15596 => x"9f",
         15597 => x"55",
         15598 => x"a7",
         15599 => x"ab",
         15600 => x"af",
         15601 => x"b3",
         15602 => x"b7",
         15603 => x"bb",
         15604 => x"bf",
         15605 => x"c3",
         15606 => x"c7",
         15607 => x"cb",
         15608 => x"cf",
         15609 => x"d3",
         15610 => x"d7",
         15611 => x"db",
         15612 => x"df",
         15613 => x"e3",
         15614 => x"e7",
         15615 => x"eb",
         15616 => x"ef",
         15617 => x"f3",
         15618 => x"f7",
         15619 => x"fb",
         15620 => x"ff",
         15621 => x"3b",
         15622 => x"2f",
         15623 => x"3a",
         15624 => x"7c",
         15625 => x"00",
         15626 => x"04",
         15627 => x"40",
         15628 => x"00",
         15629 => x"00",
         15630 => x"02",
         15631 => x"08",
         15632 => x"20",
         15633 => x"00",
         15634 => x"fc",
         15635 => x"e2",
         15636 => x"e0",
         15637 => x"e7",
         15638 => x"eb",
         15639 => x"ef",
         15640 => x"ec",
         15641 => x"c5",
         15642 => x"e6",
         15643 => x"f4",
         15644 => x"f2",
         15645 => x"f9",
         15646 => x"d6",
         15647 => x"a2",
         15648 => x"a5",
         15649 => x"92",
         15650 => x"ed",
         15651 => x"fa",
         15652 => x"d1",
         15653 => x"ba",
         15654 => x"10",
         15655 => x"bd",
         15656 => x"a1",
         15657 => x"bb",
         15658 => x"92",
         15659 => x"02",
         15660 => x"61",
         15661 => x"56",
         15662 => x"63",
         15663 => x"57",
         15664 => x"5c",
         15665 => x"10",
         15666 => x"34",
         15667 => x"1c",
         15668 => x"3c",
         15669 => x"5f",
         15670 => x"54",
         15671 => x"66",
         15672 => x"50",
         15673 => x"67",
         15674 => x"64",
         15675 => x"59",
         15676 => x"52",
         15677 => x"6b",
         15678 => x"18",
         15679 => x"88",
         15680 => x"8c",
         15681 => x"80",
         15682 => x"df",
         15683 => x"c0",
         15684 => x"c3",
         15685 => x"c4",
         15686 => x"98",
         15687 => x"b4",
         15688 => x"c6",
         15689 => x"29",
         15690 => x"b1",
         15691 => x"64",
         15692 => x"21",
         15693 => x"48",
         15694 => x"19",
         15695 => x"1a",
         15696 => x"b2",
         15697 => x"a0",
         15698 => x"1a",
         15699 => x"17",
         15700 => x"07",
         15701 => x"01",
         15702 => x"00",
         15703 => x"32",
         15704 => x"39",
         15705 => x"4a",
         15706 => x"79",
         15707 => x"80",
         15708 => x"43",
         15709 => x"82",
         15710 => x"84",
         15711 => x"86",
         15712 => x"87",
         15713 => x"8a",
         15714 => x"8b",
         15715 => x"8e",
         15716 => x"90",
         15717 => x"91",
         15718 => x"94",
         15719 => x"96",
         15720 => x"98",
         15721 => x"3d",
         15722 => x"9c",
         15723 => x"20",
         15724 => x"a0",
         15725 => x"a2",
         15726 => x"a4",
         15727 => x"a6",
         15728 => x"a7",
         15729 => x"aa",
         15730 => x"ac",
         15731 => x"ae",
         15732 => x"af",
         15733 => x"b2",
         15734 => x"b3",
         15735 => x"b5",
         15736 => x"b8",
         15737 => x"ba",
         15738 => x"bc",
         15739 => x"be",
         15740 => x"c0",
         15741 => x"c2",
         15742 => x"c4",
         15743 => x"c4",
         15744 => x"c8",
         15745 => x"ca",
         15746 => x"ca",
         15747 => x"10",
         15748 => x"01",
         15749 => x"de",
         15750 => x"f3",
         15751 => x"f1",
         15752 => x"f4",
         15753 => x"28",
         15754 => x"12",
         15755 => x"09",
         15756 => x"3b",
         15757 => x"3d",
         15758 => x"3f",
         15759 => x"41",
         15760 => x"46",
         15761 => x"53",
         15762 => x"81",
         15763 => x"55",
         15764 => x"8a",
         15765 => x"8f",
         15766 => x"90",
         15767 => x"5d",
         15768 => x"5f",
         15769 => x"61",
         15770 => x"94",
         15771 => x"65",
         15772 => x"67",
         15773 => x"96",
         15774 => x"62",
         15775 => x"6d",
         15776 => x"9c",
         15777 => x"71",
         15778 => x"73",
         15779 => x"9f",
         15780 => x"77",
         15781 => x"79",
         15782 => x"7b",
         15783 => x"64",
         15784 => x"7f",
         15785 => x"81",
         15786 => x"a9",
         15787 => x"85",
         15788 => x"87",
         15789 => x"44",
         15790 => x"b2",
         15791 => x"8d",
         15792 => x"8f",
         15793 => x"91",
         15794 => x"7b",
         15795 => x"fd",
         15796 => x"ff",
         15797 => x"04",
         15798 => x"88",
         15799 => x"8a",
         15800 => x"11",
         15801 => x"02",
         15802 => x"a3",
         15803 => x"08",
         15804 => x"03",
         15805 => x"8e",
         15806 => x"d8",
         15807 => x"f2",
         15808 => x"f9",
         15809 => x"f4",
         15810 => x"f6",
         15811 => x"f7",
         15812 => x"fa",
         15813 => x"30",
         15814 => x"50",
         15815 => x"60",
         15816 => x"8a",
         15817 => x"c1",
         15818 => x"cf",
         15819 => x"c0",
         15820 => x"44",
         15821 => x"26",
         15822 => x"00",
         15823 => x"01",
         15824 => x"00",
         15825 => x"a0",
         15826 => x"00",
         15827 => x"10",
         15828 => x"20",
         15829 => x"30",
         15830 => x"40",
         15831 => x"51",
         15832 => x"59",
         15833 => x"5b",
         15834 => x"5d",
         15835 => x"5f",
         15836 => x"08",
         15837 => x"0e",
         15838 => x"bb",
         15839 => x"c9",
         15840 => x"cb",
         15841 => x"db",
         15842 => x"f9",
         15843 => x"eb",
         15844 => x"fb",
         15845 => x"08",
         15846 => x"08",
         15847 => x"08",
         15848 => x"04",
         15849 => x"b9",
         15850 => x"bc",
         15851 => x"01",
         15852 => x"d0",
         15853 => x"e0",
         15854 => x"e5",
         15855 => x"ec",
         15856 => x"01",
         15857 => x"4e",
         15858 => x"32",
         15859 => x"10",
         15860 => x"01",
         15861 => x"d0",
         15862 => x"30",
         15863 => x"60",
         15864 => x"67",
         15865 => x"75",
         15866 => x"80",
         15867 => x"00",
         15868 => x"41",
         15869 => x"00",
         15870 => x"00",
         15871 => x"f8",
         15872 => x"00",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"00",
         15877 => x"00",
         15878 => x"00",
         15879 => x"08",
         15880 => x"00",
         15881 => x"00",
         15882 => x"00",
         15883 => x"10",
         15884 => x"00",
         15885 => x"00",
         15886 => x"00",
         15887 => x"18",
         15888 => x"00",
         15889 => x"00",
         15890 => x"00",
         15891 => x"20",
         15892 => x"00",
         15893 => x"00",
         15894 => x"00",
         15895 => x"28",
         15896 => x"00",
         15897 => x"00",
         15898 => x"00",
         15899 => x"30",
         15900 => x"00",
         15901 => x"00",
         15902 => x"00",
         15903 => x"38",
         15904 => x"00",
         15905 => x"00",
         15906 => x"00",
         15907 => x"40",
         15908 => x"00",
         15909 => x"00",
         15910 => x"00",
         15911 => x"44",
         15912 => x"00",
         15913 => x"00",
         15914 => x"00",
         15915 => x"48",
         15916 => x"00",
         15917 => x"00",
         15918 => x"00",
         15919 => x"4c",
         15920 => x"00",
         15921 => x"00",
         15922 => x"00",
         15923 => x"50",
         15924 => x"00",
         15925 => x"00",
         15926 => x"00",
         15927 => x"54",
         15928 => x"00",
         15929 => x"00",
         15930 => x"00",
         15931 => x"58",
         15932 => x"00",
         15933 => x"00",
         15934 => x"00",
         15935 => x"5c",
         15936 => x"00",
         15937 => x"00",
         15938 => x"00",
         15939 => x"64",
         15940 => x"00",
         15941 => x"00",
         15942 => x"00",
         15943 => x"68",
         15944 => x"00",
         15945 => x"00",
         15946 => x"00",
         15947 => x"70",
         15948 => x"00",
         15949 => x"00",
         15950 => x"00",
         15951 => x"78",
         15952 => x"00",
         15953 => x"00",
         15954 => x"00",
         15955 => x"80",
         15956 => x"00",
         15957 => x"00",
         15958 => x"00",
         15959 => x"88",
         15960 => x"00",
         15961 => x"00",
         15962 => x"00",
         15963 => x"8c",
         15964 => x"00",
         15965 => x"00",
         15966 => x"00",
         15967 => x"90",
         15968 => x"00",
         15969 => x"00",
         15970 => x"00",
         15971 => x"98",
         15972 => x"00",
         15973 => x"00",
         15974 => x"00",
         15975 => x"a0",
         15976 => x"00",
         15977 => x"00",
         15978 => x"00",
         15979 => x"a8",
         15980 => x"00",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"ff",
         15986 => x"00",
         15987 => x"ff",
         15988 => x"00",
         15989 => x"ff",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"ff",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"00",
         15999 => x"00",
         16000 => x"00",
         16001 => x"00",
         16002 => x"01",
         16003 => x"01",
         16004 => x"01",
         16005 => x"00",
         16006 => x"00",
         16007 => x"00",
         16008 => x"00",
         16009 => x"00",
         16010 => x"00",
         16011 => x"00",
         16012 => x"00",
         16013 => x"00",
         16014 => x"00",
         16015 => x"00",
         16016 => x"00",
         16017 => x"00",
         16018 => x"00",
         16019 => x"00",
         16020 => x"00",
         16021 => x"00",
         16022 => x"00",
         16023 => x"00",
         16024 => x"00",
         16025 => x"00",
         16026 => x"00",
         16027 => x"00",
         16028 => x"00",
         16029 => x"00",
         16030 => x"80",
         16031 => x"00",
         16032 => x"88",
         16033 => x"00",
         16034 => x"90",
         16035 => x"00",
         16036 => x"80",
         16037 => x"fd",
         16038 => x"0d",
         16039 => x"5b",
         16040 => x"f0",
         16041 => x"74",
         16042 => x"78",
         16043 => x"6c",
         16044 => x"70",
         16045 => x"64",
         16046 => x"68",
         16047 => x"34",
         16048 => x"38",
         16049 => x"20",
         16050 => x"2e",
         16051 => x"f4",
         16052 => x"2f",
         16053 => x"f0",
         16054 => x"f0",
         16055 => x"83",
         16056 => x"f0",
         16057 => x"fd",
         16058 => x"0d",
         16059 => x"5b",
         16060 => x"f0",
         16061 => x"54",
         16062 => x"58",
         16063 => x"4c",
         16064 => x"50",
         16065 => x"44",
         16066 => x"48",
         16067 => x"34",
         16068 => x"38",
         16069 => x"20",
         16070 => x"2e",
         16071 => x"f4",
         16072 => x"2f",
         16073 => x"f0",
         16074 => x"f0",
         16075 => x"83",
         16076 => x"f0",
         16077 => x"fd",
         16078 => x"0d",
         16079 => x"7b",
         16080 => x"f0",
         16081 => x"54",
         16082 => x"58",
         16083 => x"4c",
         16084 => x"50",
         16085 => x"44",
         16086 => x"48",
         16087 => x"24",
         16088 => x"28",
         16089 => x"20",
         16090 => x"3e",
         16091 => x"e1",
         16092 => x"2f",
         16093 => x"f0",
         16094 => x"f0",
         16095 => x"88",
         16096 => x"f0",
         16097 => x"fa",
         16098 => x"f0",
         16099 => x"1b",
         16100 => x"f0",
         16101 => x"14",
         16102 => x"18",
         16103 => x"0c",
         16104 => x"10",
         16105 => x"04",
         16106 => x"08",
         16107 => x"f0",
         16108 => x"f0",
         16109 => x"f0",
         16110 => x"f0",
         16111 => x"f0",
         16112 => x"1c",
         16113 => x"f0",
         16114 => x"f0",
         16115 => x"83",
         16116 => x"f0",
         16117 => x"c9",
         16118 => x"cd",
         16119 => x"b3",
         16120 => x"f0",
         16121 => x"31",
         16122 => x"dd",
         16123 => x"56",
         16124 => x"b1",
         16125 => x"48",
         16126 => x"73",
         16127 => x"3b",
         16128 => x"a2",
         16129 => x"00",
         16130 => x"b9",
         16131 => x"c1",
         16132 => x"be",
         16133 => x"f0",
         16134 => x"f0",
         16135 => x"83",
         16136 => x"f0",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"ec",
         16166 => x"00",
         16167 => x"f4",
         16168 => x"00",
         16169 => x"f8",
         16170 => x"00",
         16171 => x"fc",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"04",
         16176 => x"00",
         16177 => x"0c",
         16178 => x"00",
         16179 => x"14",
         16180 => x"00",
         16181 => x"1c",
         16182 => x"00",
         16183 => x"24",
         16184 => x"00",
         16185 => x"2c",
         16186 => x"00",
         16187 => x"34",
         16188 => x"00",
         16189 => x"3c",
         16190 => x"00",
         16191 => x"44",
         16192 => x"00",
         16193 => x"4c",
         16194 => x"00",
         16195 => x"54",
         16196 => x"00",
         16197 => x"5c",
         16198 => x"00",
         16199 => x"64",
         16200 => x"00",
         16201 => x"68",
         16202 => x"00",
         16203 => x"70",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"19",
         18206 => x"00",
         18207 => x"00",
         18208 => x"f3",
         18209 => x"f7",
         18210 => x"fb",
         18211 => x"ff",
         18212 => x"c3",
         18213 => x"e2",
         18214 => x"e6",
         18215 => x"f4",
         18216 => x"63",
         18217 => x"67",
         18218 => x"6a",
         18219 => x"2d",
         18220 => x"23",
         18221 => x"27",
         18222 => x"2c",
         18223 => x"49",
         18224 => x"03",
         18225 => x"07",
         18226 => x"0b",
         18227 => x"0f",
         18228 => x"13",
         18229 => x"17",
         18230 => x"52",
         18231 => x"3c",
         18232 => x"83",
         18233 => x"87",
         18234 => x"8b",
         18235 => x"8f",
         18236 => x"93",
         18237 => x"97",
         18238 => x"bc",
         18239 => x"c0",
         18240 => x"00",
         18241 => x"00",
         18242 => x"00",
         18243 => x"00",
         18244 => x"00",
         18245 => x"00",
         18246 => x"00",
         18247 => x"00",
         18248 => x"00",
         18249 => x"00",
         18250 => x"00",
         18251 => x"00",
         18252 => x"00",
         18253 => x"00",
         18254 => x"00",
         18255 => x"00",
         18256 => x"00",
         18257 => x"00",
         18258 => x"00",
         18259 => x"00",
         18260 => x"00",
         18261 => x"00",
         18262 => x"00",
         18263 => x"00",
         18264 => x"00",
         18265 => x"00",
         18266 => x"00",
         18267 => x"00",
         18268 => x"00",
         18269 => x"00",
         18270 => x"03",
         18271 => x"01",
         18272 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"e9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"83",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a6",
           270 => x"0b",
           271 => x"0b",
           272 => x"c6",
           273 => x"0b",
           274 => x"0b",
           275 => x"e6",
           276 => x"0b",
           277 => x"0b",
           278 => x"86",
           279 => x"0b",
           280 => x"0b",
           281 => x"a6",
           282 => x"0b",
           283 => x"0b",
           284 => x"c6",
           285 => x"0b",
           286 => x"0b",
           287 => x"e8",
           288 => x"0b",
           289 => x"0b",
           290 => x"8a",
           291 => x"0b",
           292 => x"0b",
           293 => x"ac",
           294 => x"0b",
           295 => x"0b",
           296 => x"ce",
           297 => x"0b",
           298 => x"0b",
           299 => x"f0",
           300 => x"0b",
           301 => x"0b",
           302 => x"92",
           303 => x"0b",
           304 => x"0b",
           305 => x"b4",
           306 => x"0b",
           307 => x"0b",
           308 => x"d6",
           309 => x"0b",
           310 => x"0b",
           311 => x"f8",
           312 => x"0b",
           313 => x"0b",
           314 => x"9a",
           315 => x"0b",
           316 => x"0b",
           317 => x"bc",
           318 => x"0b",
           319 => x"0b",
           320 => x"de",
           321 => x"0b",
           322 => x"0b",
           323 => x"80",
           324 => x"0b",
           325 => x"0b",
           326 => x"a2",
           327 => x"0b",
           328 => x"0b",
           329 => x"c4",
           330 => x"0b",
           331 => x"0b",
           332 => x"e6",
           333 => x"0b",
           334 => x"0b",
           335 => x"88",
           336 => x"0b",
           337 => x"0b",
           338 => x"aa",
           339 => x"0b",
           340 => x"0b",
           341 => x"cb",
           342 => x"0b",
           343 => x"0b",
           344 => x"ed",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"bb",
           386 => x"d6",
           387 => x"bb",
           388 => x"c0",
           389 => x"84",
           390 => x"a2",
           391 => x"bb",
           392 => x"c0",
           393 => x"84",
           394 => x"a0",
           395 => x"bb",
           396 => x"c0",
           397 => x"84",
           398 => x"a0",
           399 => x"bb",
           400 => x"c0",
           401 => x"84",
           402 => x"94",
           403 => x"bb",
           404 => x"c0",
           405 => x"84",
           406 => x"a1",
           407 => x"bb",
           408 => x"c0",
           409 => x"84",
           410 => x"af",
           411 => x"bb",
           412 => x"c0",
           413 => x"84",
           414 => x"ad",
           415 => x"bb",
           416 => x"c0",
           417 => x"84",
           418 => x"94",
           419 => x"bb",
           420 => x"c0",
           421 => x"84",
           422 => x"95",
           423 => x"bb",
           424 => x"c0",
           425 => x"84",
           426 => x"95",
           427 => x"bb",
           428 => x"c0",
           429 => x"84",
           430 => x"b1",
           431 => x"bb",
           432 => x"c0",
           433 => x"84",
           434 => x"80",
           435 => x"84",
           436 => x"80",
           437 => x"04",
           438 => x"0c",
           439 => x"2d",
           440 => x"08",
           441 => x"90",
           442 => x"90",
           443 => x"b8",
           444 => x"90",
           445 => x"80",
           446 => x"bb",
           447 => x"d3",
           448 => x"bb",
           449 => x"c0",
           450 => x"84",
           451 => x"82",
           452 => x"84",
           453 => x"80",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"90",
           459 => x"90",
           460 => x"c5",
           461 => x"90",
           462 => x"80",
           463 => x"bb",
           464 => x"d9",
           465 => x"bb",
           466 => x"c0",
           467 => x"84",
           468 => x"82",
           469 => x"84",
           470 => x"80",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"90",
           476 => x"90",
           477 => x"b8",
           478 => x"90",
           479 => x"80",
           480 => x"bb",
           481 => x"f2",
           482 => x"bb",
           483 => x"c0",
           484 => x"84",
           485 => x"82",
           486 => x"84",
           487 => x"80",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"90",
           493 => x"90",
           494 => x"b1",
           495 => x"90",
           496 => x"80",
           497 => x"bb",
           498 => x"ff",
           499 => x"bb",
           500 => x"c0",
           501 => x"84",
           502 => x"83",
           503 => x"84",
           504 => x"80",
           505 => x"04",
           506 => x"0c",
           507 => x"2d",
           508 => x"08",
           509 => x"90",
           510 => x"90",
           511 => x"8c",
           512 => x"90",
           513 => x"80",
           514 => x"bb",
           515 => x"96",
           516 => x"bb",
           517 => x"c0",
           518 => x"84",
           519 => x"82",
           520 => x"84",
           521 => x"80",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"90",
           527 => x"90",
           528 => x"97",
           529 => x"90",
           530 => x"80",
           531 => x"bb",
           532 => x"f6",
           533 => x"bb",
           534 => x"c0",
           535 => x"84",
           536 => x"83",
           537 => x"84",
           538 => x"80",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"90",
           544 => x"90",
           545 => x"f8",
           546 => x"90",
           547 => x"80",
           548 => x"bb",
           549 => x"c8",
           550 => x"bb",
           551 => x"c0",
           552 => x"84",
           553 => x"83",
           554 => x"84",
           555 => x"80",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"90",
           561 => x"90",
           562 => x"d4",
           563 => x"90",
           564 => x"80",
           565 => x"bb",
           566 => x"f5",
           567 => x"bb",
           568 => x"c0",
           569 => x"84",
           570 => x"81",
           571 => x"84",
           572 => x"80",
           573 => x"04",
           574 => x"0c",
           575 => x"2d",
           576 => x"08",
           577 => x"90",
           578 => x"90",
           579 => x"ba",
           580 => x"90",
           581 => x"80",
           582 => x"bb",
           583 => x"d2",
           584 => x"bb",
           585 => x"c0",
           586 => x"84",
           587 => x"80",
           588 => x"84",
           589 => x"80",
           590 => x"04",
           591 => x"0c",
           592 => x"84",
           593 => x"80",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"90",
           599 => x"90",
           600 => x"84",
           601 => x"90",
           602 => x"80",
           603 => x"bb",
           604 => x"f3",
           605 => x"bb",
           606 => x"c0",
           607 => x"84",
           608 => x"81",
           609 => x"84",
           610 => x"80",
           611 => x"04",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"04",
           621 => x"81",
           622 => x"83",
           623 => x"05",
           624 => x"10",
           625 => x"72",
           626 => x"51",
           627 => x"72",
           628 => x"06",
           629 => x"72",
           630 => x"10",
           631 => x"10",
           632 => x"ed",
           633 => x"53",
           634 => x"bb",
           635 => x"e6",
           636 => x"38",
           637 => x"84",
           638 => x"0b",
           639 => x"ec",
           640 => x"51",
           641 => x"04",
           642 => x"0d",
           643 => x"70",
           644 => x"08",
           645 => x"52",
           646 => x"08",
           647 => x"3f",
           648 => x"04",
           649 => x"78",
           650 => x"11",
           651 => x"81",
           652 => x"25",
           653 => x"55",
           654 => x"72",
           655 => x"81",
           656 => x"38",
           657 => x"74",
           658 => x"30",
           659 => x"9f",
           660 => x"55",
           661 => x"74",
           662 => x"71",
           663 => x"38",
           664 => x"fa",
           665 => x"84",
           666 => x"bb",
           667 => x"2e",
           668 => x"bb",
           669 => x"70",
           670 => x"34",
           671 => x"8a",
           672 => x"70",
           673 => x"2a",
           674 => x"54",
           675 => x"cb",
           676 => x"34",
           677 => x"84",
           678 => x"88",
           679 => x"80",
           680 => x"84",
           681 => x"0d",
           682 => x"0d",
           683 => x"02",
           684 => x"05",
           685 => x"fe",
           686 => x"3d",
           687 => x"7e",
           688 => x"e4",
           689 => x"3f",
           690 => x"80",
           691 => x"3d",
           692 => x"3d",
           693 => x"88",
           694 => x"52",
           695 => x"3f",
           696 => x"04",
           697 => x"61",
           698 => x"5d",
           699 => x"8c",
           700 => x"1e",
           701 => x"2a",
           702 => x"06",
           703 => x"ff",
           704 => x"2e",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"81",
           709 => x"06",
           710 => x"80",
           711 => x"38",
           712 => x"7e",
           713 => x"a3",
           714 => x"32",
           715 => x"80",
           716 => x"55",
           717 => x"72",
           718 => x"38",
           719 => x"70",
           720 => x"06",
           721 => x"80",
           722 => x"7a",
           723 => x"5b",
           724 => x"76",
           725 => x"8c",
           726 => x"73",
           727 => x"0c",
           728 => x"04",
           729 => x"54",
           730 => x"10",
           731 => x"70",
           732 => x"98",
           733 => x"81",
           734 => x"8b",
           735 => x"98",
           736 => x"5b",
           737 => x"79",
           738 => x"38",
           739 => x"53",
           740 => x"38",
           741 => x"58",
           742 => x"f7",
           743 => x"39",
           744 => x"09",
           745 => x"38",
           746 => x"5a",
           747 => x"7c",
           748 => x"76",
           749 => x"ff",
           750 => x"52",
           751 => x"af",
           752 => x"57",
           753 => x"38",
           754 => x"7a",
           755 => x"81",
           756 => x"78",
           757 => x"70",
           758 => x"54",
           759 => x"e0",
           760 => x"80",
           761 => x"38",
           762 => x"83",
           763 => x"54",
           764 => x"73",
           765 => x"59",
           766 => x"27",
           767 => x"52",
           768 => x"eb",
           769 => x"33",
           770 => x"fe",
           771 => x"c7",
           772 => x"59",
           773 => x"88",
           774 => x"84",
           775 => x"7d",
           776 => x"06",
           777 => x"54",
           778 => x"5e",
           779 => x"51",
           780 => x"84",
           781 => x"81",
           782 => x"bb",
           783 => x"df",
           784 => x"72",
           785 => x"38",
           786 => x"08",
           787 => x"74",
           788 => x"05",
           789 => x"52",
           790 => x"ca",
           791 => x"84",
           792 => x"bb",
           793 => x"38",
           794 => x"94",
           795 => x"7b",
           796 => x"56",
           797 => x"8f",
           798 => x"80",
           799 => x"80",
           800 => x"90",
           801 => x"7a",
           802 => x"81",
           803 => x"73",
           804 => x"38",
           805 => x"80",
           806 => x"80",
           807 => x"90",
           808 => x"77",
           809 => x"29",
           810 => x"05",
           811 => x"2c",
           812 => x"2a",
           813 => x"54",
           814 => x"2e",
           815 => x"98",
           816 => x"ff",
           817 => x"78",
           818 => x"cc",
           819 => x"ff",
           820 => x"83",
           821 => x"2a",
           822 => x"74",
           823 => x"73",
           824 => x"f0",
           825 => x"31",
           826 => x"90",
           827 => x"80",
           828 => x"53",
           829 => x"85",
           830 => x"81",
           831 => x"54",
           832 => x"38",
           833 => x"81",
           834 => x"86",
           835 => x"85",
           836 => x"54",
           837 => x"38",
           838 => x"54",
           839 => x"38",
           840 => x"81",
           841 => x"80",
           842 => x"77",
           843 => x"80",
           844 => x"80",
           845 => x"2c",
           846 => x"80",
           847 => x"38",
           848 => x"51",
           849 => x"77",
           850 => x"80",
           851 => x"80",
           852 => x"2c",
           853 => x"73",
           854 => x"38",
           855 => x"53",
           856 => x"b2",
           857 => x"81",
           858 => x"81",
           859 => x"70",
           860 => x"55",
           861 => x"25",
           862 => x"52",
           863 => x"ef",
           864 => x"81",
           865 => x"81",
           866 => x"70",
           867 => x"55",
           868 => x"24",
           869 => x"87",
           870 => x"06",
           871 => x"80",
           872 => x"38",
           873 => x"2e",
           874 => x"76",
           875 => x"81",
           876 => x"80",
           877 => x"e2",
           878 => x"bb",
           879 => x"38",
           880 => x"1e",
           881 => x"5e",
           882 => x"7d",
           883 => x"2e",
           884 => x"ec",
           885 => x"06",
           886 => x"2e",
           887 => x"77",
           888 => x"80",
           889 => x"80",
           890 => x"2c",
           891 => x"80",
           892 => x"91",
           893 => x"a0",
           894 => x"3f",
           895 => x"90",
           896 => x"a0",
           897 => x"58",
           898 => x"87",
           899 => x"39",
           900 => x"07",
           901 => x"57",
           902 => x"84",
           903 => x"7e",
           904 => x"06",
           905 => x"55",
           906 => x"39",
           907 => x"05",
           908 => x"0a",
           909 => x"33",
           910 => x"72",
           911 => x"80",
           912 => x"80",
           913 => x"90",
           914 => x"5a",
           915 => x"5f",
           916 => x"70",
           917 => x"55",
           918 => x"38",
           919 => x"80",
           920 => x"80",
           921 => x"90",
           922 => x"5f",
           923 => x"fe",
           924 => x"52",
           925 => x"f7",
           926 => x"ff",
           927 => x"ff",
           928 => x"57",
           929 => x"ff",
           930 => x"38",
           931 => x"70",
           932 => x"33",
           933 => x"3f",
           934 => x"1a",
           935 => x"ff",
           936 => x"79",
           937 => x"2e",
           938 => x"7c",
           939 => x"81",
           940 => x"51",
           941 => x"e2",
           942 => x"0a",
           943 => x"0a",
           944 => x"80",
           945 => x"80",
           946 => x"90",
           947 => x"56",
           948 => x"87",
           949 => x"06",
           950 => x"7a",
           951 => x"fe",
           952 => x"60",
           953 => x"08",
           954 => x"41",
           955 => x"24",
           956 => x"7a",
           957 => x"06",
           958 => x"94",
           959 => x"39",
           960 => x"7c",
           961 => x"76",
           962 => x"f8",
           963 => x"88",
           964 => x"7c",
           965 => x"76",
           966 => x"f8",
           967 => x"60",
           968 => x"08",
           969 => x"56",
           970 => x"72",
           971 => x"75",
           972 => x"3f",
           973 => x"08",
           974 => x"06",
           975 => x"90",
           976 => x"72",
           977 => x"fe",
           978 => x"80",
           979 => x"33",
           980 => x"f7",
           981 => x"ff",
           982 => x"84",
           983 => x"77",
           984 => x"58",
           985 => x"81",
           986 => x"51",
           987 => x"84",
           988 => x"83",
           989 => x"78",
           990 => x"2b",
           991 => x"39",
           992 => x"07",
           993 => x"5b",
           994 => x"38",
           995 => x"77",
           996 => x"80",
           997 => x"80",
           998 => x"2c",
           999 => x"80",
          1000 => x"d6",
          1001 => x"a0",
          1002 => x"3f",
          1003 => x"52",
          1004 => x"bb",
          1005 => x"2e",
          1006 => x"fa",
          1007 => x"52",
          1008 => x"ab",
          1009 => x"2a",
          1010 => x"7e",
          1011 => x"8c",
          1012 => x"39",
          1013 => x"78",
          1014 => x"2b",
          1015 => x"7d",
          1016 => x"57",
          1017 => x"73",
          1018 => x"ff",
          1019 => x"52",
          1020 => x"fb",
          1021 => x"06",
          1022 => x"2e",
          1023 => x"ff",
          1024 => x"52",
          1025 => x"51",
          1026 => x"74",
          1027 => x"7a",
          1028 => x"f1",
          1029 => x"39",
          1030 => x"98",
          1031 => x"2c",
          1032 => x"b7",
          1033 => x"ab",
          1034 => x"3f",
          1035 => x"52",
          1036 => x"bb",
          1037 => x"39",
          1038 => x"51",
          1039 => x"84",
          1040 => x"83",
          1041 => x"78",
          1042 => x"2b",
          1043 => x"f3",
          1044 => x"07",
          1045 => x"83",
          1046 => x"52",
          1047 => x"99",
          1048 => x"0d",
          1049 => x"08",
          1050 => x"74",
          1051 => x"3f",
          1052 => x"04",
          1053 => x"78",
          1054 => x"84",
          1055 => x"85",
          1056 => x"81",
          1057 => x"70",
          1058 => x"56",
          1059 => x"ff",
          1060 => x"2e",
          1061 => x"80",
          1062 => x"70",
          1063 => x"33",
          1064 => x"2e",
          1065 => x"e6",
          1066 => x"72",
          1067 => x"08",
          1068 => x"84",
          1069 => x"80",
          1070 => x"ff",
          1071 => x"81",
          1072 => x"53",
          1073 => x"88",
          1074 => x"e8",
          1075 => x"39",
          1076 => x"08",
          1077 => x"e8",
          1078 => x"51",
          1079 => x"55",
          1080 => x"bb",
          1081 => x"2e",
          1082 => x"57",
          1083 => x"84",
          1084 => x"88",
          1085 => x"fa",
          1086 => x"7a",
          1087 => x"0b",
          1088 => x"70",
          1089 => x"32",
          1090 => x"51",
          1091 => x"ff",
          1092 => x"2e",
          1093 => x"92",
          1094 => x"81",
          1095 => x"53",
          1096 => x"09",
          1097 => x"38",
          1098 => x"84",
          1099 => x"88",
          1100 => x"73",
          1101 => x"55",
          1102 => x"80",
          1103 => x"74",
          1104 => x"90",
          1105 => x"72",
          1106 => x"84",
          1107 => x"e3",
          1108 => x"70",
          1109 => x"33",
          1110 => x"e3",
          1111 => x"ff",
          1112 => x"e6",
          1113 => x"73",
          1114 => x"83",
          1115 => x"fa",
          1116 => x"7a",
          1117 => x"70",
          1118 => x"32",
          1119 => x"56",
          1120 => x"56",
          1121 => x"73",
          1122 => x"06",
          1123 => x"2e",
          1124 => x"15",
          1125 => x"88",
          1126 => x"91",
          1127 => x"56",
          1128 => x"74",
          1129 => x"75",
          1130 => x"08",
          1131 => x"8c",
          1132 => x"56",
          1133 => x"84",
          1134 => x"0d",
          1135 => x"76",
          1136 => x"51",
          1137 => x"54",
          1138 => x"56",
          1139 => x"08",
          1140 => x"15",
          1141 => x"8c",
          1142 => x"56",
          1143 => x"3d",
          1144 => x"11",
          1145 => x"ff",
          1146 => x"32",
          1147 => x"55",
          1148 => x"54",
          1149 => x"72",
          1150 => x"06",
          1151 => x"38",
          1152 => x"81",
          1153 => x"80",
          1154 => x"38",
          1155 => x"33",
          1156 => x"80",
          1157 => x"38",
          1158 => x"0c",
          1159 => x"81",
          1160 => x"0c",
          1161 => x"06",
          1162 => x"bb",
          1163 => x"3d",
          1164 => x"ff",
          1165 => x"72",
          1166 => x"8c",
          1167 => x"05",
          1168 => x"84",
          1169 => x"bb",
          1170 => x"3d",
          1171 => x"51",
          1172 => x"55",
          1173 => x"bb",
          1174 => x"84",
          1175 => x"80",
          1176 => x"38",
          1177 => x"70",
          1178 => x"52",
          1179 => x"08",
          1180 => x"38",
          1181 => x"53",
          1182 => x"34",
          1183 => x"84",
          1184 => x"87",
          1185 => x"74",
          1186 => x"72",
          1187 => x"ff",
          1188 => x"fd",
          1189 => x"77",
          1190 => x"54",
          1191 => x"05",
          1192 => x"70",
          1193 => x"12",
          1194 => x"81",
          1195 => x"51",
          1196 => x"81",
          1197 => x"70",
          1198 => x"84",
          1199 => x"85",
          1200 => x"fc",
          1201 => x"79",
          1202 => x"55",
          1203 => x"80",
          1204 => x"73",
          1205 => x"38",
          1206 => x"93",
          1207 => x"81",
          1208 => x"73",
          1209 => x"55",
          1210 => x"51",
          1211 => x"73",
          1212 => x"0c",
          1213 => x"04",
          1214 => x"73",
          1215 => x"38",
          1216 => x"53",
          1217 => x"ff",
          1218 => x"71",
          1219 => x"ff",
          1220 => x"80",
          1221 => x"ff",
          1222 => x"53",
          1223 => x"73",
          1224 => x"51",
          1225 => x"c7",
          1226 => x"0d",
          1227 => x"53",
          1228 => x"05",
          1229 => x"70",
          1230 => x"12",
          1231 => x"84",
          1232 => x"51",
          1233 => x"04",
          1234 => x"75",
          1235 => x"54",
          1236 => x"81",
          1237 => x"51",
          1238 => x"81",
          1239 => x"70",
          1240 => x"84",
          1241 => x"85",
          1242 => x"fd",
          1243 => x"78",
          1244 => x"55",
          1245 => x"80",
          1246 => x"71",
          1247 => x"53",
          1248 => x"81",
          1249 => x"ff",
          1250 => x"ef",
          1251 => x"bb",
          1252 => x"3d",
          1253 => x"3d",
          1254 => x"7a",
          1255 => x"72",
          1256 => x"38",
          1257 => x"70",
          1258 => x"33",
          1259 => x"71",
          1260 => x"06",
          1261 => x"14",
          1262 => x"2e",
          1263 => x"13",
          1264 => x"38",
          1265 => x"84",
          1266 => x"86",
          1267 => x"72",
          1268 => x"38",
          1269 => x"ff",
          1270 => x"2e",
          1271 => x"15",
          1272 => x"51",
          1273 => x"de",
          1274 => x"31",
          1275 => x"0c",
          1276 => x"04",
          1277 => x"84",
          1278 => x"0d",
          1279 => x"0d",
          1280 => x"70",
          1281 => x"c1",
          1282 => x"84",
          1283 => x"84",
          1284 => x"52",
          1285 => x"b2",
          1286 => x"84",
          1287 => x"bb",
          1288 => x"2e",
          1289 => x"bb",
          1290 => x"54",
          1291 => x"74",
          1292 => x"84",
          1293 => x"51",
          1294 => x"84",
          1295 => x"54",
          1296 => x"84",
          1297 => x"0d",
          1298 => x"0d",
          1299 => x"71",
          1300 => x"54",
          1301 => x"9f",
          1302 => x"81",
          1303 => x"51",
          1304 => x"8c",
          1305 => x"52",
          1306 => x"09",
          1307 => x"38",
          1308 => x"75",
          1309 => x"70",
          1310 => x"0c",
          1311 => x"04",
          1312 => x"75",
          1313 => x"55",
          1314 => x"70",
          1315 => x"38",
          1316 => x"81",
          1317 => x"ff",
          1318 => x"f4",
          1319 => x"bb",
          1320 => x"3d",
          1321 => x"3d",
          1322 => x"58",
          1323 => x"76",
          1324 => x"38",
          1325 => x"f5",
          1326 => x"84",
          1327 => x"12",
          1328 => x"2e",
          1329 => x"51",
          1330 => x"71",
          1331 => x"08",
          1332 => x"52",
          1333 => x"80",
          1334 => x"52",
          1335 => x"80",
          1336 => x"13",
          1337 => x"a0",
          1338 => x"71",
          1339 => x"54",
          1340 => x"74",
          1341 => x"38",
          1342 => x"9f",
          1343 => x"10",
          1344 => x"72",
          1345 => x"9f",
          1346 => x"06",
          1347 => x"75",
          1348 => x"1c",
          1349 => x"52",
          1350 => x"53",
          1351 => x"73",
          1352 => x"52",
          1353 => x"84",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"80",
          1357 => x"30",
          1358 => x"80",
          1359 => x"2b",
          1360 => x"75",
          1361 => x"83",
          1362 => x"70",
          1363 => x"25",
          1364 => x"71",
          1365 => x"2a",
          1366 => x"06",
          1367 => x"80",
          1368 => x"84",
          1369 => x"71",
          1370 => x"75",
          1371 => x"8c",
          1372 => x"70",
          1373 => x"82",
          1374 => x"71",
          1375 => x"2a",
          1376 => x"81",
          1377 => x"82",
          1378 => x"75",
          1379 => x"bb",
          1380 => x"52",
          1381 => x"54",
          1382 => x"55",
          1383 => x"56",
          1384 => x"51",
          1385 => x"52",
          1386 => x"04",
          1387 => x"75",
          1388 => x"71",
          1389 => x"81",
          1390 => x"bb",
          1391 => x"29",
          1392 => x"84",
          1393 => x"53",
          1394 => x"04",
          1395 => x"78",
          1396 => x"a0",
          1397 => x"2e",
          1398 => x"51",
          1399 => x"84",
          1400 => x"53",
          1401 => x"73",
          1402 => x"38",
          1403 => x"bd",
          1404 => x"bb",
          1405 => x"52",
          1406 => x"9f",
          1407 => x"38",
          1408 => x"9f",
          1409 => x"81",
          1410 => x"2a",
          1411 => x"76",
          1412 => x"54",
          1413 => x"56",
          1414 => x"a8",
          1415 => x"74",
          1416 => x"74",
          1417 => x"78",
          1418 => x"11",
          1419 => x"81",
          1420 => x"06",
          1421 => x"ff",
          1422 => x"52",
          1423 => x"55",
          1424 => x"38",
          1425 => x"84",
          1426 => x"0d",
          1427 => x"0d",
          1428 => x"7a",
          1429 => x"9f",
          1430 => x"7c",
          1431 => x"32",
          1432 => x"71",
          1433 => x"72",
          1434 => x"59",
          1435 => x"56",
          1436 => x"84",
          1437 => x"75",
          1438 => x"84",
          1439 => x"88",
          1440 => x"f7",
          1441 => x"7d",
          1442 => x"70",
          1443 => x"08",
          1444 => x"56",
          1445 => x"2e",
          1446 => x"8f",
          1447 => x"70",
          1448 => x"33",
          1449 => x"a0",
          1450 => x"73",
          1451 => x"f5",
          1452 => x"2e",
          1453 => x"d0",
          1454 => x"56",
          1455 => x"80",
          1456 => x"58",
          1457 => x"74",
          1458 => x"38",
          1459 => x"27",
          1460 => x"14",
          1461 => x"06",
          1462 => x"14",
          1463 => x"06",
          1464 => x"73",
          1465 => x"f9",
          1466 => x"ff",
          1467 => x"89",
          1468 => x"89",
          1469 => x"27",
          1470 => x"77",
          1471 => x"81",
          1472 => x"0c",
          1473 => x"56",
          1474 => x"26",
          1475 => x"78",
          1476 => x"38",
          1477 => x"75",
          1478 => x"56",
          1479 => x"84",
          1480 => x"0d",
          1481 => x"16",
          1482 => x"70",
          1483 => x"59",
          1484 => x"09",
          1485 => x"ff",
          1486 => x"70",
          1487 => x"33",
          1488 => x"80",
          1489 => x"38",
          1490 => x"80",
          1491 => x"38",
          1492 => x"74",
          1493 => x"d0",
          1494 => x"56",
          1495 => x"73",
          1496 => x"38",
          1497 => x"84",
          1498 => x"0d",
          1499 => x"81",
          1500 => x"0c",
          1501 => x"55",
          1502 => x"ca",
          1503 => x"84",
          1504 => x"8b",
          1505 => x"f7",
          1506 => x"7d",
          1507 => x"70",
          1508 => x"08",
          1509 => x"56",
          1510 => x"2e",
          1511 => x"8f",
          1512 => x"70",
          1513 => x"33",
          1514 => x"a0",
          1515 => x"73",
          1516 => x"f5",
          1517 => x"2e",
          1518 => x"d0",
          1519 => x"56",
          1520 => x"80",
          1521 => x"58",
          1522 => x"74",
          1523 => x"38",
          1524 => x"27",
          1525 => x"14",
          1526 => x"06",
          1527 => x"14",
          1528 => x"06",
          1529 => x"73",
          1530 => x"f9",
          1531 => x"ff",
          1532 => x"89",
          1533 => x"89",
          1534 => x"27",
          1535 => x"77",
          1536 => x"81",
          1537 => x"0c",
          1538 => x"56",
          1539 => x"26",
          1540 => x"78",
          1541 => x"38",
          1542 => x"75",
          1543 => x"56",
          1544 => x"84",
          1545 => x"0d",
          1546 => x"16",
          1547 => x"70",
          1548 => x"59",
          1549 => x"09",
          1550 => x"ff",
          1551 => x"70",
          1552 => x"33",
          1553 => x"80",
          1554 => x"38",
          1555 => x"80",
          1556 => x"38",
          1557 => x"74",
          1558 => x"d0",
          1559 => x"56",
          1560 => x"73",
          1561 => x"38",
          1562 => x"84",
          1563 => x"0d",
          1564 => x"81",
          1565 => x"0c",
          1566 => x"55",
          1567 => x"ca",
          1568 => x"84",
          1569 => x"8b",
          1570 => x"80",
          1571 => x"84",
          1572 => x"81",
          1573 => x"bb",
          1574 => x"ff",
          1575 => x"52",
          1576 => x"8c",
          1577 => x"10",
          1578 => x"05",
          1579 => x"04",
          1580 => x"51",
          1581 => x"83",
          1582 => x"83",
          1583 => x"ef",
          1584 => x"3d",
          1585 => x"cf",
          1586 => x"a8",
          1587 => x"0d",
          1588 => x"ec",
          1589 => x"3f",
          1590 => x"04",
          1591 => x"51",
          1592 => x"83",
          1593 => x"83",
          1594 => x"ef",
          1595 => x"3d",
          1596 => x"d0",
          1597 => x"fc",
          1598 => x"0d",
          1599 => x"c4",
          1600 => x"3f",
          1601 => x"04",
          1602 => x"51",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ee",
          1606 => x"3d",
          1607 => x"d1",
          1608 => x"d0",
          1609 => x"0d",
          1610 => x"b4",
          1611 => x"3f",
          1612 => x"04",
          1613 => x"51",
          1614 => x"83",
          1615 => x"83",
          1616 => x"ee",
          1617 => x"3d",
          1618 => x"d1",
          1619 => x"a4",
          1620 => x"0d",
          1621 => x"88",
          1622 => x"3f",
          1623 => x"04",
          1624 => x"51",
          1625 => x"83",
          1626 => x"83",
          1627 => x"ee",
          1628 => x"3d",
          1629 => x"d2",
          1630 => x"f8",
          1631 => x"0d",
          1632 => x"c8",
          1633 => x"3f",
          1634 => x"04",
          1635 => x"51",
          1636 => x"83",
          1637 => x"fe",
          1638 => x"81",
          1639 => x"02",
          1640 => x"e3",
          1641 => x"58",
          1642 => x"99",
          1643 => x"30",
          1644 => x"73",
          1645 => x"57",
          1646 => x"75",
          1647 => x"83",
          1648 => x"74",
          1649 => x"81",
          1650 => x"55",
          1651 => x"80",
          1652 => x"53",
          1653 => x"3d",
          1654 => x"82",
          1655 => x"84",
          1656 => x"57",
          1657 => x"08",
          1658 => x"d1",
          1659 => x"82",
          1660 => x"76",
          1661 => x"07",
          1662 => x"30",
          1663 => x"72",
          1664 => x"57",
          1665 => x"2e",
          1666 => x"c0",
          1667 => x"55",
          1668 => x"26",
          1669 => x"74",
          1670 => x"e8",
          1671 => x"86",
          1672 => x"84",
          1673 => x"d3",
          1674 => x"52",
          1675 => x"51",
          1676 => x"76",
          1677 => x"0c",
          1678 => x"0d",
          1679 => x"84",
          1680 => x"98",
          1681 => x"bb",
          1682 => x"81",
          1683 => x"d4",
          1684 => x"80",
          1685 => x"77",
          1686 => x"ea",
          1687 => x"84",
          1688 => x"bb",
          1689 => x"85",
          1690 => x"74",
          1691 => x"fd",
          1692 => x"75",
          1693 => x"d3",
          1694 => x"52",
          1695 => x"a6",
          1696 => x"84",
          1697 => x"51",
          1698 => x"84",
          1699 => x"54",
          1700 => x"53",
          1701 => x"d2",
          1702 => x"ed",
          1703 => x"39",
          1704 => x"7c",
          1705 => x"b7",
          1706 => x"59",
          1707 => x"53",
          1708 => x"51",
          1709 => x"84",
          1710 => x"8b",
          1711 => x"2e",
          1712 => x"81",
          1713 => x"77",
          1714 => x"0c",
          1715 => x"04",
          1716 => x"e6",
          1717 => x"55",
          1718 => x"bb",
          1719 => x"52",
          1720 => x"2d",
          1721 => x"08",
          1722 => x"0c",
          1723 => x"04",
          1724 => x"7f",
          1725 => x"8c",
          1726 => x"05",
          1727 => x"15",
          1728 => x"5c",
          1729 => x"5e",
          1730 => x"83",
          1731 => x"52",
          1732 => x"51",
          1733 => x"83",
          1734 => x"dd",
          1735 => x"54",
          1736 => x"b2",
          1737 => x"2e",
          1738 => x"7c",
          1739 => x"a8",
          1740 => x"53",
          1741 => x"81",
          1742 => x"33",
          1743 => x"98",
          1744 => x"3f",
          1745 => x"e6",
          1746 => x"54",
          1747 => x"9f",
          1748 => x"26",
          1749 => x"d3",
          1750 => x"ad",
          1751 => x"75",
          1752 => x"c0",
          1753 => x"70",
          1754 => x"80",
          1755 => x"27",
          1756 => x"55",
          1757 => x"74",
          1758 => x"81",
          1759 => x"06",
          1760 => x"06",
          1761 => x"80",
          1762 => x"80",
          1763 => x"81",
          1764 => x"e6",
          1765 => x"a0",
          1766 => x"3f",
          1767 => x"78",
          1768 => x"38",
          1769 => x"51",
          1770 => x"78",
          1771 => x"5c",
          1772 => x"9d",
          1773 => x"bb",
          1774 => x"2b",
          1775 => x"58",
          1776 => x"2e",
          1777 => x"76",
          1778 => x"c3",
          1779 => x"57",
          1780 => x"fe",
          1781 => x"0b",
          1782 => x"0c",
          1783 => x"04",
          1784 => x"51",
          1785 => x"81",
          1786 => x"e8",
          1787 => x"a0",
          1788 => x"3f",
          1789 => x"fe",
          1790 => x"da",
          1791 => x"b8",
          1792 => x"3f",
          1793 => x"e6",
          1794 => x"54",
          1795 => x"df",
          1796 => x"27",
          1797 => x"73",
          1798 => x"7a",
          1799 => x"72",
          1800 => x"d3",
          1801 => x"e1",
          1802 => x"84",
          1803 => x"53",
          1804 => x"ea",
          1805 => x"74",
          1806 => x"fe",
          1807 => x"d3",
          1808 => x"c5",
          1809 => x"84",
          1810 => x"53",
          1811 => x"ea",
          1812 => x"79",
          1813 => x"38",
          1814 => x"72",
          1815 => x"38",
          1816 => x"83",
          1817 => x"db",
          1818 => x"14",
          1819 => x"08",
          1820 => x"51",
          1821 => x"78",
          1822 => x"38",
          1823 => x"84",
          1824 => x"52",
          1825 => x"e7",
          1826 => x"56",
          1827 => x"80",
          1828 => x"84",
          1829 => x"81",
          1830 => x"88",
          1831 => x"2e",
          1832 => x"a0",
          1833 => x"d0",
          1834 => x"06",
          1835 => x"90",
          1836 => x"39",
          1837 => x"c5",
          1838 => x"84",
          1839 => x"70",
          1840 => x"a0",
          1841 => x"72",
          1842 => x"30",
          1843 => x"73",
          1844 => x"51",
          1845 => x"57",
          1846 => x"80",
          1847 => x"38",
          1848 => x"99",
          1849 => x"84",
          1850 => x"70",
          1851 => x"a0",
          1852 => x"72",
          1853 => x"30",
          1854 => x"73",
          1855 => x"51",
          1856 => x"57",
          1857 => x"73",
          1858 => x"38",
          1859 => x"80",
          1860 => x"84",
          1861 => x"0d",
          1862 => x"0d",
          1863 => x"80",
          1864 => x"dd",
          1865 => x"9d",
          1866 => x"d4",
          1867 => x"9e",
          1868 => x"9d",
          1869 => x"81",
          1870 => x"06",
          1871 => x"82",
          1872 => x"82",
          1873 => x"06",
          1874 => x"82",
          1875 => x"83",
          1876 => x"06",
          1877 => x"81",
          1878 => x"84",
          1879 => x"06",
          1880 => x"81",
          1881 => x"85",
          1882 => x"06",
          1883 => x"80",
          1884 => x"86",
          1885 => x"06",
          1886 => x"80",
          1887 => x"87",
          1888 => x"06",
          1889 => x"a9",
          1890 => x"2a",
          1891 => x"72",
          1892 => x"f5",
          1893 => x"0d",
          1894 => x"9c",
          1895 => x"d4",
          1896 => x"aa",
          1897 => x"9c",
          1898 => x"dd",
          1899 => x"0d",
          1900 => x"9c",
          1901 => x"d4",
          1902 => x"92",
          1903 => x"9b",
          1904 => x"88",
          1905 => x"53",
          1906 => x"c6",
          1907 => x"81",
          1908 => x"3f",
          1909 => x"51",
          1910 => x"80",
          1911 => x"3f",
          1912 => x"70",
          1913 => x"52",
          1914 => x"ff",
          1915 => x"39",
          1916 => x"c2",
          1917 => x"a4",
          1918 => x"3f",
          1919 => x"b6",
          1920 => x"2a",
          1921 => x"51",
          1922 => x"2e",
          1923 => x"ff",
          1924 => x"51",
          1925 => x"83",
          1926 => x"9b",
          1927 => x"51",
          1928 => x"72",
          1929 => x"81",
          1930 => x"71",
          1931 => x"c2",
          1932 => x"39",
          1933 => x"fe",
          1934 => x"cc",
          1935 => x"3f",
          1936 => x"f2",
          1937 => x"2a",
          1938 => x"51",
          1939 => x"2e",
          1940 => x"ff",
          1941 => x"51",
          1942 => x"83",
          1943 => x"9a",
          1944 => x"51",
          1945 => x"72",
          1946 => x"81",
          1947 => x"71",
          1948 => x"e6",
          1949 => x"39",
          1950 => x"ba",
          1951 => x"f0",
          1952 => x"3f",
          1953 => x"ae",
          1954 => x"2a",
          1955 => x"51",
          1956 => x"2e",
          1957 => x"ff",
          1958 => x"3d",
          1959 => x"41",
          1960 => x"84",
          1961 => x"42",
          1962 => x"51",
          1963 => x"3f",
          1964 => x"08",
          1965 => x"9b",
          1966 => x"78",
          1967 => x"b5",
          1968 => x"c4",
          1969 => x"3f",
          1970 => x"83",
          1971 => x"d6",
          1972 => x"48",
          1973 => x"80",
          1974 => x"eb",
          1975 => x"0b",
          1976 => x"33",
          1977 => x"06",
          1978 => x"80",
          1979 => x"38",
          1980 => x"83",
          1981 => x"81",
          1982 => x"7d",
          1983 => x"c1",
          1984 => x"5a",
          1985 => x"2e",
          1986 => x"79",
          1987 => x"a0",
          1988 => x"06",
          1989 => x"1a",
          1990 => x"5a",
          1991 => x"f6",
          1992 => x"7b",
          1993 => x"38",
          1994 => x"83",
          1995 => x"70",
          1996 => x"e7",
          1997 => x"bb",
          1998 => x"bb",
          1999 => x"7a",
          2000 => x"52",
          2001 => x"3f",
          2002 => x"08",
          2003 => x"1b",
          2004 => x"81",
          2005 => x"38",
          2006 => x"81",
          2007 => x"5b",
          2008 => x"c4",
          2009 => x"33",
          2010 => x"2e",
          2011 => x"80",
          2012 => x"51",
          2013 => x"84",
          2014 => x"5e",
          2015 => x"08",
          2016 => x"ce",
          2017 => x"84",
          2018 => x"3d",
          2019 => x"51",
          2020 => x"84",
          2021 => x"60",
          2022 => x"5c",
          2023 => x"81",
          2024 => x"bb",
          2025 => x"e7",
          2026 => x"bb",
          2027 => x"26",
          2028 => x"81",
          2029 => x"5e",
          2030 => x"2e",
          2031 => x"7a",
          2032 => x"e7",
          2033 => x"2e",
          2034 => x"7b",
          2035 => x"83",
          2036 => x"7c",
          2037 => x"3f",
          2038 => x"58",
          2039 => x"57",
          2040 => x"55",
          2041 => x"80",
          2042 => x"80",
          2043 => x"51",
          2044 => x"84",
          2045 => x"84",
          2046 => x"09",
          2047 => x"72",
          2048 => x"51",
          2049 => x"80",
          2050 => x"26",
          2051 => x"5a",
          2052 => x"59",
          2053 => x"8d",
          2054 => x"70",
          2055 => x"5c",
          2056 => x"95",
          2057 => x"32",
          2058 => x"07",
          2059 => x"f2",
          2060 => x"2e",
          2061 => x"7d",
          2062 => x"9e",
          2063 => x"fc",
          2064 => x"3f",
          2065 => x"f8",
          2066 => x"7e",
          2067 => x"3f",
          2068 => x"ef",
          2069 => x"81",
          2070 => x"59",
          2071 => x"38",
          2072 => x"d6",
          2073 => x"de",
          2074 => x"8a",
          2075 => x"bb",
          2076 => x"c5",
          2077 => x"0b",
          2078 => x"f8",
          2079 => x"94",
          2080 => x"52",
          2081 => x"f7",
          2082 => x"bb",
          2083 => x"2e",
          2084 => x"bb",
          2085 => x"df",
          2086 => x"0b",
          2087 => x"33",
          2088 => x"06",
          2089 => x"82",
          2090 => x"06",
          2091 => x"91",
          2092 => x"94",
          2093 => x"d2",
          2094 => x"0b",
          2095 => x"f8",
          2096 => x"83",
          2097 => x"80",
          2098 => x"52",
          2099 => x"d7",
          2100 => x"5a",
          2101 => x"b3",
          2102 => x"7c",
          2103 => x"85",
          2104 => x"78",
          2105 => x"fc",
          2106 => x"10",
          2107 => x"e4",
          2108 => x"08",
          2109 => x"83",
          2110 => x"7e",
          2111 => x"3f",
          2112 => x"52",
          2113 => x"51",
          2114 => x"3f",
          2115 => x"08",
          2116 => x"81",
          2117 => x"38",
          2118 => x"3d",
          2119 => x"fb",
          2120 => x"d7",
          2121 => x"cc",
          2122 => x"81",
          2123 => x"fe",
          2124 => x"d7",
          2125 => x"55",
          2126 => x"54",
          2127 => x"d7",
          2128 => x"51",
          2129 => x"fd",
          2130 => x"8d",
          2131 => x"fb",
          2132 => x"3f",
          2133 => x"81",
          2134 => x"80",
          2135 => x"fa",
          2136 => x"8f",
          2137 => x"e3",
          2138 => x"b4",
          2139 => x"3f",
          2140 => x"04",
          2141 => x"51",
          2142 => x"d0",
          2143 => x"cb",
          2144 => x"ff",
          2145 => x"ff",
          2146 => x"eb",
          2147 => x"bb",
          2148 => x"2e",
          2149 => x"68",
          2150 => x"e4",
          2151 => x"3f",
          2152 => x"2d",
          2153 => x"08",
          2154 => x"9f",
          2155 => x"84",
          2156 => x"d8",
          2157 => x"d1",
          2158 => x"39",
          2159 => x"84",
          2160 => x"80",
          2161 => x"bf",
          2162 => x"84",
          2163 => x"f9",
          2164 => x"52",
          2165 => x"51",
          2166 => x"68",
          2167 => x"b8",
          2168 => x"11",
          2169 => x"05",
          2170 => x"3f",
          2171 => x"08",
          2172 => x"d7",
          2173 => x"fe",
          2174 => x"ff",
          2175 => x"e9",
          2176 => x"bb",
          2177 => x"d0",
          2178 => x"78",
          2179 => x"52",
          2180 => x"51",
          2181 => x"84",
          2182 => x"53",
          2183 => x"7e",
          2184 => x"3f",
          2185 => x"33",
          2186 => x"2e",
          2187 => x"78",
          2188 => x"d3",
          2189 => x"05",
          2190 => x"cf",
          2191 => x"fe",
          2192 => x"ff",
          2193 => x"e8",
          2194 => x"bb",
          2195 => x"2e",
          2196 => x"b8",
          2197 => x"11",
          2198 => x"05",
          2199 => x"3f",
          2200 => x"08",
          2201 => x"64",
          2202 => x"53",
          2203 => x"d8",
          2204 => x"95",
          2205 => x"e4",
          2206 => x"f8",
          2207 => x"cf",
          2208 => x"48",
          2209 => x"78",
          2210 => x"bf",
          2211 => x"26",
          2212 => x"64",
          2213 => x"46",
          2214 => x"b8",
          2215 => x"11",
          2216 => x"05",
          2217 => x"3f",
          2218 => x"08",
          2219 => x"9b",
          2220 => x"fe",
          2221 => x"ff",
          2222 => x"e9",
          2223 => x"bb",
          2224 => x"2e",
          2225 => x"b8",
          2226 => x"11",
          2227 => x"05",
          2228 => x"3f",
          2229 => x"08",
          2230 => x"ef",
          2231 => x"d4",
          2232 => x"3f",
          2233 => x"59",
          2234 => x"83",
          2235 => x"70",
          2236 => x"5f",
          2237 => x"7d",
          2238 => x"7a",
          2239 => x"78",
          2240 => x"52",
          2241 => x"51",
          2242 => x"66",
          2243 => x"81",
          2244 => x"47",
          2245 => x"b8",
          2246 => x"11",
          2247 => x"05",
          2248 => x"3f",
          2249 => x"08",
          2250 => x"9f",
          2251 => x"fe",
          2252 => x"ff",
          2253 => x"e8",
          2254 => x"bb",
          2255 => x"2e",
          2256 => x"b8",
          2257 => x"11",
          2258 => x"05",
          2259 => x"3f",
          2260 => x"08",
          2261 => x"f3",
          2262 => x"80",
          2263 => x"3f",
          2264 => x"67",
          2265 => x"38",
          2266 => x"70",
          2267 => x"33",
          2268 => x"81",
          2269 => x"39",
          2270 => x"84",
          2271 => x"80",
          2272 => x"83",
          2273 => x"84",
          2274 => x"f6",
          2275 => x"3d",
          2276 => x"53",
          2277 => x"51",
          2278 => x"84",
          2279 => x"b1",
          2280 => x"33",
          2281 => x"d9",
          2282 => x"dd",
          2283 => x"e4",
          2284 => x"f8",
          2285 => x"cc",
          2286 => x"48",
          2287 => x"78",
          2288 => x"87",
          2289 => x"26",
          2290 => x"68",
          2291 => x"d1",
          2292 => x"02",
          2293 => x"33",
          2294 => x"81",
          2295 => x"3d",
          2296 => x"53",
          2297 => x"51",
          2298 => x"84",
          2299 => x"80",
          2300 => x"38",
          2301 => x"80",
          2302 => x"79",
          2303 => x"05",
          2304 => x"fe",
          2305 => x"ff",
          2306 => x"e6",
          2307 => x"bb",
          2308 => x"bd",
          2309 => x"39",
          2310 => x"84",
          2311 => x"80",
          2312 => x"e3",
          2313 => x"84",
          2314 => x"f5",
          2315 => x"3d",
          2316 => x"53",
          2317 => x"51",
          2318 => x"84",
          2319 => x"80",
          2320 => x"38",
          2321 => x"f8",
          2322 => x"80",
          2323 => x"b7",
          2324 => x"84",
          2325 => x"84",
          2326 => x"46",
          2327 => x"51",
          2328 => x"68",
          2329 => x"78",
          2330 => x"38",
          2331 => x"79",
          2332 => x"5b",
          2333 => x"26",
          2334 => x"51",
          2335 => x"f4",
          2336 => x"3d",
          2337 => x"51",
          2338 => x"84",
          2339 => x"b9",
          2340 => x"05",
          2341 => x"f3",
          2342 => x"84",
          2343 => x"52",
          2344 => x"f3",
          2345 => x"84",
          2346 => x"f4",
          2347 => x"bb",
          2348 => x"e7",
          2349 => x"93",
          2350 => x"ff",
          2351 => x"ff",
          2352 => x"e5",
          2353 => x"bb",
          2354 => x"38",
          2355 => x"33",
          2356 => x"2e",
          2357 => x"83",
          2358 => x"49",
          2359 => x"fc",
          2360 => x"80",
          2361 => x"9f",
          2362 => x"84",
          2363 => x"83",
          2364 => x"5a",
          2365 => x"83",
          2366 => x"f3",
          2367 => x"b8",
          2368 => x"11",
          2369 => x"05",
          2370 => x"3f",
          2371 => x"08",
          2372 => x"38",
          2373 => x"5c",
          2374 => x"83",
          2375 => x"7a",
          2376 => x"30",
          2377 => x"9f",
          2378 => x"5c",
          2379 => x"80",
          2380 => x"7a",
          2381 => x"38",
          2382 => x"d9",
          2383 => x"b4",
          2384 => x"68",
          2385 => x"66",
          2386 => x"eb",
          2387 => x"d9",
          2388 => x"a0",
          2389 => x"39",
          2390 => x"0c",
          2391 => x"05",
          2392 => x"fe",
          2393 => x"ff",
          2394 => x"e2",
          2395 => x"bb",
          2396 => x"2e",
          2397 => x"64",
          2398 => x"59",
          2399 => x"45",
          2400 => x"f0",
          2401 => x"80",
          2402 => x"f7",
          2403 => x"84",
          2404 => x"f2",
          2405 => x"5e",
          2406 => x"05",
          2407 => x"82",
          2408 => x"7d",
          2409 => x"fe",
          2410 => x"ff",
          2411 => x"e1",
          2412 => x"bb",
          2413 => x"2e",
          2414 => x"64",
          2415 => x"ce",
          2416 => x"70",
          2417 => x"23",
          2418 => x"3d",
          2419 => x"53",
          2420 => x"51",
          2421 => x"84",
          2422 => x"ff",
          2423 => x"eb",
          2424 => x"fe",
          2425 => x"ff",
          2426 => x"e3",
          2427 => x"bb",
          2428 => x"2e",
          2429 => x"68",
          2430 => x"db",
          2431 => x"34",
          2432 => x"49",
          2433 => x"b8",
          2434 => x"11",
          2435 => x"05",
          2436 => x"3f",
          2437 => x"08",
          2438 => x"98",
          2439 => x"71",
          2440 => x"84",
          2441 => x"59",
          2442 => x"7a",
          2443 => x"81",
          2444 => x"38",
          2445 => x"d7",
          2446 => x"53",
          2447 => x"52",
          2448 => x"e5",
          2449 => x"39",
          2450 => x"51",
          2451 => x"f3",
          2452 => x"d9",
          2453 => x"9c",
          2454 => x"39",
          2455 => x"f0",
          2456 => x"80",
          2457 => x"9b",
          2458 => x"84",
          2459 => x"b8",
          2460 => x"02",
          2461 => x"22",
          2462 => x"05",
          2463 => x"45",
          2464 => x"83",
          2465 => x"5c",
          2466 => x"80",
          2467 => x"f3",
          2468 => x"fc",
          2469 => x"f4",
          2470 => x"7b",
          2471 => x"38",
          2472 => x"08",
          2473 => x"39",
          2474 => x"51",
          2475 => x"64",
          2476 => x"39",
          2477 => x"51",
          2478 => x"64",
          2479 => x"39",
          2480 => x"33",
          2481 => x"2e",
          2482 => x"f3",
          2483 => x"fc",
          2484 => x"d9",
          2485 => x"9c",
          2486 => x"39",
          2487 => x"33",
          2488 => x"2e",
          2489 => x"f3",
          2490 => x"fc",
          2491 => x"f4",
          2492 => x"7d",
          2493 => x"38",
          2494 => x"08",
          2495 => x"39",
          2496 => x"33",
          2497 => x"2e",
          2498 => x"f3",
          2499 => x"fb",
          2500 => x"f4",
          2501 => x"7c",
          2502 => x"38",
          2503 => x"08",
          2504 => x"39",
          2505 => x"33",
          2506 => x"2e",
          2507 => x"f3",
          2508 => x"fb",
          2509 => x"f3",
          2510 => x"80",
          2511 => x"9c",
          2512 => x"f0",
          2513 => x"47",
          2514 => x"f3",
          2515 => x"0b",
          2516 => x"34",
          2517 => x"8c",
          2518 => x"57",
          2519 => x"52",
          2520 => x"c2",
          2521 => x"84",
          2522 => x"77",
          2523 => x"87",
          2524 => x"75",
          2525 => x"3f",
          2526 => x"84",
          2527 => x"0c",
          2528 => x"9c",
          2529 => x"57",
          2530 => x"52",
          2531 => x"96",
          2532 => x"84",
          2533 => x"77",
          2534 => x"87",
          2535 => x"75",
          2536 => x"3f",
          2537 => x"84",
          2538 => x"0c",
          2539 => x"0b",
          2540 => x"84",
          2541 => x"83",
          2542 => x"94",
          2543 => x"be",
          2544 => x"c9",
          2545 => x"02",
          2546 => x"05",
          2547 => x"84",
          2548 => x"89",
          2549 => x"13",
          2550 => x"0c",
          2551 => x"0c",
          2552 => x"3f",
          2553 => x"95",
          2554 => x"98",
          2555 => x"3f",
          2556 => x"52",
          2557 => x"51",
          2558 => x"83",
          2559 => x"22",
          2560 => x"98",
          2561 => x"cc",
          2562 => x"d8",
          2563 => x"33",
          2564 => x"e0",
          2565 => x"3f",
          2566 => x"83",
          2567 => x"d0",
          2568 => x"52",
          2569 => x"51",
          2570 => x"90",
          2571 => x"83",
          2572 => x"c3",
          2573 => x"e2",
          2574 => x"fb",
          2575 => x"70",
          2576 => x"80",
          2577 => x"74",
          2578 => x"83",
          2579 => x"70",
          2580 => x"52",
          2581 => x"2e",
          2582 => x"91",
          2583 => x"70",
          2584 => x"ff",
          2585 => x"55",
          2586 => x"f1",
          2587 => x"ff",
          2588 => x"a2",
          2589 => x"38",
          2590 => x"81",
          2591 => x"38",
          2592 => x"70",
          2593 => x"53",
          2594 => x"a0",
          2595 => x"81",
          2596 => x"2e",
          2597 => x"80",
          2598 => x"81",
          2599 => x"39",
          2600 => x"ff",
          2601 => x"70",
          2602 => x"81",
          2603 => x"81",
          2604 => x"32",
          2605 => x"80",
          2606 => x"52",
          2607 => x"80",
          2608 => x"80",
          2609 => x"05",
          2610 => x"76",
          2611 => x"70",
          2612 => x"0c",
          2613 => x"04",
          2614 => x"c4",
          2615 => x"2e",
          2616 => x"81",
          2617 => x"72",
          2618 => x"ff",
          2619 => x"54",
          2620 => x"e4",
          2621 => x"e0",
          2622 => x"55",
          2623 => x"53",
          2624 => x"09",
          2625 => x"f8",
          2626 => x"fc",
          2627 => x"53",
          2628 => x"38",
          2629 => x"bb",
          2630 => x"3d",
          2631 => x"3d",
          2632 => x"72",
          2633 => x"3f",
          2634 => x"08",
          2635 => x"38",
          2636 => x"84",
          2637 => x"0d",
          2638 => x"0d",
          2639 => x"33",
          2640 => x"53",
          2641 => x"8b",
          2642 => x"38",
          2643 => x"ff",
          2644 => x"52",
          2645 => x"81",
          2646 => x"13",
          2647 => x"52",
          2648 => x"80",
          2649 => x"13",
          2650 => x"52",
          2651 => x"80",
          2652 => x"13",
          2653 => x"52",
          2654 => x"80",
          2655 => x"13",
          2656 => x"52",
          2657 => x"26",
          2658 => x"8a",
          2659 => x"87",
          2660 => x"e7",
          2661 => x"38",
          2662 => x"c0",
          2663 => x"72",
          2664 => x"98",
          2665 => x"13",
          2666 => x"98",
          2667 => x"13",
          2668 => x"98",
          2669 => x"13",
          2670 => x"98",
          2671 => x"13",
          2672 => x"98",
          2673 => x"13",
          2674 => x"98",
          2675 => x"87",
          2676 => x"0c",
          2677 => x"98",
          2678 => x"0b",
          2679 => x"9c",
          2680 => x"71",
          2681 => x"0c",
          2682 => x"04",
          2683 => x"7f",
          2684 => x"98",
          2685 => x"7d",
          2686 => x"98",
          2687 => x"7d",
          2688 => x"c0",
          2689 => x"5c",
          2690 => x"34",
          2691 => x"b4",
          2692 => x"83",
          2693 => x"c0",
          2694 => x"5c",
          2695 => x"34",
          2696 => x"ac",
          2697 => x"85",
          2698 => x"c0",
          2699 => x"5c",
          2700 => x"34",
          2701 => x"a4",
          2702 => x"88",
          2703 => x"c0",
          2704 => x"5a",
          2705 => x"23",
          2706 => x"79",
          2707 => x"06",
          2708 => x"ff",
          2709 => x"86",
          2710 => x"85",
          2711 => x"84",
          2712 => x"83",
          2713 => x"82",
          2714 => x"7d",
          2715 => x"06",
          2716 => x"fc",
          2717 => x"91",
          2718 => x"0d",
          2719 => x"0d",
          2720 => x"33",
          2721 => x"2e",
          2722 => x"51",
          2723 => x"3f",
          2724 => x"08",
          2725 => x"98",
          2726 => x"71",
          2727 => x"81",
          2728 => x"72",
          2729 => x"38",
          2730 => x"84",
          2731 => x"0d",
          2732 => x"80",
          2733 => x"84",
          2734 => x"98",
          2735 => x"2c",
          2736 => x"ff",
          2737 => x"06",
          2738 => x"51",
          2739 => x"3f",
          2740 => x"08",
          2741 => x"98",
          2742 => x"71",
          2743 => x"38",
          2744 => x"3d",
          2745 => x"54",
          2746 => x"2b",
          2747 => x"80",
          2748 => x"84",
          2749 => x"98",
          2750 => x"2c",
          2751 => x"ff",
          2752 => x"73",
          2753 => x"14",
          2754 => x"73",
          2755 => x"71",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"02",
          2759 => x"83",
          2760 => x"70",
          2761 => x"53",
          2762 => x"80",
          2763 => x"38",
          2764 => x"94",
          2765 => x"2a",
          2766 => x"53",
          2767 => x"80",
          2768 => x"71",
          2769 => x"81",
          2770 => x"70",
          2771 => x"81",
          2772 => x"53",
          2773 => x"8a",
          2774 => x"2a",
          2775 => x"71",
          2776 => x"81",
          2777 => x"87",
          2778 => x"52",
          2779 => x"86",
          2780 => x"94",
          2781 => x"72",
          2782 => x"bb",
          2783 => x"3d",
          2784 => x"91",
          2785 => x"06",
          2786 => x"97",
          2787 => x"32",
          2788 => x"72",
          2789 => x"38",
          2790 => x"81",
          2791 => x"80",
          2792 => x"87",
          2793 => x"08",
          2794 => x"70",
          2795 => x"54",
          2796 => x"38",
          2797 => x"3d",
          2798 => x"05",
          2799 => x"70",
          2800 => x"52",
          2801 => x"f3",
          2802 => x"3d",
          2803 => x"3d",
          2804 => x"80",
          2805 => x"56",
          2806 => x"77",
          2807 => x"38",
          2808 => x"f3",
          2809 => x"81",
          2810 => x"57",
          2811 => x"2e",
          2812 => x"87",
          2813 => x"08",
          2814 => x"70",
          2815 => x"54",
          2816 => x"2e",
          2817 => x"91",
          2818 => x"06",
          2819 => x"e3",
          2820 => x"32",
          2821 => x"72",
          2822 => x"38",
          2823 => x"81",
          2824 => x"cf",
          2825 => x"ff",
          2826 => x"c0",
          2827 => x"70",
          2828 => x"38",
          2829 => x"90",
          2830 => x"0c",
          2831 => x"33",
          2832 => x"ff",
          2833 => x"84",
          2834 => x"88",
          2835 => x"71",
          2836 => x"81",
          2837 => x"70",
          2838 => x"81",
          2839 => x"53",
          2840 => x"c1",
          2841 => x"2a",
          2842 => x"71",
          2843 => x"b5",
          2844 => x"94",
          2845 => x"96",
          2846 => x"06",
          2847 => x"70",
          2848 => x"39",
          2849 => x"87",
          2850 => x"08",
          2851 => x"8a",
          2852 => x"70",
          2853 => x"ab",
          2854 => x"9e",
          2855 => x"f3",
          2856 => x"c0",
          2857 => x"83",
          2858 => x"87",
          2859 => x"08",
          2860 => x"0c",
          2861 => x"98",
          2862 => x"cc",
          2863 => x"9e",
          2864 => x"f3",
          2865 => x"c0",
          2866 => x"83",
          2867 => x"87",
          2868 => x"08",
          2869 => x"0c",
          2870 => x"b0",
          2871 => x"dc",
          2872 => x"9e",
          2873 => x"f3",
          2874 => x"c0",
          2875 => x"83",
          2876 => x"87",
          2877 => x"08",
          2878 => x"0c",
          2879 => x"c0",
          2880 => x"ec",
          2881 => x"9e",
          2882 => x"f3",
          2883 => x"c0",
          2884 => x"52",
          2885 => x"f4",
          2886 => x"9e",
          2887 => x"f3",
          2888 => x"c0",
          2889 => x"83",
          2890 => x"87",
          2891 => x"08",
          2892 => x"0c",
          2893 => x"f4",
          2894 => x"0b",
          2895 => x"90",
          2896 => x"80",
          2897 => x"52",
          2898 => x"fb",
          2899 => x"f4",
          2900 => x"0b",
          2901 => x"90",
          2902 => x"80",
          2903 => x"52",
          2904 => x"2e",
          2905 => x"52",
          2906 => x"86",
          2907 => x"87",
          2908 => x"08",
          2909 => x"0a",
          2910 => x"52",
          2911 => x"83",
          2912 => x"71",
          2913 => x"34",
          2914 => x"c0",
          2915 => x"70",
          2916 => x"06",
          2917 => x"70",
          2918 => x"38",
          2919 => x"83",
          2920 => x"80",
          2921 => x"9e",
          2922 => x"a0",
          2923 => x"51",
          2924 => x"80",
          2925 => x"81",
          2926 => x"f4",
          2927 => x"0b",
          2928 => x"90",
          2929 => x"80",
          2930 => x"52",
          2931 => x"2e",
          2932 => x"52",
          2933 => x"8a",
          2934 => x"87",
          2935 => x"08",
          2936 => x"80",
          2937 => x"52",
          2938 => x"83",
          2939 => x"71",
          2940 => x"34",
          2941 => x"c0",
          2942 => x"70",
          2943 => x"06",
          2944 => x"70",
          2945 => x"38",
          2946 => x"83",
          2947 => x"80",
          2948 => x"9e",
          2949 => x"81",
          2950 => x"51",
          2951 => x"80",
          2952 => x"81",
          2953 => x"f4",
          2954 => x"0b",
          2955 => x"90",
          2956 => x"c0",
          2957 => x"52",
          2958 => x"2e",
          2959 => x"52",
          2960 => x"8e",
          2961 => x"87",
          2962 => x"08",
          2963 => x"06",
          2964 => x"70",
          2965 => x"38",
          2966 => x"83",
          2967 => x"87",
          2968 => x"08",
          2969 => x"70",
          2970 => x"51",
          2971 => x"90",
          2972 => x"87",
          2973 => x"08",
          2974 => x"06",
          2975 => x"70",
          2976 => x"38",
          2977 => x"83",
          2978 => x"87",
          2979 => x"08",
          2980 => x"70",
          2981 => x"51",
          2982 => x"92",
          2983 => x"87",
          2984 => x"08",
          2985 => x"51",
          2986 => x"80",
          2987 => x"81",
          2988 => x"f4",
          2989 => x"c0",
          2990 => x"87",
          2991 => x"83",
          2992 => x"83",
          2993 => x"81",
          2994 => x"39",
          2995 => x"83",
          2996 => x"ff",
          2997 => x"83",
          2998 => x"54",
          2999 => x"38",
          3000 => x"51",
          3001 => x"83",
          3002 => x"55",
          3003 => x"38",
          3004 => x"33",
          3005 => x"c7",
          3006 => x"88",
          3007 => x"85",
          3008 => x"f4",
          3009 => x"74",
          3010 => x"83",
          3011 => x"54",
          3012 => x"38",
          3013 => x"33",
          3014 => x"a9",
          3015 => x"93",
          3016 => x"84",
          3017 => x"f4",
          3018 => x"74",
          3019 => x"83",
          3020 => x"56",
          3021 => x"38",
          3022 => x"33",
          3023 => x"a7",
          3024 => x"8c",
          3025 => x"83",
          3026 => x"f4",
          3027 => x"75",
          3028 => x"83",
          3029 => x"54",
          3030 => x"38",
          3031 => x"51",
          3032 => x"83",
          3033 => x"52",
          3034 => x"51",
          3035 => x"3f",
          3036 => x"08",
          3037 => x"f4",
          3038 => x"8d",
          3039 => x"f0",
          3040 => x"db",
          3041 => x"b5",
          3042 => x"db",
          3043 => x"e4",
          3044 => x"f4",
          3045 => x"db",
          3046 => x"b4",
          3047 => x"f3",
          3048 => x"bd",
          3049 => x"75",
          3050 => x"3f",
          3051 => x"08",
          3052 => x"29",
          3053 => x"54",
          3054 => x"84",
          3055 => x"db",
          3056 => x"b4",
          3057 => x"f4",
          3058 => x"74",
          3059 => x"f4",
          3060 => x"74",
          3061 => x"3d",
          3062 => x"f4",
          3063 => x"bd",
          3064 => x"75",
          3065 => x"3f",
          3066 => x"08",
          3067 => x"29",
          3068 => x"54",
          3069 => x"84",
          3070 => x"dc",
          3071 => x"b4",
          3072 => x"3d",
          3073 => x"f3",
          3074 => x"bd",
          3075 => x"75",
          3076 => x"3f",
          3077 => x"08",
          3078 => x"29",
          3079 => x"54",
          3080 => x"84",
          3081 => x"dc",
          3082 => x"b3",
          3083 => x"f4",
          3084 => x"74",
          3085 => x"9e",
          3086 => x"39",
          3087 => x"51",
          3088 => x"83",
          3089 => x"c0",
          3090 => x"f3",
          3091 => x"83",
          3092 => x"ff",
          3093 => x"83",
          3094 => x"52",
          3095 => x"51",
          3096 => x"3f",
          3097 => x"08",
          3098 => x"9c",
          3099 => x"99",
          3100 => x"c4",
          3101 => x"fc",
          3102 => x"f4",
          3103 => x"db",
          3104 => x"b3",
          3105 => x"f3",
          3106 => x"bd",
          3107 => x"75",
          3108 => x"3f",
          3109 => x"08",
          3110 => x"29",
          3111 => x"54",
          3112 => x"84",
          3113 => x"db",
          3114 => x"b2",
          3115 => x"f4",
          3116 => x"74",
          3117 => x"96",
          3118 => x"39",
          3119 => x"51",
          3120 => x"3f",
          3121 => x"33",
          3122 => x"2e",
          3123 => x"fe",
          3124 => x"dd",
          3125 => x"bf",
          3126 => x"f4",
          3127 => x"75",
          3128 => x"ef",
          3129 => x"83",
          3130 => x"ff",
          3131 => x"83",
          3132 => x"55",
          3133 => x"fc",
          3134 => x"39",
          3135 => x"51",
          3136 => x"3f",
          3137 => x"33",
          3138 => x"2e",
          3139 => x"d7",
          3140 => x"92",
          3141 => x"dd",
          3142 => x"b1",
          3143 => x"f4",
          3144 => x"75",
          3145 => x"90",
          3146 => x"83",
          3147 => x"52",
          3148 => x"51",
          3149 => x"3f",
          3150 => x"33",
          3151 => x"2e",
          3152 => x"cd",
          3153 => x"90",
          3154 => x"dd",
          3155 => x"b1",
          3156 => x"f4",
          3157 => x"73",
          3158 => x"ca",
          3159 => x"83",
          3160 => x"83",
          3161 => x"11",
          3162 => x"de",
          3163 => x"b1",
          3164 => x"f4",
          3165 => x"75",
          3166 => x"a1",
          3167 => x"83",
          3168 => x"83",
          3169 => x"11",
          3170 => x"de",
          3171 => x"b0",
          3172 => x"f4",
          3173 => x"73",
          3174 => x"f8",
          3175 => x"83",
          3176 => x"83",
          3177 => x"11",
          3178 => x"de",
          3179 => x"b0",
          3180 => x"f4",
          3181 => x"74",
          3182 => x"cf",
          3183 => x"83",
          3184 => x"83",
          3185 => x"11",
          3186 => x"de",
          3187 => x"b0",
          3188 => x"f4",
          3189 => x"75",
          3190 => x"a6",
          3191 => x"83",
          3192 => x"83",
          3193 => x"11",
          3194 => x"df",
          3195 => x"b0",
          3196 => x"f4",
          3197 => x"73",
          3198 => x"fd",
          3199 => x"83",
          3200 => x"ff",
          3201 => x"83",
          3202 => x"ff",
          3203 => x"83",
          3204 => x"55",
          3205 => x"f9",
          3206 => x"39",
          3207 => x"02",
          3208 => x"52",
          3209 => x"8c",
          3210 => x"10",
          3211 => x"05",
          3212 => x"04",
          3213 => x"51",
          3214 => x"3f",
          3215 => x"04",
          3216 => x"51",
          3217 => x"3f",
          3218 => x"04",
          3219 => x"51",
          3220 => x"3f",
          3221 => x"04",
          3222 => x"51",
          3223 => x"3f",
          3224 => x"04",
          3225 => x"51",
          3226 => x"3f",
          3227 => x"04",
          3228 => x"51",
          3229 => x"3f",
          3230 => x"04",
          3231 => x"0c",
          3232 => x"87",
          3233 => x"0c",
          3234 => x"98",
          3235 => x"96",
          3236 => x"d9",
          3237 => x"3d",
          3238 => x"08",
          3239 => x"70",
          3240 => x"52",
          3241 => x"08",
          3242 => x"fb",
          3243 => x"84",
          3244 => x"38",
          3245 => x"ff",
          3246 => x"ec",
          3247 => x"80",
          3248 => x"51",
          3249 => x"3f",
          3250 => x"08",
          3251 => x"38",
          3252 => x"d5",
          3253 => x"84",
          3254 => x"57",
          3255 => x"84",
          3256 => x"25",
          3257 => x"bb",
          3258 => x"05",
          3259 => x"55",
          3260 => x"74",
          3261 => x"70",
          3262 => x"2a",
          3263 => x"78",
          3264 => x"38",
          3265 => x"38",
          3266 => x"08",
          3267 => x"53",
          3268 => x"93",
          3269 => x"84",
          3270 => x"78",
          3271 => x"38",
          3272 => x"84",
          3273 => x"0d",
          3274 => x"b8",
          3275 => x"d9",
          3276 => x"2e",
          3277 => x"e8",
          3278 => x"79",
          3279 => x"3f",
          3280 => x"bf",
          3281 => x"3d",
          3282 => x"bb",
          3283 => x"34",
          3284 => x"e3",
          3285 => x"ad",
          3286 => x"0b",
          3287 => x"0c",
          3288 => x"04",
          3289 => x"ab",
          3290 => x"3d",
          3291 => x"5d",
          3292 => x"57",
          3293 => x"a0",
          3294 => x"38",
          3295 => x"3d",
          3296 => x"10",
          3297 => x"f4",
          3298 => x"08",
          3299 => x"bf",
          3300 => x"bb",
          3301 => x"79",
          3302 => x"51",
          3303 => x"3f",
          3304 => x"08",
          3305 => x"14",
          3306 => x"81",
          3307 => x"38",
          3308 => x"99",
          3309 => x"70",
          3310 => x"57",
          3311 => x"27",
          3312 => x"54",
          3313 => x"84",
          3314 => x"0d",
          3315 => x"5a",
          3316 => x"84",
          3317 => x"80",
          3318 => x"ab",
          3319 => x"84",
          3320 => x"d1",
          3321 => x"53",
          3322 => x"51",
          3323 => x"84",
          3324 => x"81",
          3325 => x"73",
          3326 => x"38",
          3327 => x"81",
          3328 => x"54",
          3329 => x"fe",
          3330 => x"b6",
          3331 => x"77",
          3332 => x"76",
          3333 => x"38",
          3334 => x"5b",
          3335 => x"55",
          3336 => x"09",
          3337 => x"d4",
          3338 => x"26",
          3339 => x"0b",
          3340 => x"56",
          3341 => x"73",
          3342 => x"08",
          3343 => x"ec",
          3344 => x"82",
          3345 => x"84",
          3346 => x"80",
          3347 => x"f4",
          3348 => x"80",
          3349 => x"51",
          3350 => x"3f",
          3351 => x"08",
          3352 => x"38",
          3353 => x"bd",
          3354 => x"bb",
          3355 => x"80",
          3356 => x"84",
          3357 => x"38",
          3358 => x"08",
          3359 => x"19",
          3360 => x"77",
          3361 => x"75",
          3362 => x"83",
          3363 => x"56",
          3364 => x"3f",
          3365 => x"09",
          3366 => x"b2",
          3367 => x"84",
          3368 => x"aa",
          3369 => x"cd",
          3370 => x"3d",
          3371 => x"08",
          3372 => x"bc",
          3373 => x"3d",
          3374 => x"58",
          3375 => x"0b",
          3376 => x"83",
          3377 => x"5d",
          3378 => x"f0",
          3379 => x"ec",
          3380 => x"9e",
          3381 => x"81",
          3382 => x"57",
          3383 => x"82",
          3384 => x"80",
          3385 => x"38",
          3386 => x"06",
          3387 => x"90",
          3388 => x"80",
          3389 => x"38",
          3390 => x"3d",
          3391 => x"51",
          3392 => x"84",
          3393 => x"98",
          3394 => x"2c",
          3395 => x"ff",
          3396 => x"38",
          3397 => x"06",
          3398 => x"33",
          3399 => x"70",
          3400 => x"e2",
          3401 => x"98",
          3402 => x"2c",
          3403 => x"05",
          3404 => x"83",
          3405 => x"70",
          3406 => x"33",
          3407 => x"5d",
          3408 => x"58",
          3409 => x"57",
          3410 => x"80",
          3411 => x"75",
          3412 => x"38",
          3413 => x"0a",
          3414 => x"0a",
          3415 => x"2c",
          3416 => x"76",
          3417 => x"38",
          3418 => x"70",
          3419 => x"57",
          3420 => x"df",
          3421 => x"43",
          3422 => x"25",
          3423 => x"df",
          3424 => x"18",
          3425 => x"42",
          3426 => x"81",
          3427 => x"80",
          3428 => x"75",
          3429 => x"34",
          3430 => x"80",
          3431 => x"38",
          3432 => x"98",
          3433 => x"2c",
          3434 => x"33",
          3435 => x"70",
          3436 => x"98",
          3437 => x"82",
          3438 => x"e4",
          3439 => x"53",
          3440 => x"5d",
          3441 => x"78",
          3442 => x"38",
          3443 => x"c0",
          3444 => x"e9",
          3445 => x"bb",
          3446 => x"2b",
          3447 => x"5b",
          3448 => x"2e",
          3449 => x"fe",
          3450 => x"80",
          3451 => x"38",
          3452 => x"8a",
          3453 => x"76",
          3454 => x"75",
          3455 => x"29",
          3456 => x"05",
          3457 => x"70",
          3458 => x"59",
          3459 => x"95",
          3460 => x"38",
          3461 => x"70",
          3462 => x"55",
          3463 => x"df",
          3464 => x"43",
          3465 => x"25",
          3466 => x"df",
          3467 => x"18",
          3468 => x"55",
          3469 => x"ff",
          3470 => x"80",
          3471 => x"38",
          3472 => x"81",
          3473 => x"2e",
          3474 => x"fe",
          3475 => x"57",
          3476 => x"80",
          3477 => x"c8",
          3478 => x"e2",
          3479 => x"84",
          3480 => x"79",
          3481 => x"60",
          3482 => x"74",
          3483 => x"8e",
          3484 => x"10",
          3485 => x"05",
          3486 => x"04",
          3487 => x"15",
          3488 => x"80",
          3489 => x"c0",
          3490 => x"84",
          3491 => x"d9",
          3492 => x"c8",
          3493 => x"80",
          3494 => x"38",
          3495 => x"08",
          3496 => x"ff",
          3497 => x"84",
          3498 => x"ff",
          3499 => x"84",
          3500 => x"fc",
          3501 => x"e2",
          3502 => x"81",
          3503 => x"e2",
          3504 => x"57",
          3505 => x"27",
          3506 => x"84",
          3507 => x"52",
          3508 => x"61",
          3509 => x"34",
          3510 => x"33",
          3511 => x"b5",
          3512 => x"9a",
          3513 => x"2e",
          3514 => x"7c",
          3515 => x"38",
          3516 => x"83",
          3517 => x"70",
          3518 => x"75",
          3519 => x"80",
          3520 => x"c4",
          3521 => x"34",
          3522 => x"33",
          3523 => x"33",
          3524 => x"80",
          3525 => x"84",
          3526 => x"52",
          3527 => x"b4",
          3528 => x"e6",
          3529 => x"a0",
          3530 => x"c3",
          3531 => x"e8",
          3532 => x"51",
          3533 => x"3f",
          3534 => x"33",
          3535 => x"78",
          3536 => x"34",
          3537 => x"06",
          3538 => x"38",
          3539 => x"a5",
          3540 => x"84",
          3541 => x"fb",
          3542 => x"8a",
          3543 => x"e8",
          3544 => x"8c",
          3545 => x"1d",
          3546 => x"06",
          3547 => x"92",
          3548 => x"7c",
          3549 => x"f4",
          3550 => x"08",
          3551 => x"8d",
          3552 => x"93",
          3553 => x"38",
          3554 => x"83",
          3555 => x"70",
          3556 => x"75",
          3557 => x"e6",
          3558 => x"ff",
          3559 => x"84",
          3560 => x"84",
          3561 => x"84",
          3562 => x"81",
          3563 => x"05",
          3564 => x"7b",
          3565 => x"b3",
          3566 => x"c4",
          3567 => x"c8",
          3568 => x"74",
          3569 => x"84",
          3570 => x"e8",
          3571 => x"51",
          3572 => x"3f",
          3573 => x"08",
          3574 => x"ff",
          3575 => x"84",
          3576 => x"52",
          3577 => x"b3",
          3578 => x"e2",
          3579 => x"05",
          3580 => x"e2",
          3581 => x"81",
          3582 => x"c7",
          3583 => x"c8",
          3584 => x"ff",
          3585 => x"c4",
          3586 => x"55",
          3587 => x"f9",
          3588 => x"e6",
          3589 => x"81",
          3590 => x"84",
          3591 => x"7b",
          3592 => x"52",
          3593 => x"c7",
          3594 => x"c8",
          3595 => x"ff",
          3596 => x"c4",
          3597 => x"55",
          3598 => x"f9",
          3599 => x"e6",
          3600 => x"81",
          3601 => x"84",
          3602 => x"7b",
          3603 => x"52",
          3604 => x"9b",
          3605 => x"c8",
          3606 => x"ff",
          3607 => x"c4",
          3608 => x"55",
          3609 => x"ff",
          3610 => x"92",
          3611 => x"c8",
          3612 => x"c4",
          3613 => x"74",
          3614 => x"82",
          3615 => x"5b",
          3616 => x"c4",
          3617 => x"2b",
          3618 => x"7c",
          3619 => x"44",
          3620 => x"76",
          3621 => x"38",
          3622 => x"08",
          3623 => x"ff",
          3624 => x"84",
          3625 => x"70",
          3626 => x"98",
          3627 => x"c4",
          3628 => x"43",
          3629 => x"24",
          3630 => x"84",
          3631 => x"52",
          3632 => x"b1",
          3633 => x"81",
          3634 => x"81",
          3635 => x"70",
          3636 => x"e2",
          3637 => x"56",
          3638 => x"24",
          3639 => x"84",
          3640 => x"52",
          3641 => x"b1",
          3642 => x"81",
          3643 => x"81",
          3644 => x"70",
          3645 => x"e2",
          3646 => x"56",
          3647 => x"25",
          3648 => x"f7",
          3649 => x"16",
          3650 => x"33",
          3651 => x"e6",
          3652 => x"77",
          3653 => x"b0",
          3654 => x"81",
          3655 => x"81",
          3656 => x"70",
          3657 => x"e2",
          3658 => x"57",
          3659 => x"25",
          3660 => x"7b",
          3661 => x"18",
          3662 => x"84",
          3663 => x"52",
          3664 => x"ff",
          3665 => x"75",
          3666 => x"29",
          3667 => x"05",
          3668 => x"84",
          3669 => x"5c",
          3670 => x"76",
          3671 => x"38",
          3672 => x"84",
          3673 => x"55",
          3674 => x"f7",
          3675 => x"e6",
          3676 => x"88",
          3677 => x"f7",
          3678 => x"c8",
          3679 => x"57",
          3680 => x"c8",
          3681 => x"ff",
          3682 => x"39",
          3683 => x"33",
          3684 => x"80",
          3685 => x"e6",
          3686 => x"8a",
          3687 => x"cf",
          3688 => x"c4",
          3689 => x"f3",
          3690 => x"bb",
          3691 => x"ff",
          3692 => x"8a",
          3693 => x"e2",
          3694 => x"76",
          3695 => x"f0",
          3696 => x"f4",
          3697 => x"10",
          3698 => x"05",
          3699 => x"41",
          3700 => x"c2",
          3701 => x"2b",
          3702 => x"83",
          3703 => x"81",
          3704 => x"57",
          3705 => x"e2",
          3706 => x"84",
          3707 => x"83",
          3708 => x"70",
          3709 => x"f4",
          3710 => x"08",
          3711 => x"e3",
          3712 => x"ff",
          3713 => x"83",
          3714 => x"70",
          3715 => x"f4",
          3716 => x"08",
          3717 => x"74",
          3718 => x"83",
          3719 => x"56",
          3720 => x"8c",
          3721 => x"f0",
          3722 => x"80",
          3723 => x"38",
          3724 => x"e2",
          3725 => x"0b",
          3726 => x"34",
          3727 => x"84",
          3728 => x"0d",
          3729 => x"c8",
          3730 => x"80",
          3731 => x"84",
          3732 => x"52",
          3733 => x"ae",
          3734 => x"e6",
          3735 => x"a0",
          3736 => x"8b",
          3737 => x"e8",
          3738 => x"51",
          3739 => x"3f",
          3740 => x"33",
          3741 => x"61",
          3742 => x"34",
          3743 => x"06",
          3744 => x"38",
          3745 => x"51",
          3746 => x"3f",
          3747 => x"e2",
          3748 => x"0b",
          3749 => x"34",
          3750 => x"84",
          3751 => x"70",
          3752 => x"5c",
          3753 => x"2e",
          3754 => x"84",
          3755 => x"ff",
          3756 => x"84",
          3757 => x"ff",
          3758 => x"84",
          3759 => x"84",
          3760 => x"52",
          3761 => x"ad",
          3762 => x"e2",
          3763 => x"98",
          3764 => x"2c",
          3765 => x"33",
          3766 => x"56",
          3767 => x"80",
          3768 => x"e6",
          3769 => x"a0",
          3770 => x"83",
          3771 => x"c8",
          3772 => x"2b",
          3773 => x"84",
          3774 => x"5c",
          3775 => x"74",
          3776 => x"fa",
          3777 => x"e8",
          3778 => x"51",
          3779 => x"3f",
          3780 => x"0a",
          3781 => x"0a",
          3782 => x"2c",
          3783 => x"33",
          3784 => x"74",
          3785 => x"d6",
          3786 => x"e8",
          3787 => x"51",
          3788 => x"3f",
          3789 => x"0a",
          3790 => x"0a",
          3791 => x"2c",
          3792 => x"33",
          3793 => x"79",
          3794 => x"b9",
          3795 => x"39",
          3796 => x"81",
          3797 => x"34",
          3798 => x"08",
          3799 => x"51",
          3800 => x"3f",
          3801 => x"0a",
          3802 => x"0a",
          3803 => x"2c",
          3804 => x"33",
          3805 => x"75",
          3806 => x"e6",
          3807 => x"57",
          3808 => x"77",
          3809 => x"e8",
          3810 => x"33",
          3811 => x"df",
          3812 => x"80",
          3813 => x"80",
          3814 => x"98",
          3815 => x"c4",
          3816 => x"5b",
          3817 => x"ff",
          3818 => x"b6",
          3819 => x"34",
          3820 => x"1d",
          3821 => x"c8",
          3822 => x"80",
          3823 => x"84",
          3824 => x"52",
          3825 => x"ab",
          3826 => x"e6",
          3827 => x"a0",
          3828 => x"9b",
          3829 => x"e8",
          3830 => x"51",
          3831 => x"3f",
          3832 => x"33",
          3833 => x"7c",
          3834 => x"34",
          3835 => x"06",
          3836 => x"38",
          3837 => x"51",
          3838 => x"3f",
          3839 => x"e2",
          3840 => x"0b",
          3841 => x"34",
          3842 => x"84",
          3843 => x"0d",
          3844 => x"c8",
          3845 => x"ff",
          3846 => x"76",
          3847 => x"de",
          3848 => x"c4",
          3849 => x"75",
          3850 => x"74",
          3851 => x"98",
          3852 => x"76",
          3853 => x"38",
          3854 => x"7a",
          3855 => x"34",
          3856 => x"0a",
          3857 => x"0a",
          3858 => x"2c",
          3859 => x"33",
          3860 => x"75",
          3861 => x"38",
          3862 => x"74",
          3863 => x"34",
          3864 => x"06",
          3865 => x"b4",
          3866 => x"34",
          3867 => x"33",
          3868 => x"25",
          3869 => x"17",
          3870 => x"e2",
          3871 => x"57",
          3872 => x"33",
          3873 => x"0a",
          3874 => x"0a",
          3875 => x"2c",
          3876 => x"06",
          3877 => x"58",
          3878 => x"81",
          3879 => x"98",
          3880 => x"2c",
          3881 => x"06",
          3882 => x"75",
          3883 => x"ce",
          3884 => x"e8",
          3885 => x"51",
          3886 => x"3f",
          3887 => x"0a",
          3888 => x"0a",
          3889 => x"2c",
          3890 => x"33",
          3891 => x"75",
          3892 => x"aa",
          3893 => x"e8",
          3894 => x"51",
          3895 => x"3f",
          3896 => x"0a",
          3897 => x"0a",
          3898 => x"2c",
          3899 => x"33",
          3900 => x"74",
          3901 => x"b9",
          3902 => x"39",
          3903 => x"80",
          3904 => x"84",
          3905 => x"83",
          3906 => x"84",
          3907 => x"52",
          3908 => x"51",
          3909 => x"3f",
          3910 => x"08",
          3911 => x"a6",
          3912 => x"f4",
          3913 => x"ef",
          3914 => x"c3",
          3915 => x"e8",
          3916 => x"16",
          3917 => x"58",
          3918 => x"3f",
          3919 => x"0a",
          3920 => x"0a",
          3921 => x"2c",
          3922 => x"33",
          3923 => x"76",
          3924 => x"38",
          3925 => x"33",
          3926 => x"70",
          3927 => x"81",
          3928 => x"58",
          3929 => x"79",
          3930 => x"38",
          3931 => x"83",
          3932 => x"80",
          3933 => x"38",
          3934 => x"57",
          3935 => x"08",
          3936 => x"38",
          3937 => x"18",
          3938 => x"80",
          3939 => x"80",
          3940 => x"f4",
          3941 => x"ec",
          3942 => x"80",
          3943 => x"38",
          3944 => x"e7",
          3945 => x"f4",
          3946 => x"80",
          3947 => x"80",
          3948 => x"ec",
          3949 => x"b5",
          3950 => x"ee",
          3951 => x"51",
          3952 => x"3f",
          3953 => x"ff",
          3954 => x"58",
          3955 => x"25",
          3956 => x"ff",
          3957 => x"51",
          3958 => x"3f",
          3959 => x"08",
          3960 => x"34",
          3961 => x"08",
          3962 => x"81",
          3963 => x"52",
          3964 => x"aa",
          3965 => x"0b",
          3966 => x"33",
          3967 => x"33",
          3968 => x"74",
          3969 => x"c4",
          3970 => x"e8",
          3971 => x"51",
          3972 => x"3f",
          3973 => x"08",
          3974 => x"ff",
          3975 => x"84",
          3976 => x"52",
          3977 => x"a6",
          3978 => x"e2",
          3979 => x"05",
          3980 => x"e2",
          3981 => x"81",
          3982 => x"c7",
          3983 => x"ff",
          3984 => x"84",
          3985 => x"84",
          3986 => x"84",
          3987 => x"81",
          3988 => x"05",
          3989 => x"7b",
          3990 => x"8f",
          3991 => x"e2",
          3992 => x"e2",
          3993 => x"57",
          3994 => x"2e",
          3995 => x"84",
          3996 => x"52",
          3997 => x"a5",
          3998 => x"e6",
          3999 => x"a0",
          4000 => x"eb",
          4001 => x"e8",
          4002 => x"51",
          4003 => x"3f",
          4004 => x"33",
          4005 => x"76",
          4006 => x"34",
          4007 => x"06",
          4008 => x"75",
          4009 => x"81",
          4010 => x"84",
          4011 => x"c4",
          4012 => x"84",
          4013 => x"06",
          4014 => x"75",
          4015 => x"ff",
          4016 => x"81",
          4017 => x"ff",
          4018 => x"c4",
          4019 => x"c8",
          4020 => x"5e",
          4021 => x"2e",
          4022 => x"84",
          4023 => x"52",
          4024 => x"a5",
          4025 => x"e6",
          4026 => x"a0",
          4027 => x"ff",
          4028 => x"e8",
          4029 => x"51",
          4030 => x"3f",
          4031 => x"33",
          4032 => x"7a",
          4033 => x"34",
          4034 => x"06",
          4035 => x"80",
          4036 => x"0b",
          4037 => x"34",
          4038 => x"e2",
          4039 => x"84",
          4040 => x"b5",
          4041 => x"83",
          4042 => x"56",
          4043 => x"ef",
          4044 => x"51",
          4045 => x"3f",
          4046 => x"08",
          4047 => x"34",
          4048 => x"08",
          4049 => x"81",
          4050 => x"52",
          4051 => x"a8",
          4052 => x"e2",
          4053 => x"e2",
          4054 => x"56",
          4055 => x"ef",
          4056 => x"e6",
          4057 => x"88",
          4058 => x"83",
          4059 => x"e8",
          4060 => x"51",
          4061 => x"3f",
          4062 => x"08",
          4063 => x"ff",
          4064 => x"84",
          4065 => x"ff",
          4066 => x"84",
          4067 => x"78",
          4068 => x"55",
          4069 => x"51",
          4070 => x"3f",
          4071 => x"33",
          4072 => x"87",
          4073 => x"f4",
          4074 => x"19",
          4075 => x"5a",
          4076 => x"96",
          4077 => x"84",
          4078 => x"83",
          4079 => x"70",
          4080 => x"f4",
          4081 => x"08",
          4082 => x"e3",
          4083 => x"ff",
          4084 => x"83",
          4085 => x"70",
          4086 => x"f4",
          4087 => x"08",
          4088 => x"74",
          4089 => x"b3",
          4090 => x"7b",
          4091 => x"ff",
          4092 => x"83",
          4093 => x"81",
          4094 => x"ff",
          4095 => x"93",
          4096 => x"9f",
          4097 => x"f4",
          4098 => x"8f",
          4099 => x"fe",
          4100 => x"76",
          4101 => x"75",
          4102 => x"8a",
          4103 => x"ec",
          4104 => x"51",
          4105 => x"3f",
          4106 => x"08",
          4107 => x"89",
          4108 => x"84",
          4109 => x"80",
          4110 => x"c4",
          4111 => x"bb",
          4112 => x"3d",
          4113 => x"53",
          4114 => x"51",
          4115 => x"3f",
          4116 => x"08",
          4117 => x"84",
          4118 => x"97",
          4119 => x"83",
          4120 => x"53",
          4121 => x"7a",
          4122 => x"e9",
          4123 => x"84",
          4124 => x"bb",
          4125 => x"2e",
          4126 => x"e8",
          4127 => x"bb",
          4128 => x"ff",
          4129 => x"84",
          4130 => x"57",
          4131 => x"bb",
          4132 => x"80",
          4133 => x"bb",
          4134 => x"05",
          4135 => x"57",
          4136 => x"76",
          4137 => x"83",
          4138 => x"70",
          4139 => x"f4",
          4140 => x"08",
          4141 => x"59",
          4142 => x"38",
          4143 => x"87",
          4144 => x"f4",
          4145 => x"1a",
          4146 => x"5f",
          4147 => x"3f",
          4148 => x"08",
          4149 => x"f4",
          4150 => x"10",
          4151 => x"9c",
          4152 => x"54",
          4153 => x"94",
          4154 => x"92",
          4155 => x"f4",
          4156 => x"10",
          4157 => x"9c",
          4158 => x"57",
          4159 => x"a0",
          4160 => x"70",
          4161 => x"5e",
          4162 => x"27",
          4163 => x"5d",
          4164 => x"09",
          4165 => x"c7",
          4166 => x"dc",
          4167 => x"39",
          4168 => x"52",
          4169 => x"a4",
          4170 => x"f4",
          4171 => x"05",
          4172 => x"06",
          4173 => x"7a",
          4174 => x"38",
          4175 => x"f4",
          4176 => x"bd",
          4177 => x"80",
          4178 => x"83",
          4179 => x"70",
          4180 => x"fc",
          4181 => x"9c",
          4182 => x"70",
          4183 => x"56",
          4184 => x"3f",
          4185 => x"08",
          4186 => x"f4",
          4187 => x"10",
          4188 => x"9c",
          4189 => x"54",
          4190 => x"94",
          4191 => x"91",
          4192 => x"f4",
          4193 => x"10",
          4194 => x"9c",
          4195 => x"57",
          4196 => x"80",
          4197 => x"38",
          4198 => x"75",
          4199 => x"34",
          4200 => x"75",
          4201 => x"34",
          4202 => x"83",
          4203 => x"ff",
          4204 => x"77",
          4205 => x"f7",
          4206 => x"3d",
          4207 => x"c3",
          4208 => x"84",
          4209 => x"05",
          4210 => x"72",
          4211 => x"8d",
          4212 => x"2e",
          4213 => x"81",
          4214 => x"9e",
          4215 => x"2e",
          4216 => x"86",
          4217 => x"59",
          4218 => x"80",
          4219 => x"80",
          4220 => x"58",
          4221 => x"90",
          4222 => x"fa",
          4223 => x"83",
          4224 => x"75",
          4225 => x"23",
          4226 => x"33",
          4227 => x"71",
          4228 => x"71",
          4229 => x"71",
          4230 => x"56",
          4231 => x"78",
          4232 => x"38",
          4233 => x"84",
          4234 => x"74",
          4235 => x"05",
          4236 => x"74",
          4237 => x"75",
          4238 => x"38",
          4239 => x"33",
          4240 => x"17",
          4241 => x"55",
          4242 => x"0b",
          4243 => x"34",
          4244 => x"81",
          4245 => x"ff",
          4246 => x"ee",
          4247 => x"0d",
          4248 => x"a0",
          4249 => x"fa",
          4250 => x"10",
          4251 => x"fa",
          4252 => x"90",
          4253 => x"05",
          4254 => x"40",
          4255 => x"b0",
          4256 => x"b8",
          4257 => x"81",
          4258 => x"b8",
          4259 => x"81",
          4260 => x"fa",
          4261 => x"83",
          4262 => x"70",
          4263 => x"59",
          4264 => x"57",
          4265 => x"73",
          4266 => x"72",
          4267 => x"29",
          4268 => x"ff",
          4269 => x"ff",
          4270 => x"ff",
          4271 => x"ff",
          4272 => x"81",
          4273 => x"75",
          4274 => x"42",
          4275 => x"5c",
          4276 => x"8f",
          4277 => x"b4",
          4278 => x"31",
          4279 => x"29",
          4280 => x"76",
          4281 => x"7b",
          4282 => x"9c",
          4283 => x"55",
          4284 => x"26",
          4285 => x"80",
          4286 => x"05",
          4287 => x"fa",
          4288 => x"70",
          4289 => x"34",
          4290 => x"c7",
          4291 => x"86",
          4292 => x"70",
          4293 => x"33",
          4294 => x"06",
          4295 => x"33",
          4296 => x"06",
          4297 => x"22",
          4298 => x"5d",
          4299 => x"5e",
          4300 => x"74",
          4301 => x"df",
          4302 => x"ff",
          4303 => x"ff",
          4304 => x"29",
          4305 => x"54",
          4306 => x"fd",
          4307 => x"0b",
          4308 => x"34",
          4309 => x"fa",
          4310 => x"fa",
          4311 => x"98",
          4312 => x"2b",
          4313 => x"2b",
          4314 => x"7a",
          4315 => x"56",
          4316 => x"26",
          4317 => x"fd",
          4318 => x"fc",
          4319 => x"fa",
          4320 => x"81",
          4321 => x"10",
          4322 => x"fa",
          4323 => x"90",
          4324 => x"c7",
          4325 => x"5e",
          4326 => x"56",
          4327 => x"b0",
          4328 => x"84",
          4329 => x"70",
          4330 => x"84",
          4331 => x"70",
          4332 => x"83",
          4333 => x"70",
          4334 => x"06",
          4335 => x"60",
          4336 => x"41",
          4337 => x"40",
          4338 => x"73",
          4339 => x"72",
          4340 => x"70",
          4341 => x"57",
          4342 => x"ff",
          4343 => x"ff",
          4344 => x"29",
          4345 => x"ff",
          4346 => x"ff",
          4347 => x"29",
          4348 => x"5c",
          4349 => x"78",
          4350 => x"77",
          4351 => x"79",
          4352 => x"79",
          4353 => x"58",
          4354 => x"38",
          4355 => x"5c",
          4356 => x"38",
          4357 => x"74",
          4358 => x"29",
          4359 => x"39",
          4360 => x"87",
          4361 => x"53",
          4362 => x"34",
          4363 => x"85",
          4364 => x"73",
          4365 => x"80",
          4366 => x"f4",
          4367 => x"b0",
          4368 => x"8e",
          4369 => x"80",
          4370 => x"76",
          4371 => x"80",
          4372 => x"74",
          4373 => x"34",
          4374 => x"34",
          4375 => x"51",
          4376 => x"86",
          4377 => x"70",
          4378 => x"81",
          4379 => x"c0",
          4380 => x"77",
          4381 => x"54",
          4382 => x"34",
          4383 => x"80",
          4384 => x"c0",
          4385 => x"72",
          4386 => x"c0",
          4387 => x"70",
          4388 => x"07",
          4389 => x"86",
          4390 => x"34",
          4391 => x"f7",
          4392 => x"53",
          4393 => x"80",
          4394 => x"b8",
          4395 => x"0b",
          4396 => x"0c",
          4397 => x"04",
          4398 => x"33",
          4399 => x"0c",
          4400 => x"0d",
          4401 => x"33",
          4402 => x"b3",
          4403 => x"b8",
          4404 => x"59",
          4405 => x"75",
          4406 => x"da",
          4407 => x"f8",
          4408 => x"b5",
          4409 => x"b4",
          4410 => x"29",
          4411 => x"a0",
          4412 => x"fa",
          4413 => x"51",
          4414 => x"7c",
          4415 => x"83",
          4416 => x"83",
          4417 => x"53",
          4418 => x"72",
          4419 => x"c4",
          4420 => x"b2",
          4421 => x"55",
          4422 => x"b2",
          4423 => x"b4",
          4424 => x"70",
          4425 => x"7a",
          4426 => x"55",
          4427 => x"7a",
          4428 => x"38",
          4429 => x"72",
          4430 => x"34",
          4431 => x"22",
          4432 => x"ff",
          4433 => x"f6",
          4434 => x"57",
          4435 => x"82",
          4436 => x"b8",
          4437 => x"71",
          4438 => x"80",
          4439 => x"9f",
          4440 => x"84",
          4441 => x"14",
          4442 => x"e0",
          4443 => x"e0",
          4444 => x"70",
          4445 => x"33",
          4446 => x"05",
          4447 => x"14",
          4448 => x"f5",
          4449 => x"38",
          4450 => x"26",
          4451 => x"fa",
          4452 => x"99",
          4453 => x"55",
          4454 => x"e0",
          4455 => x"73",
          4456 => x"55",
          4457 => x"54",
          4458 => x"27",
          4459 => x"b8",
          4460 => x"05",
          4461 => x"fa",
          4462 => x"57",
          4463 => x"06",
          4464 => x"ff",
          4465 => x"73",
          4466 => x"fd",
          4467 => x"31",
          4468 => x"b8",
          4469 => x"71",
          4470 => x"57",
          4471 => x"c7",
          4472 => x"86",
          4473 => x"79",
          4474 => x"75",
          4475 => x"71",
          4476 => x"5c",
          4477 => x"75",
          4478 => x"38",
          4479 => x"16",
          4480 => x"14",
          4481 => x"b9",
          4482 => x"78",
          4483 => x"5a",
          4484 => x"81",
          4485 => x"77",
          4486 => x"59",
          4487 => x"84",
          4488 => x"84",
          4489 => x"71",
          4490 => x"56",
          4491 => x"72",
          4492 => x"38",
          4493 => x"84",
          4494 => x"8b",
          4495 => x"74",
          4496 => x"34",
          4497 => x"22",
          4498 => x"ff",
          4499 => x"f6",
          4500 => x"57",
          4501 => x"fd",
          4502 => x"80",
          4503 => x"38",
          4504 => x"06",
          4505 => x"fa",
          4506 => x"53",
          4507 => x"09",
          4508 => x"c8",
          4509 => x"31",
          4510 => x"b8",
          4511 => x"71",
          4512 => x"29",
          4513 => x"59",
          4514 => x"27",
          4515 => x"83",
          4516 => x"84",
          4517 => x"74",
          4518 => x"56",
          4519 => x"e0",
          4520 => x"75",
          4521 => x"05",
          4522 => x"13",
          4523 => x"2e",
          4524 => x"a0",
          4525 => x"16",
          4526 => x"70",
          4527 => x"34",
          4528 => x"72",
          4529 => x"f4",
          4530 => x"84",
          4531 => x"55",
          4532 => x"39",
          4533 => x"15",
          4534 => x"b9",
          4535 => x"74",
          4536 => x"f7",
          4537 => x"a9",
          4538 => x"0d",
          4539 => x"05",
          4540 => x"53",
          4541 => x"26",
          4542 => x"10",
          4543 => x"fc",
          4544 => x"08",
          4545 => x"f8",
          4546 => x"71",
          4547 => x"71",
          4548 => x"34",
          4549 => x"bb",
          4550 => x"3d",
          4551 => x"0b",
          4552 => x"34",
          4553 => x"33",
          4554 => x"06",
          4555 => x"80",
          4556 => x"ff",
          4557 => x"83",
          4558 => x"80",
          4559 => x"84",
          4560 => x"0d",
          4561 => x"b4",
          4562 => x"31",
          4563 => x"9f",
          4564 => x"54",
          4565 => x"70",
          4566 => x"34",
          4567 => x"fa",
          4568 => x"05",
          4569 => x"33",
          4570 => x"56",
          4571 => x"25",
          4572 => x"53",
          4573 => x"b4",
          4574 => x"84",
          4575 => x"86",
          4576 => x"83",
          4577 => x"70",
          4578 => x"09",
          4579 => x"72",
          4580 => x"53",
          4581 => x"fa",
          4582 => x"0b",
          4583 => x"0c",
          4584 => x"04",
          4585 => x"33",
          4586 => x"b8",
          4587 => x"11",
          4588 => x"70",
          4589 => x"38",
          4590 => x"83",
          4591 => x"80",
          4592 => x"84",
          4593 => x"0d",
          4594 => x"83",
          4595 => x"83",
          4596 => x"84",
          4597 => x"ff",
          4598 => x"71",
          4599 => x"b4",
          4600 => x"51",
          4601 => x"b4",
          4602 => x"39",
          4603 => x"02",
          4604 => x"51",
          4605 => x"b3",
          4606 => x"10",
          4607 => x"05",
          4608 => x"04",
          4609 => x"33",
          4610 => x"06",
          4611 => x"80",
          4612 => x"72",
          4613 => x"51",
          4614 => x"71",
          4615 => x"09",
          4616 => x"38",
          4617 => x"83",
          4618 => x"80",
          4619 => x"84",
          4620 => x"0d",
          4621 => x"b0",
          4622 => x"06",
          4623 => x"70",
          4624 => x"34",
          4625 => x"bb",
          4626 => x"3d",
          4627 => x"fa",
          4628 => x"f0",
          4629 => x"83",
          4630 => x"e8",
          4631 => x"b0",
          4632 => x"06",
          4633 => x"70",
          4634 => x"34",
          4635 => x"f1",
          4636 => x"b0",
          4637 => x"84",
          4638 => x"83",
          4639 => x"83",
          4640 => x"81",
          4641 => x"07",
          4642 => x"fa",
          4643 => x"b4",
          4644 => x"b0",
          4645 => x"51",
          4646 => x"b0",
          4647 => x"39",
          4648 => x"33",
          4649 => x"85",
          4650 => x"83",
          4651 => x"ff",
          4652 => x"fa",
          4653 => x"fb",
          4654 => x"51",
          4655 => x"b0",
          4656 => x"39",
          4657 => x"33",
          4658 => x"81",
          4659 => x"83",
          4660 => x"fe",
          4661 => x"fa",
          4662 => x"f8",
          4663 => x"83",
          4664 => x"fe",
          4665 => x"fa",
          4666 => x"df",
          4667 => x"07",
          4668 => x"fa",
          4669 => x"cc",
          4670 => x"b0",
          4671 => x"06",
          4672 => x"70",
          4673 => x"34",
          4674 => x"83",
          4675 => x"81",
          4676 => x"e0",
          4677 => x"83",
          4678 => x"fe",
          4679 => x"fa",
          4680 => x"cf",
          4681 => x"07",
          4682 => x"fa",
          4683 => x"94",
          4684 => x"b0",
          4685 => x"06",
          4686 => x"70",
          4687 => x"34",
          4688 => x"83",
          4689 => x"81",
          4690 => x"70",
          4691 => x"34",
          4692 => x"83",
          4693 => x"81",
          4694 => x"07",
          4695 => x"fa",
          4696 => x"e0",
          4697 => x"0d",
          4698 => x"33",
          4699 => x"80",
          4700 => x"83",
          4701 => x"83",
          4702 => x"83",
          4703 => x"84",
          4704 => x"43",
          4705 => x"5b",
          4706 => x"2e",
          4707 => x"78",
          4708 => x"38",
          4709 => x"81",
          4710 => x"84",
          4711 => x"80",
          4712 => x"fc",
          4713 => x"fa",
          4714 => x"83",
          4715 => x"7c",
          4716 => x"34",
          4717 => x"04",
          4718 => x"09",
          4719 => x"38",
          4720 => x"b8",
          4721 => x"0b",
          4722 => x"34",
          4723 => x"fa",
          4724 => x"0b",
          4725 => x"34",
          4726 => x"fa",
          4727 => x"58",
          4728 => x"33",
          4729 => x"f7",
          4730 => x"b8",
          4731 => x"7b",
          4732 => x"7a",
          4733 => x"f8",
          4734 => x"8d",
          4735 => x"b8",
          4736 => x"0b",
          4737 => x"34",
          4738 => x"b4",
          4739 => x"fa",
          4740 => x"83",
          4741 => x"8f",
          4742 => x"80",
          4743 => x"fa",
          4744 => x"84",
          4745 => x"80",
          4746 => x"b4",
          4747 => x"83",
          4748 => x"80",
          4749 => x"b2",
          4750 => x"87",
          4751 => x"ba",
          4752 => x"84",
          4753 => x"56",
          4754 => x"54",
          4755 => x"52",
          4756 => x"51",
          4757 => x"3f",
          4758 => x"ba",
          4759 => x"5a",
          4760 => x"a5",
          4761 => x"84",
          4762 => x"70",
          4763 => x"83",
          4764 => x"fe",
          4765 => x"81",
          4766 => x"ff",
          4767 => x"85",
          4768 => x"59",
          4769 => x"dd",
          4770 => x"b4",
          4771 => x"f9",
          4772 => x"b8",
          4773 => x"0b",
          4774 => x"34",
          4775 => x"b4",
          4776 => x"fa",
          4777 => x"83",
          4778 => x"8f",
          4779 => x"80",
          4780 => x"fa",
          4781 => x"84",
          4782 => x"81",
          4783 => x"b4",
          4784 => x"83",
          4785 => x"81",
          4786 => x"b2",
          4787 => x"e8",
          4788 => x"d5",
          4789 => x"84",
          4790 => x"e5",
          4791 => x"fe",
          4792 => x"59",
          4793 => x"51",
          4794 => x"3f",
          4795 => x"84",
          4796 => x"a6",
          4797 => x"e8",
          4798 => x"83",
          4799 => x"fe",
          4800 => x"81",
          4801 => x"ff",
          4802 => x"d8",
          4803 => x"0d",
          4804 => x"05",
          4805 => x"84",
          4806 => x"83",
          4807 => x"83",
          4808 => x"72",
          4809 => x"86",
          4810 => x"11",
          4811 => x"22",
          4812 => x"5c",
          4813 => x"05",
          4814 => x"ff",
          4815 => x"8a",
          4816 => x"51",
          4817 => x"72",
          4818 => x"e9",
          4819 => x"2e",
          4820 => x"75",
          4821 => x"b9",
          4822 => x"2e",
          4823 => x"75",
          4824 => x"d5",
          4825 => x"f8",
          4826 => x"b4",
          4827 => x"b5",
          4828 => x"29",
          4829 => x"54",
          4830 => x"16",
          4831 => x"a0",
          4832 => x"84",
          4833 => x"83",
          4834 => x"83",
          4835 => x"72",
          4836 => x"5a",
          4837 => x"75",
          4838 => x"18",
          4839 => x"b4",
          4840 => x"29",
          4841 => x"83",
          4842 => x"86",
          4843 => x"18",
          4844 => x"f8",
          4845 => x"ff",
          4846 => x"b2",
          4847 => x"b5",
          4848 => x"29",
          4849 => x"57",
          4850 => x"fa",
          4851 => x"99",
          4852 => x"81",
          4853 => x"ff",
          4854 => x"73",
          4855 => x"99",
          4856 => x"f9",
          4857 => x"81",
          4858 => x"17",
          4859 => x"fa",
          4860 => x"b8",
          4861 => x"72",
          4862 => x"38",
          4863 => x"33",
          4864 => x"2e",
          4865 => x"80",
          4866 => x"84",
          4867 => x"0d",
          4868 => x"2e",
          4869 => x"8d",
          4870 => x"38",
          4871 => x"09",
          4872 => x"c1",
          4873 => x"81",
          4874 => x"3f",
          4875 => x"fa",
          4876 => x"be",
          4877 => x"b6",
          4878 => x"84",
          4879 => x"33",
          4880 => x"89",
          4881 => x"06",
          4882 => x"80",
          4883 => x"a0",
          4884 => x"3f",
          4885 => x"81",
          4886 => x"54",
          4887 => x"ff",
          4888 => x"52",
          4889 => x"a5",
          4890 => x"70",
          4891 => x"54",
          4892 => x"27",
          4893 => x"fa",
          4894 => x"fa",
          4895 => x"f2",
          4896 => x"83",
          4897 => x"3f",
          4898 => x"bb",
          4899 => x"3d",
          4900 => x"80",
          4901 => x"81",
          4902 => x"38",
          4903 => x"33",
          4904 => x"06",
          4905 => x"53",
          4906 => x"73",
          4907 => x"fa",
          4908 => x"52",
          4909 => x"d5",
          4910 => x"b5",
          4911 => x"ff",
          4912 => x"05",
          4913 => x"a5",
          4914 => x"72",
          4915 => x"34",
          4916 => x"80",
          4917 => x"b5",
          4918 => x"81",
          4919 => x"3f",
          4920 => x"80",
          4921 => x"ef",
          4922 => x"86",
          4923 => x"0d",
          4924 => x"05",
          4925 => x"80",
          4926 => x"75",
          4927 => x"b8",
          4928 => x"2e",
          4929 => x"78",
          4930 => x"b5",
          4931 => x"24",
          4932 => x"78",
          4933 => x"b9",
          4934 => x"2e",
          4935 => x"84",
          4936 => x"83",
          4937 => x"83",
          4938 => x"72",
          4939 => x"58",
          4940 => x"b9",
          4941 => x"86",
          4942 => x"17",
          4943 => x"f8",
          4944 => x"b5",
          4945 => x"b2",
          4946 => x"29",
          4947 => x"42",
          4948 => x"fa",
          4949 => x"83",
          4950 => x"60",
          4951 => x"05",
          4952 => x"fa",
          4953 => x"86",
          4954 => x"05",
          4955 => x"f8",
          4956 => x"ff",
          4957 => x"b2",
          4958 => x"b5",
          4959 => x"29",
          4960 => x"5d",
          4961 => x"fa",
          4962 => x"99",
          4963 => x"81",
          4964 => x"ff",
          4965 => x"76",
          4966 => x"b8",
          4967 => x"f9",
          4968 => x"86",
          4969 => x"19",
          4970 => x"fa",
          4971 => x"0b",
          4972 => x"0c",
          4973 => x"04",
          4974 => x"84",
          4975 => x"79",
          4976 => x"38",
          4977 => x"9b",
          4978 => x"80",
          4979 => x"cc",
          4980 => x"84",
          4981 => x"84",
          4982 => x"83",
          4983 => x"83",
          4984 => x"72",
          4985 => x"5e",
          4986 => x"b9",
          4987 => x"86",
          4988 => x"1d",
          4989 => x"f8",
          4990 => x"b5",
          4991 => x"b2",
          4992 => x"29",
          4993 => x"59",
          4994 => x"fa",
          4995 => x"83",
          4996 => x"76",
          4997 => x"5b",
          4998 => x"b0",
          4999 => x"b0",
          5000 => x"84",
          5001 => x"70",
          5002 => x"83",
          5003 => x"83",
          5004 => x"72",
          5005 => x"44",
          5006 => x"59",
          5007 => x"33",
          5008 => x"d6",
          5009 => x"1f",
          5010 => x"ff",
          5011 => x"77",
          5012 => x"38",
          5013 => x"b5",
          5014 => x"84",
          5015 => x"9c",
          5016 => x"78",
          5017 => x"b7",
          5018 => x"24",
          5019 => x"78",
          5020 => x"81",
          5021 => x"38",
          5022 => x"fa",
          5023 => x"0b",
          5024 => x"0c",
          5025 => x"04",
          5026 => x"82",
          5027 => x"19",
          5028 => x"26",
          5029 => x"84",
          5030 => x"81",
          5031 => x"77",
          5032 => x"34",
          5033 => x"88",
          5034 => x"81",
          5035 => x"80",
          5036 => x"88",
          5037 => x"0b",
          5038 => x"0c",
          5039 => x"04",
          5040 => x"fd",
          5041 => x"0b",
          5042 => x"0c",
          5043 => x"33",
          5044 => x"33",
          5045 => x"33",
          5046 => x"05",
          5047 => x"84",
          5048 => x"33",
          5049 => x"80",
          5050 => x"b8",
          5051 => x"fa",
          5052 => x"fa",
          5053 => x"71",
          5054 => x"5f",
          5055 => x"83",
          5056 => x"34",
          5057 => x"33",
          5058 => x"19",
          5059 => x"fa",
          5060 => x"c7",
          5061 => x"34",
          5062 => x"33",
          5063 => x"06",
          5064 => x"22",
          5065 => x"33",
          5066 => x"11",
          5067 => x"58",
          5068 => x"b0",
          5069 => x"99",
          5070 => x"81",
          5071 => x"89",
          5072 => x"81",
          5073 => x"3f",
          5074 => x"fa",
          5075 => x"ae",
          5076 => x"f8",
          5077 => x"b5",
          5078 => x"ff",
          5079 => x"b4",
          5080 => x"29",
          5081 => x"a0",
          5082 => x"fa",
          5083 => x"51",
          5084 => x"29",
          5085 => x"ff",
          5086 => x"f9",
          5087 => x"51",
          5088 => x"75",
          5089 => x"a4",
          5090 => x"ff",
          5091 => x"57",
          5092 => x"95",
          5093 => x"75",
          5094 => x"34",
          5095 => x"80",
          5096 => x"84",
          5097 => x"84",
          5098 => x"80",
          5099 => x"86",
          5100 => x"84",
          5101 => x"81",
          5102 => x"80",
          5103 => x"84",
          5104 => x"9c",
          5105 => x"83",
          5106 => x"84",
          5107 => x"83",
          5108 => x"84",
          5109 => x"83",
          5110 => x"84",
          5111 => x"80",
          5112 => x"80",
          5113 => x"84",
          5114 => x"9c",
          5115 => x"78",
          5116 => x"09",
          5117 => x"a7",
          5118 => x"b4",
          5119 => x"f8",
          5120 => x"ff",
          5121 => x"b5",
          5122 => x"ff",
          5123 => x"29",
          5124 => x"a0",
          5125 => x"fa",
          5126 => x"40",
          5127 => x"05",
          5128 => x"ff",
          5129 => x"8a",
          5130 => x"43",
          5131 => x"5c",
          5132 => x"85",
          5133 => x"81",
          5134 => x"1a",
          5135 => x"83",
          5136 => x"76",
          5137 => x"34",
          5138 => x"06",
          5139 => x"06",
          5140 => x"06",
          5141 => x"05",
          5142 => x"84",
          5143 => x"86",
          5144 => x"1e",
          5145 => x"f8",
          5146 => x"b5",
          5147 => x"b2",
          5148 => x"29",
          5149 => x"42",
          5150 => x"83",
          5151 => x"34",
          5152 => x"33",
          5153 => x"62",
          5154 => x"83",
          5155 => x"86",
          5156 => x"1a",
          5157 => x"f8",
          5158 => x"ff",
          5159 => x"b2",
          5160 => x"b5",
          5161 => x"29",
          5162 => x"5a",
          5163 => x"fa",
          5164 => x"84",
          5165 => x"34",
          5166 => x"81",
          5167 => x"58",
          5168 => x"95",
          5169 => x"b8",
          5170 => x"79",
          5171 => x"ff",
          5172 => x"83",
          5173 => x"83",
          5174 => x"70",
          5175 => x"58",
          5176 => x"fd",
          5177 => x"bb",
          5178 => x"38",
          5179 => x"83",
          5180 => x"bf",
          5181 => x"38",
          5182 => x"33",
          5183 => x"f9",
          5184 => x"19",
          5185 => x"26",
          5186 => x"75",
          5187 => x"c6",
          5188 => x"77",
          5189 => x"0b",
          5190 => x"34",
          5191 => x"51",
          5192 => x"80",
          5193 => x"84",
          5194 => x"0d",
          5195 => x"b4",
          5196 => x"f8",
          5197 => x"ff",
          5198 => x"b5",
          5199 => x"ff",
          5200 => x"29",
          5201 => x"a0",
          5202 => x"fa",
          5203 => x"41",
          5204 => x"05",
          5205 => x"ff",
          5206 => x"8a",
          5207 => x"45",
          5208 => x"5b",
          5209 => x"82",
          5210 => x"5c",
          5211 => x"06",
          5212 => x"06",
          5213 => x"06",
          5214 => x"05",
          5215 => x"84",
          5216 => x"86",
          5217 => x"1b",
          5218 => x"f8",
          5219 => x"b5",
          5220 => x"b2",
          5221 => x"29",
          5222 => x"5e",
          5223 => x"83",
          5224 => x"34",
          5225 => x"33",
          5226 => x"1e",
          5227 => x"fa",
          5228 => x"c7",
          5229 => x"34",
          5230 => x"33",
          5231 => x"06",
          5232 => x"22",
          5233 => x"33",
          5234 => x"11",
          5235 => x"40",
          5236 => x"b0",
          5237 => x"d6",
          5238 => x"81",
          5239 => x"ff",
          5240 => x"7e",
          5241 => x"ac",
          5242 => x"f9",
          5243 => x"92",
          5244 => x"19",
          5245 => x"fa",
          5246 => x"1c",
          5247 => x"06",
          5248 => x"83",
          5249 => x"38",
          5250 => x"33",
          5251 => x"33",
          5252 => x"33",
          5253 => x"06",
          5254 => x"06",
          5255 => x"06",
          5256 => x"05",
          5257 => x"5b",
          5258 => x"b9",
          5259 => x"c7",
          5260 => x"34",
          5261 => x"33",
          5262 => x"33",
          5263 => x"22",
          5264 => x"12",
          5265 => x"56",
          5266 => x"fa",
          5267 => x"83",
          5268 => x"76",
          5269 => x"5a",
          5270 => x"b0",
          5271 => x"b0",
          5272 => x"84",
          5273 => x"70",
          5274 => x"83",
          5275 => x"83",
          5276 => x"72",
          5277 => x"5b",
          5278 => x"59",
          5279 => x"33",
          5280 => x"18",
          5281 => x"05",
          5282 => x"06",
          5283 => x"7f",
          5284 => x"38",
          5285 => x"b5",
          5286 => x"39",
          5287 => x"ba",
          5288 => x"0b",
          5289 => x"0c",
          5290 => x"04",
          5291 => x"17",
          5292 => x"b9",
          5293 => x"7a",
          5294 => x"b5",
          5295 => x"ff",
          5296 => x"05",
          5297 => x"39",
          5298 => x"ba",
          5299 => x"0b",
          5300 => x"0c",
          5301 => x"04",
          5302 => x"17",
          5303 => x"b9",
          5304 => x"7c",
          5305 => x"b4",
          5306 => x"f8",
          5307 => x"b5",
          5308 => x"5b",
          5309 => x"f4",
          5310 => x"88",
          5311 => x"dc",
          5312 => x"05",
          5313 => x"ff",
          5314 => x"84",
          5315 => x"fb",
          5316 => x"ba",
          5317 => x"11",
          5318 => x"84",
          5319 => x"79",
          5320 => x"06",
          5321 => x"ca",
          5322 => x"84",
          5323 => x"23",
          5324 => x"83",
          5325 => x"33",
          5326 => x"80",
          5327 => x"34",
          5328 => x"33",
          5329 => x"33",
          5330 => x"33",
          5331 => x"f9",
          5332 => x"b8",
          5333 => x"fa",
          5334 => x"fa",
          5335 => x"72",
          5336 => x"5d",
          5337 => x"80",
          5338 => x"86",
          5339 => x"05",
          5340 => x"f8",
          5341 => x"b5",
          5342 => x"b2",
          5343 => x"29",
          5344 => x"5b",
          5345 => x"fa",
          5346 => x"83",
          5347 => x"76",
          5348 => x"41",
          5349 => x"b0",
          5350 => x"c7",
          5351 => x"34",
          5352 => x"33",
          5353 => x"06",
          5354 => x"22",
          5355 => x"33",
          5356 => x"11",
          5357 => x"42",
          5358 => x"b0",
          5359 => x"d6",
          5360 => x"1c",
          5361 => x"06",
          5362 => x"7b",
          5363 => x"38",
          5364 => x"33",
          5365 => x"e2",
          5366 => x"56",
          5367 => x"b5",
          5368 => x"84",
          5369 => x"84",
          5370 => x"40",
          5371 => x"f3",
          5372 => x"b8",
          5373 => x"75",
          5374 => x"78",
          5375 => x"ea",
          5376 => x"0b",
          5377 => x"0c",
          5378 => x"04",
          5379 => x"33",
          5380 => x"34",
          5381 => x"33",
          5382 => x"34",
          5383 => x"33",
          5384 => x"fa",
          5385 => x"b9",
          5386 => x"b4",
          5387 => x"ec",
          5388 => x"b5",
          5389 => x"ed",
          5390 => x"b3",
          5391 => x"ee",
          5392 => x"39",
          5393 => x"33",
          5394 => x"2e",
          5395 => x"84",
          5396 => x"5d",
          5397 => x"09",
          5398 => x"85",
          5399 => x"b5",
          5400 => x"55",
          5401 => x"33",
          5402 => x"9b",
          5403 => x"c0",
          5404 => x"70",
          5405 => x"ec",
          5406 => x"51",
          5407 => x"3f",
          5408 => x"08",
          5409 => x"83",
          5410 => x"57",
          5411 => x"60",
          5412 => x"cd",
          5413 => x"83",
          5414 => x"fe",
          5415 => x"fe",
          5416 => x"0b",
          5417 => x"33",
          5418 => x"81",
          5419 => x"77",
          5420 => x"ad",
          5421 => x"84",
          5422 => x"81",
          5423 => x"41",
          5424 => x"8a",
          5425 => x"10",
          5426 => x"b4",
          5427 => x"08",
          5428 => x"85",
          5429 => x"80",
          5430 => x"38",
          5431 => x"33",
          5432 => x"33",
          5433 => x"70",
          5434 => x"2c",
          5435 => x"42",
          5436 => x"75",
          5437 => x"34",
          5438 => x"84",
          5439 => x"56",
          5440 => x"8e",
          5441 => x"ba",
          5442 => x"05",
          5443 => x"06",
          5444 => x"33",
          5445 => x"75",
          5446 => x"c5",
          5447 => x"fa",
          5448 => x"bd",
          5449 => x"83",
          5450 => x"83",
          5451 => x"70",
          5452 => x"5d",
          5453 => x"2e",
          5454 => x"ff",
          5455 => x"83",
          5456 => x"fd",
          5457 => x"0b",
          5458 => x"34",
          5459 => x"33",
          5460 => x"33",
          5461 => x"57",
          5462 => x"fd",
          5463 => x"17",
          5464 => x"fa",
          5465 => x"f9",
          5466 => x"85",
          5467 => x"80",
          5468 => x"38",
          5469 => x"33",
          5470 => x"33",
          5471 => x"70",
          5472 => x"2c",
          5473 => x"41",
          5474 => x"75",
          5475 => x"34",
          5476 => x"84",
          5477 => x"5b",
          5478 => x"fc",
          5479 => x"ba",
          5480 => x"60",
          5481 => x"81",
          5482 => x"38",
          5483 => x"33",
          5484 => x"33",
          5485 => x"33",
          5486 => x"12",
          5487 => x"80",
          5488 => x"b2",
          5489 => x"5a",
          5490 => x"29",
          5491 => x"ff",
          5492 => x"f9",
          5493 => x"ff",
          5494 => x"42",
          5495 => x"7e",
          5496 => x"2e",
          5497 => x"80",
          5498 => x"89",
          5499 => x"39",
          5500 => x"33",
          5501 => x"2e",
          5502 => x"84",
          5503 => x"58",
          5504 => x"09",
          5505 => x"d9",
          5506 => x"83",
          5507 => x"fb",
          5508 => x"ba",
          5509 => x"75",
          5510 => x"be",
          5511 => x"d9",
          5512 => x"b5",
          5513 => x"05",
          5514 => x"33",
          5515 => x"5e",
          5516 => x"25",
          5517 => x"57",
          5518 => x"b5",
          5519 => x"39",
          5520 => x"33",
          5521 => x"2e",
          5522 => x"84",
          5523 => x"83",
          5524 => x"42",
          5525 => x"b8",
          5526 => x"11",
          5527 => x"75",
          5528 => x"38",
          5529 => x"83",
          5530 => x"fa",
          5531 => x"e5",
          5532 => x"e7",
          5533 => x"0b",
          5534 => x"33",
          5535 => x"76",
          5536 => x"38",
          5537 => x"ba",
          5538 => x"22",
          5539 => x"e5",
          5540 => x"e6",
          5541 => x"17",
          5542 => x"06",
          5543 => x"33",
          5544 => x"da",
          5545 => x"84",
          5546 => x"5f",
          5547 => x"2e",
          5548 => x"ba",
          5549 => x"75",
          5550 => x"38",
          5551 => x"52",
          5552 => x"06",
          5553 => x"3f",
          5554 => x"84",
          5555 => x"57",
          5556 => x"8e",
          5557 => x"ba",
          5558 => x"05",
          5559 => x"06",
          5560 => x"33",
          5561 => x"81",
          5562 => x"b8",
          5563 => x"81",
          5564 => x"11",
          5565 => x"5b",
          5566 => x"77",
          5567 => x"38",
          5568 => x"83",
          5569 => x"76",
          5570 => x"ff",
          5571 => x"77",
          5572 => x"38",
          5573 => x"83",
          5574 => x"84",
          5575 => x"ff",
          5576 => x"7a",
          5577 => x"b4",
          5578 => x"75",
          5579 => x"34",
          5580 => x"84",
          5581 => x"5f",
          5582 => x"8a",
          5583 => x"ba",
          5584 => x"b8",
          5585 => x"5b",
          5586 => x"f9",
          5587 => x"fa",
          5588 => x"b8",
          5589 => x"81",
          5590 => x"fa",
          5591 => x"74",
          5592 => x"c7",
          5593 => x"83",
          5594 => x"5f",
          5595 => x"29",
          5596 => x"ff",
          5597 => x"f9",
          5598 => x"52",
          5599 => x"5d",
          5600 => x"84",
          5601 => x"83",
          5602 => x"70",
          5603 => x"57",
          5604 => x"8e",
          5605 => x"b8",
          5606 => x"76",
          5607 => x"d6",
          5608 => x"56",
          5609 => x"b2",
          5610 => x"ff",
          5611 => x"31",
          5612 => x"60",
          5613 => x"38",
          5614 => x"33",
          5615 => x"27",
          5616 => x"ff",
          5617 => x"83",
          5618 => x"7e",
          5619 => x"83",
          5620 => x"57",
          5621 => x"76",
          5622 => x"38",
          5623 => x"81",
          5624 => x"ff",
          5625 => x"29",
          5626 => x"79",
          5627 => x"a0",
          5628 => x"c7",
          5629 => x"81",
          5630 => x"81",
          5631 => x"71",
          5632 => x"58",
          5633 => x"7f",
          5634 => x"38",
          5635 => x"1a",
          5636 => x"17",
          5637 => x"b9",
          5638 => x"7b",
          5639 => x"5d",
          5640 => x"81",
          5641 => x"7c",
          5642 => x"5e",
          5643 => x"84",
          5644 => x"84",
          5645 => x"71",
          5646 => x"43",
          5647 => x"77",
          5648 => x"9d",
          5649 => x"17",
          5650 => x"b9",
          5651 => x"7b",
          5652 => x"5d",
          5653 => x"81",
          5654 => x"7c",
          5655 => x"5e",
          5656 => x"84",
          5657 => x"84",
          5658 => x"71",
          5659 => x"43",
          5660 => x"7f",
          5661 => x"99",
          5662 => x"39",
          5663 => x"33",
          5664 => x"2e",
          5665 => x"80",
          5666 => x"d9",
          5667 => x"b1",
          5668 => x"39",
          5669 => x"b8",
          5670 => x"11",
          5671 => x"33",
          5672 => x"58",
          5673 => x"94",
          5674 => x"d8",
          5675 => x"78",
          5676 => x"06",
          5677 => x"83",
          5678 => x"58",
          5679 => x"06",
          5680 => x"33",
          5681 => x"5c",
          5682 => x"81",
          5683 => x"b8",
          5684 => x"7a",
          5685 => x"89",
          5686 => x"ff",
          5687 => x"76",
          5688 => x"38",
          5689 => x"61",
          5690 => x"57",
          5691 => x"38",
          5692 => x"1b",
          5693 => x"62",
          5694 => x"a0",
          5695 => x"1f",
          5696 => x"c7",
          5697 => x"79",
          5698 => x"51",
          5699 => x"ac",
          5700 => x"06",
          5701 => x"a4",
          5702 => x"b0",
          5703 => x"2b",
          5704 => x"07",
          5705 => x"07",
          5706 => x"7f",
          5707 => x"57",
          5708 => x"9e",
          5709 => x"70",
          5710 => x"0c",
          5711 => x"84",
          5712 => x"79",
          5713 => x"38",
          5714 => x"33",
          5715 => x"33",
          5716 => x"81",
          5717 => x"81",
          5718 => x"fa",
          5719 => x"73",
          5720 => x"59",
          5721 => x"77",
          5722 => x"38",
          5723 => x"1b",
          5724 => x"62",
          5725 => x"75",
          5726 => x"57",
          5727 => x"f4",
          5728 => x"fa",
          5729 => x"99",
          5730 => x"5a",
          5731 => x"e0",
          5732 => x"78",
          5733 => x"5a",
          5734 => x"57",
          5735 => x"f4",
          5736 => x"0b",
          5737 => x"34",
          5738 => x"81",
          5739 => x"81",
          5740 => x"77",
          5741 => x"f4",
          5742 => x"1f",
          5743 => x"06",
          5744 => x"8a",
          5745 => x"b0",
          5746 => x"f0",
          5747 => x"2b",
          5748 => x"71",
          5749 => x"58",
          5750 => x"80",
          5751 => x"81",
          5752 => x"80",
          5753 => x"fa",
          5754 => x"18",
          5755 => x"06",
          5756 => x"b6",
          5757 => x"b6",
          5758 => x"84",
          5759 => x"33",
          5760 => x"fa",
          5761 => x"b8",
          5762 => x"fa",
          5763 => x"b8",
          5764 => x"5c",
          5765 => x"ee",
          5766 => x"b0",
          5767 => x"56",
          5768 => x"b0",
          5769 => x"70",
          5770 => x"59",
          5771 => x"39",
          5772 => x"33",
          5773 => x"85",
          5774 => x"83",
          5775 => x"e5",
          5776 => x"b0",
          5777 => x"06",
          5778 => x"75",
          5779 => x"34",
          5780 => x"fa",
          5781 => x"f9",
          5782 => x"56",
          5783 => x"b0",
          5784 => x"83",
          5785 => x"81",
          5786 => x"07",
          5787 => x"fa",
          5788 => x"b1",
          5789 => x"0b",
          5790 => x"34",
          5791 => x"81",
          5792 => x"56",
          5793 => x"83",
          5794 => x"81",
          5795 => x"75",
          5796 => x"34",
          5797 => x"83",
          5798 => x"81",
          5799 => x"07",
          5800 => x"fa",
          5801 => x"fd",
          5802 => x"b0",
          5803 => x"06",
          5804 => x"56",
          5805 => x"b0",
          5806 => x"39",
          5807 => x"33",
          5808 => x"80",
          5809 => x"75",
          5810 => x"34",
          5811 => x"83",
          5812 => x"81",
          5813 => x"07",
          5814 => x"fa",
          5815 => x"c5",
          5816 => x"b0",
          5817 => x"06",
          5818 => x"75",
          5819 => x"34",
          5820 => x"83",
          5821 => x"81",
          5822 => x"07",
          5823 => x"fa",
          5824 => x"a1",
          5825 => x"b0",
          5826 => x"06",
          5827 => x"75",
          5828 => x"34",
          5829 => x"83",
          5830 => x"81",
          5831 => x"75",
          5832 => x"34",
          5833 => x"83",
          5834 => x"80",
          5835 => x"75",
          5836 => x"34",
          5837 => x"83",
          5838 => x"80",
          5839 => x"75",
          5840 => x"34",
          5841 => x"83",
          5842 => x"81",
          5843 => x"d0",
          5844 => x"83",
          5845 => x"fd",
          5846 => x"fa",
          5847 => x"bf",
          5848 => x"56",
          5849 => x"b0",
          5850 => x"39",
          5851 => x"fa",
          5852 => x"52",
          5853 => x"c9",
          5854 => x"39",
          5855 => x"33",
          5856 => x"34",
          5857 => x"33",
          5858 => x"34",
          5859 => x"33",
          5860 => x"fa",
          5861 => x"0b",
          5862 => x"0c",
          5863 => x"81",
          5864 => x"87",
          5865 => x"84",
          5866 => x"9c",
          5867 => x"77",
          5868 => x"34",
          5869 => x"33",
          5870 => x"06",
          5871 => x"56",
          5872 => x"84",
          5873 => x"9c",
          5874 => x"53",
          5875 => x"fe",
          5876 => x"84",
          5877 => x"a1",
          5878 => x"84",
          5879 => x"80",
          5880 => x"84",
          5881 => x"80",
          5882 => x"84",
          5883 => x"0d",
          5884 => x"fa",
          5885 => x"e9",
          5886 => x"85",
          5887 => x"5c",
          5888 => x"ba",
          5889 => x"10",
          5890 => x"5d",
          5891 => x"05",
          5892 => x"d8",
          5893 => x"0b",
          5894 => x"34",
          5895 => x"0b",
          5896 => x"34",
          5897 => x"51",
          5898 => x"83",
          5899 => x"70",
          5900 => x"58",
          5901 => x"e6",
          5902 => x"0b",
          5903 => x"34",
          5904 => x"51",
          5905 => x"ef",
          5906 => x"51",
          5907 => x"3f",
          5908 => x"83",
          5909 => x"ff",
          5910 => x"70",
          5911 => x"06",
          5912 => x"f2",
          5913 => x"52",
          5914 => x"39",
          5915 => x"33",
          5916 => x"27",
          5917 => x"75",
          5918 => x"34",
          5919 => x"83",
          5920 => x"ff",
          5921 => x"70",
          5922 => x"06",
          5923 => x"f0",
          5924 => x"fa",
          5925 => x"05",
          5926 => x"33",
          5927 => x"59",
          5928 => x"25",
          5929 => x"75",
          5930 => x"39",
          5931 => x"33",
          5932 => x"06",
          5933 => x"77",
          5934 => x"38",
          5935 => x"33",
          5936 => x"33",
          5937 => x"06",
          5938 => x"33",
          5939 => x"11",
          5940 => x"80",
          5941 => x"b2",
          5942 => x"71",
          5943 => x"70",
          5944 => x"06",
          5945 => x"33",
          5946 => x"42",
          5947 => x"81",
          5948 => x"38",
          5949 => x"ff",
          5950 => x"5c",
          5951 => x"24",
          5952 => x"84",
          5953 => x"56",
          5954 => x"83",
          5955 => x"16",
          5956 => x"fa",
          5957 => x"81",
          5958 => x"11",
          5959 => x"76",
          5960 => x"38",
          5961 => x"33",
          5962 => x"27",
          5963 => x"ff",
          5964 => x"83",
          5965 => x"7b",
          5966 => x"83",
          5967 => x"57",
          5968 => x"76",
          5969 => x"38",
          5970 => x"81",
          5971 => x"ff",
          5972 => x"29",
          5973 => x"79",
          5974 => x"a0",
          5975 => x"c7",
          5976 => x"81",
          5977 => x"81",
          5978 => x"71",
          5979 => x"42",
          5980 => x"7e",
          5981 => x"38",
          5982 => x"1a",
          5983 => x"17",
          5984 => x"b9",
          5985 => x"7b",
          5986 => x"5d",
          5987 => x"81",
          5988 => x"7d",
          5989 => x"5f",
          5990 => x"84",
          5991 => x"84",
          5992 => x"71",
          5993 => x"59",
          5994 => x"77",
          5995 => x"b1",
          5996 => x"17",
          5997 => x"b9",
          5998 => x"7b",
          5999 => x"5d",
          6000 => x"81",
          6001 => x"7d",
          6002 => x"5f",
          6003 => x"84",
          6004 => x"84",
          6005 => x"71",
          6006 => x"59",
          6007 => x"75",
          6008 => x"99",
          6009 => x"39",
          6010 => x"17",
          6011 => x"b9",
          6012 => x"7b",
          6013 => x"b4",
          6014 => x"f8",
          6015 => x"b2",
          6016 => x"f7",
          6017 => x"5f",
          6018 => x"39",
          6019 => x"38",
          6020 => x"33",
          6021 => x"06",
          6022 => x"42",
          6023 => x"27",
          6024 => x"5a",
          6025 => x"b2",
          6026 => x"ff",
          6027 => x"58",
          6028 => x"27",
          6029 => x"57",
          6030 => x"b4",
          6031 => x"f8",
          6032 => x"ff",
          6033 => x"52",
          6034 => x"78",
          6035 => x"38",
          6036 => x"83",
          6037 => x"eb",
          6038 => x"fa",
          6039 => x"05",
          6040 => x"33",
          6041 => x"40",
          6042 => x"25",
          6043 => x"75",
          6044 => x"39",
          6045 => x"09",
          6046 => x"c0",
          6047 => x"b5",
          6048 => x"ff",
          6049 => x"b4",
          6050 => x"5d",
          6051 => x"ff",
          6052 => x"06",
          6053 => x"f6",
          6054 => x"1d",
          6055 => x"fa",
          6056 => x"93",
          6057 => x"56",
          6058 => x"b2",
          6059 => x"39",
          6060 => x"56",
          6061 => x"b4",
          6062 => x"39",
          6063 => x"56",
          6064 => x"f5",
          6065 => x"76",
          6066 => x"58",
          6067 => x"b0",
          6068 => x"81",
          6069 => x"75",
          6070 => x"ec",
          6071 => x"70",
          6072 => x"34",
          6073 => x"33",
          6074 => x"05",
          6075 => x"76",
          6076 => x"f4",
          6077 => x"7b",
          6078 => x"83",
          6079 => x"f1",
          6080 => x"0b",
          6081 => x"34",
          6082 => x"7e",
          6083 => x"23",
          6084 => x"80",
          6085 => x"b2",
          6086 => x"39",
          6087 => x"fa",
          6088 => x"a7",
          6089 => x"b6",
          6090 => x"84",
          6091 => x"33",
          6092 => x"0b",
          6093 => x"34",
          6094 => x"fd",
          6095 => x"97",
          6096 => x"b8",
          6097 => x"54",
          6098 => x"90",
          6099 => x"db",
          6100 => x"0b",
          6101 => x"0c",
          6102 => x"04",
          6103 => x"51",
          6104 => x"80",
          6105 => x"84",
          6106 => x"0d",
          6107 => x"0d",
          6108 => x"33",
          6109 => x"83",
          6110 => x"70",
          6111 => x"83",
          6112 => x"33",
          6113 => x"59",
          6114 => x"80",
          6115 => x"14",
          6116 => x"f9",
          6117 => x"59",
          6118 => x"84",
          6119 => x"0d",
          6120 => x"e4",
          6121 => x"53",
          6122 => x"91",
          6123 => x"32",
          6124 => x"07",
          6125 => x"9f",
          6126 => x"5e",
          6127 => x"f8",
          6128 => x"59",
          6129 => x"81",
          6130 => x"06",
          6131 => x"54",
          6132 => x"70",
          6133 => x"25",
          6134 => x"5c",
          6135 => x"2e",
          6136 => x"84",
          6137 => x"83",
          6138 => x"83",
          6139 => x"72",
          6140 => x"86",
          6141 => x"05",
          6142 => x"22",
          6143 => x"71",
          6144 => x"70",
          6145 => x"06",
          6146 => x"33",
          6147 => x"58",
          6148 => x"83",
          6149 => x"f0",
          6150 => x"8e",
          6151 => x"80",
          6152 => x"98",
          6153 => x"c0",
          6154 => x"56",
          6155 => x"f6",
          6156 => x"80",
          6157 => x"76",
          6158 => x"15",
          6159 => x"70",
          6160 => x"55",
          6161 => x"74",
          6162 => x"80",
          6163 => x"a4",
          6164 => x"81",
          6165 => x"f8",
          6166 => x"58",
          6167 => x"76",
          6168 => x"38",
          6169 => x"2e",
          6170 => x"74",
          6171 => x"15",
          6172 => x"ff",
          6173 => x"81",
          6174 => x"cd",
          6175 => x"f8",
          6176 => x"83",
          6177 => x"33",
          6178 => x"15",
          6179 => x"70",
          6180 => x"55",
          6181 => x"27",
          6182 => x"83",
          6183 => x"70",
          6184 => x"80",
          6185 => x"54",
          6186 => x"dc",
          6187 => x"ff",
          6188 => x"2a",
          6189 => x"81",
          6190 => x"58",
          6191 => x"85",
          6192 => x"0b",
          6193 => x"34",
          6194 => x"06",
          6195 => x"2e",
          6196 => x"81",
          6197 => x"de",
          6198 => x"83",
          6199 => x"83",
          6200 => x"83",
          6201 => x"70",
          6202 => x"33",
          6203 => x"33",
          6204 => x"5e",
          6205 => x"83",
          6206 => x"33",
          6207 => x"ff",
          6208 => x"83",
          6209 => x"33",
          6210 => x"2e",
          6211 => x"83",
          6212 => x"33",
          6213 => x"ff",
          6214 => x"83",
          6215 => x"33",
          6216 => x"ec",
          6217 => x"ff",
          6218 => x"81",
          6219 => x"38",
          6220 => x"16",
          6221 => x"81",
          6222 => x"38",
          6223 => x"06",
          6224 => x"ff",
          6225 => x"38",
          6226 => x"16",
          6227 => x"74",
          6228 => x"38",
          6229 => x"08",
          6230 => x"87",
          6231 => x"08",
          6232 => x"73",
          6233 => x"38",
          6234 => x"c0",
          6235 => x"83",
          6236 => x"58",
          6237 => x"81",
          6238 => x"54",
          6239 => x"fe",
          6240 => x"83",
          6241 => x"77",
          6242 => x"34",
          6243 => x"53",
          6244 => x"82",
          6245 => x"10",
          6246 => x"fc",
          6247 => x"08",
          6248 => x"8c",
          6249 => x"80",
          6250 => x"83",
          6251 => x"c0",
          6252 => x"5e",
          6253 => x"27",
          6254 => x"80",
          6255 => x"8a",
          6256 => x"72",
          6257 => x"38",
          6258 => x"83",
          6259 => x"87",
          6260 => x"08",
          6261 => x"0c",
          6262 => x"06",
          6263 => x"2e",
          6264 => x"fa",
          6265 => x"54",
          6266 => x"14",
          6267 => x"81",
          6268 => x"a5",
          6269 => x"e4",
          6270 => x"80",
          6271 => x"38",
          6272 => x"83",
          6273 => x"c3",
          6274 => x"f0",
          6275 => x"39",
          6276 => x"e0",
          6277 => x"56",
          6278 => x"7c",
          6279 => x"38",
          6280 => x"09",
          6281 => x"b4",
          6282 => x"2e",
          6283 => x"79",
          6284 => x"d7",
          6285 => x"ff",
          6286 => x"77",
          6287 => x"2b",
          6288 => x"80",
          6289 => x"73",
          6290 => x"38",
          6291 => x"81",
          6292 => x"10",
          6293 => x"87",
          6294 => x"98",
          6295 => x"57",
          6296 => x"73",
          6297 => x"78",
          6298 => x"79",
          6299 => x"11",
          6300 => x"05",
          6301 => x"05",
          6302 => x"56",
          6303 => x"c0",
          6304 => x"83",
          6305 => x"57",
          6306 => x"80",
          6307 => x"2e",
          6308 => x"79",
          6309 => x"59",
          6310 => x"82",
          6311 => x"39",
          6312 => x"fa",
          6313 => x"0b",
          6314 => x"33",
          6315 => x"81",
          6316 => x"38",
          6317 => x"70",
          6318 => x"25",
          6319 => x"59",
          6320 => x"38",
          6321 => x"09",
          6322 => x"cc",
          6323 => x"2e",
          6324 => x"80",
          6325 => x"10",
          6326 => x"90",
          6327 => x"5d",
          6328 => x"2e",
          6329 => x"81",
          6330 => x"ff",
          6331 => x"93",
          6332 => x"38",
          6333 => x"33",
          6334 => x"2e",
          6335 => x"84",
          6336 => x"55",
          6337 => x"38",
          6338 => x"06",
          6339 => x"cc",
          6340 => x"84",
          6341 => x"8f",
          6342 => x"be",
          6343 => x"f0",
          6344 => x"39",
          6345 => x"2e",
          6346 => x"f8",
          6347 => x"81",
          6348 => x"83",
          6349 => x"34",
          6350 => x"80",
          6351 => x"cc",
          6352 => x"0b",
          6353 => x"15",
          6354 => x"83",
          6355 => x"34",
          6356 => x"74",
          6357 => x"53",
          6358 => x"2e",
          6359 => x"83",
          6360 => x"33",
          6361 => x"27",
          6362 => x"77",
          6363 => x"54",
          6364 => x"09",
          6365 => x"fc",
          6366 => x"d8",
          6367 => x"05",
          6368 => x"9c",
          6369 => x"74",
          6370 => x"e8",
          6371 => x"98",
          6372 => x"f8",
          6373 => x"81",
          6374 => x"fb",
          6375 => x"0b",
          6376 => x"15",
          6377 => x"39",
          6378 => x"dd",
          6379 => x"81",
          6380 => x"fa",
          6381 => x"83",
          6382 => x"80",
          6383 => x"dd",
          6384 => x"e4",
          6385 => x"de",
          6386 => x"f8",
          6387 => x"f8",
          6388 => x"5d",
          6389 => x"5e",
          6390 => x"39",
          6391 => x"09",
          6392 => x"cb",
          6393 => x"7a",
          6394 => x"ce",
          6395 => x"2e",
          6396 => x"fc",
          6397 => x"93",
          6398 => x"34",
          6399 => x"f8",
          6400 => x"0b",
          6401 => x"33",
          6402 => x"83",
          6403 => x"73",
          6404 => x"34",
          6405 => x"ac",
          6406 => x"84",
          6407 => x"58",
          6408 => x"38",
          6409 => x"84",
          6410 => x"ff",
          6411 => x"39",
          6412 => x"f8",
          6413 => x"2e",
          6414 => x"84",
          6415 => x"e4",
          6416 => x"39",
          6417 => x"33",
          6418 => x"06",
          6419 => x"5a",
          6420 => x"27",
          6421 => x"55",
          6422 => x"b2",
          6423 => x"ff",
          6424 => x"55",
          6425 => x"27",
          6426 => x"54",
          6427 => x"b4",
          6428 => x"f8",
          6429 => x"ff",
          6430 => x"05",
          6431 => x"27",
          6432 => x"53",
          6433 => x"b5",
          6434 => x"f6",
          6435 => x"52",
          6436 => x"ba",
          6437 => x"59",
          6438 => x"72",
          6439 => x"39",
          6440 => x"52",
          6441 => x"51",
          6442 => x"3f",
          6443 => x"f9",
          6444 => x"f8",
          6445 => x"fc",
          6446 => x"3d",
          6447 => x"f5",
          6448 => x"3d",
          6449 => x"3d",
          6450 => x"83",
          6451 => x"53",
          6452 => x"05",
          6453 => x"34",
          6454 => x"08",
          6455 => x"71",
          6456 => x"83",
          6457 => x"55",
          6458 => x"81",
          6459 => x"0b",
          6460 => x"e8",
          6461 => x"98",
          6462 => x"f5",
          6463 => x"80",
          6464 => x"53",
          6465 => x"9c",
          6466 => x"c0",
          6467 => x"51",
          6468 => x"f6",
          6469 => x"33",
          6470 => x"9c",
          6471 => x"74",
          6472 => x"38",
          6473 => x"2e",
          6474 => x"c0",
          6475 => x"51",
          6476 => x"73",
          6477 => x"38",
          6478 => x"ff",
          6479 => x"38",
          6480 => x"9c",
          6481 => x"90",
          6482 => x"c0",
          6483 => x"52",
          6484 => x"9c",
          6485 => x"72",
          6486 => x"81",
          6487 => x"c0",
          6488 => x"52",
          6489 => x"27",
          6490 => x"81",
          6491 => x"38",
          6492 => x"a4",
          6493 => x"75",
          6494 => x"ff",
          6495 => x"ff",
          6496 => x"ff",
          6497 => x"75",
          6498 => x"38",
          6499 => x"06",
          6500 => x"d5",
          6501 => x"2e",
          6502 => x"84",
          6503 => x"88",
          6504 => x"81",
          6505 => x"84",
          6506 => x"0d",
          6507 => x"0d",
          6508 => x"05",
          6509 => x"56",
          6510 => x"83",
          6511 => x"73",
          6512 => x"fc",
          6513 => x"70",
          6514 => x"07",
          6515 => x"57",
          6516 => x"34",
          6517 => x"51",
          6518 => x"34",
          6519 => x"56",
          6520 => x"34",
          6521 => x"34",
          6522 => x"08",
          6523 => x"13",
          6524 => x"90",
          6525 => x"e1",
          6526 => x"0b",
          6527 => x"08",
          6528 => x"0b",
          6529 => x"80",
          6530 => x"80",
          6531 => x"c0",
          6532 => x"83",
          6533 => x"55",
          6534 => x"05",
          6535 => x"98",
          6536 => x"87",
          6537 => x"08",
          6538 => x"2e",
          6539 => x"14",
          6540 => x"98",
          6541 => x"52",
          6542 => x"87",
          6543 => x"fe",
          6544 => x"87",
          6545 => x"08",
          6546 => x"70",
          6547 => x"c8",
          6548 => x"71",
          6549 => x"c0",
          6550 => x"98",
          6551 => x"ce",
          6552 => x"87",
          6553 => x"08",
          6554 => x"98",
          6555 => x"74",
          6556 => x"38",
          6557 => x"87",
          6558 => x"08",
          6559 => x"73",
          6560 => x"71",
          6561 => x"db",
          6562 => x"98",
          6563 => x"72",
          6564 => x"38",
          6565 => x"55",
          6566 => x"81",
          6567 => x"53",
          6568 => x"80",
          6569 => x"81",
          6570 => x"71",
          6571 => x"74",
          6572 => x"ff",
          6573 => x"aa",
          6574 => x"14",
          6575 => x"11",
          6576 => x"70",
          6577 => x"38",
          6578 => x"05",
          6579 => x"70",
          6580 => x"34",
          6581 => x"f0",
          6582 => x"bb",
          6583 => x"3d",
          6584 => x"0b",
          6585 => x"0c",
          6586 => x"04",
          6587 => x"39",
          6588 => x"79",
          6589 => x"a3",
          6590 => x"56",
          6591 => x"f5",
          6592 => x"88",
          6593 => x"80",
          6594 => x"79",
          6595 => x"51",
          6596 => x"75",
          6597 => x"72",
          6598 => x"70",
          6599 => x"75",
          6600 => x"71",
          6601 => x"72",
          6602 => x"7a",
          6603 => x"08",
          6604 => x"84",
          6605 => x"54",
          6606 => x"73",
          6607 => x"70",
          6608 => x"52",
          6609 => x"81",
          6610 => x"72",
          6611 => x"38",
          6612 => x"08",
          6613 => x"15",
          6614 => x"90",
          6615 => x"e2",
          6616 => x"0b",
          6617 => x"08",
          6618 => x"0b",
          6619 => x"80",
          6620 => x"80",
          6621 => x"c0",
          6622 => x"83",
          6623 => x"55",
          6624 => x"05",
          6625 => x"98",
          6626 => x"87",
          6627 => x"08",
          6628 => x"2e",
          6629 => x"14",
          6630 => x"98",
          6631 => x"52",
          6632 => x"87",
          6633 => x"fe",
          6634 => x"87",
          6635 => x"08",
          6636 => x"70",
          6637 => x"c8",
          6638 => x"71",
          6639 => x"c0",
          6640 => x"98",
          6641 => x"ce",
          6642 => x"87",
          6643 => x"08",
          6644 => x"98",
          6645 => x"74",
          6646 => x"38",
          6647 => x"87",
          6648 => x"08",
          6649 => x"73",
          6650 => x"71",
          6651 => x"db",
          6652 => x"98",
          6653 => x"72",
          6654 => x"38",
          6655 => x"55",
          6656 => x"81",
          6657 => x"53",
          6658 => x"a1",
          6659 => x"ff",
          6660 => x"fe",
          6661 => x"51",
          6662 => x"06",
          6663 => x"2e",
          6664 => x"57",
          6665 => x"84",
          6666 => x"0d",
          6667 => x"e8",
          6668 => x"0d",
          6669 => x"08",
          6670 => x"71",
          6671 => x"83",
          6672 => x"56",
          6673 => x"81",
          6674 => x"0b",
          6675 => x"e8",
          6676 => x"98",
          6677 => x"f5",
          6678 => x"80",
          6679 => x"54",
          6680 => x"9c",
          6681 => x"c0",
          6682 => x"53",
          6683 => x"f6",
          6684 => x"33",
          6685 => x"9c",
          6686 => x"70",
          6687 => x"38",
          6688 => x"2e",
          6689 => x"c0",
          6690 => x"51",
          6691 => x"74",
          6692 => x"38",
          6693 => x"ff",
          6694 => x"38",
          6695 => x"9c",
          6696 => x"90",
          6697 => x"c0",
          6698 => x"52",
          6699 => x"9c",
          6700 => x"72",
          6701 => x"81",
          6702 => x"c0",
          6703 => x"55",
          6704 => x"27",
          6705 => x"81",
          6706 => x"38",
          6707 => x"a4",
          6708 => x"71",
          6709 => x"ff",
          6710 => x"ff",
          6711 => x"ff",
          6712 => x"75",
          6713 => x"38",
          6714 => x"06",
          6715 => x"d5",
          6716 => x"80",
          6717 => x"e6",
          6718 => x"ce",
          6719 => x"3d",
          6720 => x"3d",
          6721 => x"f4",
          6722 => x"31",
          6723 => x"83",
          6724 => x"70",
          6725 => x"11",
          6726 => x"12",
          6727 => x"2b",
          6728 => x"07",
          6729 => x"33",
          6730 => x"71",
          6731 => x"90",
          6732 => x"54",
          6733 => x"5d",
          6734 => x"56",
          6735 => x"71",
          6736 => x"38",
          6737 => x"11",
          6738 => x"33",
          6739 => x"71",
          6740 => x"76",
          6741 => x"81",
          6742 => x"98",
          6743 => x"2b",
          6744 => x"5c",
          6745 => x"52",
          6746 => x"83",
          6747 => x"13",
          6748 => x"33",
          6749 => x"71",
          6750 => x"75",
          6751 => x"2a",
          6752 => x"57",
          6753 => x"34",
          6754 => x"06",
          6755 => x"13",
          6756 => x"f4",
          6757 => x"84",
          6758 => x"13",
          6759 => x"2b",
          6760 => x"2a",
          6761 => x"54",
          6762 => x"14",
          6763 => x"14",
          6764 => x"f4",
          6765 => x"80",
          6766 => x"34",
          6767 => x"13",
          6768 => x"f4",
          6769 => x"84",
          6770 => x"85",
          6771 => x"ba",
          6772 => x"70",
          6773 => x"33",
          6774 => x"07",
          6775 => x"07",
          6776 => x"58",
          6777 => x"74",
          6778 => x"81",
          6779 => x"3d",
          6780 => x"12",
          6781 => x"33",
          6782 => x"71",
          6783 => x"75",
          6784 => x"33",
          6785 => x"71",
          6786 => x"70",
          6787 => x"58",
          6788 => x"58",
          6789 => x"12",
          6790 => x"12",
          6791 => x"f4",
          6792 => x"84",
          6793 => x"12",
          6794 => x"2b",
          6795 => x"07",
          6796 => x"52",
          6797 => x"12",
          6798 => x"33",
          6799 => x"07",
          6800 => x"52",
          6801 => x"77",
          6802 => x"72",
          6803 => x"84",
          6804 => x"15",
          6805 => x"12",
          6806 => x"2b",
          6807 => x"ff",
          6808 => x"2a",
          6809 => x"52",
          6810 => x"77",
          6811 => x"84",
          6812 => x"70",
          6813 => x"81",
          6814 => x"8b",
          6815 => x"2b",
          6816 => x"70",
          6817 => x"33",
          6818 => x"07",
          6819 => x"8f",
          6820 => x"77",
          6821 => x"2a",
          6822 => x"54",
          6823 => x"54",
          6824 => x"14",
          6825 => x"14",
          6826 => x"f4",
          6827 => x"70",
          6828 => x"33",
          6829 => x"71",
          6830 => x"74",
          6831 => x"81",
          6832 => x"88",
          6833 => x"ff",
          6834 => x"88",
          6835 => x"53",
          6836 => x"54",
          6837 => x"34",
          6838 => x"34",
          6839 => x"08",
          6840 => x"11",
          6841 => x"33",
          6842 => x"71",
          6843 => x"74",
          6844 => x"81",
          6845 => x"98",
          6846 => x"2b",
          6847 => x"5d",
          6848 => x"53",
          6849 => x"25",
          6850 => x"71",
          6851 => x"33",
          6852 => x"07",
          6853 => x"07",
          6854 => x"59",
          6855 => x"75",
          6856 => x"16",
          6857 => x"f4",
          6858 => x"70",
          6859 => x"33",
          6860 => x"71",
          6861 => x"74",
          6862 => x"33",
          6863 => x"71",
          6864 => x"70",
          6865 => x"5c",
          6866 => x"56",
          6867 => x"82",
          6868 => x"83",
          6869 => x"3d",
          6870 => x"3d",
          6871 => x"ba",
          6872 => x"58",
          6873 => x"8f",
          6874 => x"2e",
          6875 => x"51",
          6876 => x"89",
          6877 => x"84",
          6878 => x"84",
          6879 => x"a0",
          6880 => x"ba",
          6881 => x"80",
          6882 => x"52",
          6883 => x"51",
          6884 => x"3f",
          6885 => x"08",
          6886 => x"34",
          6887 => x"16",
          6888 => x"f4",
          6889 => x"84",
          6890 => x"0b",
          6891 => x"84",
          6892 => x"56",
          6893 => x"34",
          6894 => x"17",
          6895 => x"f4",
          6896 => x"f0",
          6897 => x"fe",
          6898 => x"70",
          6899 => x"06",
          6900 => x"58",
          6901 => x"74",
          6902 => x"73",
          6903 => x"84",
          6904 => x"70",
          6905 => x"84",
          6906 => x"05",
          6907 => x"55",
          6908 => x"34",
          6909 => x"15",
          6910 => x"39",
          6911 => x"7b",
          6912 => x"81",
          6913 => x"27",
          6914 => x"12",
          6915 => x"05",
          6916 => x"ff",
          6917 => x"70",
          6918 => x"06",
          6919 => x"08",
          6920 => x"85",
          6921 => x"88",
          6922 => x"52",
          6923 => x"55",
          6924 => x"54",
          6925 => x"80",
          6926 => x"10",
          6927 => x"70",
          6928 => x"33",
          6929 => x"07",
          6930 => x"ff",
          6931 => x"70",
          6932 => x"06",
          6933 => x"56",
          6934 => x"54",
          6935 => x"27",
          6936 => x"80",
          6937 => x"75",
          6938 => x"84",
          6939 => x"13",
          6940 => x"2b",
          6941 => x"75",
          6942 => x"81",
          6943 => x"85",
          6944 => x"54",
          6945 => x"83",
          6946 => x"70",
          6947 => x"33",
          6948 => x"07",
          6949 => x"ff",
          6950 => x"5d",
          6951 => x"70",
          6952 => x"38",
          6953 => x"51",
          6954 => x"82",
          6955 => x"51",
          6956 => x"82",
          6957 => x"75",
          6958 => x"38",
          6959 => x"83",
          6960 => x"74",
          6961 => x"07",
          6962 => x"5b",
          6963 => x"5a",
          6964 => x"78",
          6965 => x"84",
          6966 => x"15",
          6967 => x"53",
          6968 => x"14",
          6969 => x"14",
          6970 => x"f4",
          6971 => x"70",
          6972 => x"33",
          6973 => x"07",
          6974 => x"8f",
          6975 => x"74",
          6976 => x"ff",
          6977 => x"88",
          6978 => x"53",
          6979 => x"52",
          6980 => x"34",
          6981 => x"06",
          6982 => x"12",
          6983 => x"f4",
          6984 => x"75",
          6985 => x"81",
          6986 => x"ba",
          6987 => x"19",
          6988 => x"87",
          6989 => x"8b",
          6990 => x"2b",
          6991 => x"58",
          6992 => x"57",
          6993 => x"34",
          6994 => x"34",
          6995 => x"08",
          6996 => x"78",
          6997 => x"33",
          6998 => x"71",
          6999 => x"70",
          7000 => x"54",
          7001 => x"86",
          7002 => x"87",
          7003 => x"ba",
          7004 => x"19",
          7005 => x"85",
          7006 => x"8b",
          7007 => x"2b",
          7008 => x"58",
          7009 => x"52",
          7010 => x"34",
          7011 => x"34",
          7012 => x"08",
          7013 => x"78",
          7014 => x"33",
          7015 => x"71",
          7016 => x"70",
          7017 => x"5c",
          7018 => x"84",
          7019 => x"85",
          7020 => x"ba",
          7021 => x"84",
          7022 => x"84",
          7023 => x"8b",
          7024 => x"86",
          7025 => x"15",
          7026 => x"2b",
          7027 => x"07",
          7028 => x"17",
          7029 => x"33",
          7030 => x"07",
          7031 => x"5a",
          7032 => x"54",
          7033 => x"12",
          7034 => x"12",
          7035 => x"f4",
          7036 => x"84",
          7037 => x"12",
          7038 => x"2b",
          7039 => x"07",
          7040 => x"14",
          7041 => x"33",
          7042 => x"07",
          7043 => x"58",
          7044 => x"56",
          7045 => x"70",
          7046 => x"76",
          7047 => x"84",
          7048 => x"18",
          7049 => x"12",
          7050 => x"2b",
          7051 => x"ff",
          7052 => x"2a",
          7053 => x"57",
          7054 => x"74",
          7055 => x"84",
          7056 => x"18",
          7057 => x"fe",
          7058 => x"3d",
          7059 => x"ba",
          7060 => x"58",
          7061 => x"a0",
          7062 => x"77",
          7063 => x"84",
          7064 => x"89",
          7065 => x"77",
          7066 => x"3f",
          7067 => x"08",
          7068 => x"0c",
          7069 => x"04",
          7070 => x"0b",
          7071 => x"0c",
          7072 => x"84",
          7073 => x"82",
          7074 => x"76",
          7075 => x"f4",
          7076 => x"ec",
          7077 => x"f4",
          7078 => x"75",
          7079 => x"81",
          7080 => x"ba",
          7081 => x"76",
          7082 => x"81",
          7083 => x"34",
          7084 => x"08",
          7085 => x"17",
          7086 => x"87",
          7087 => x"ba",
          7088 => x"ba",
          7089 => x"05",
          7090 => x"07",
          7091 => x"ff",
          7092 => x"2a",
          7093 => x"56",
          7094 => x"34",
          7095 => x"34",
          7096 => x"22",
          7097 => x"10",
          7098 => x"08",
          7099 => x"55",
          7100 => x"15",
          7101 => x"83",
          7102 => x"54",
          7103 => x"fe",
          7104 => x"e3",
          7105 => x"0d",
          7106 => x"5f",
          7107 => x"ba",
          7108 => x"45",
          7109 => x"2e",
          7110 => x"7e",
          7111 => x"af",
          7112 => x"2e",
          7113 => x"81",
          7114 => x"27",
          7115 => x"fb",
          7116 => x"82",
          7117 => x"ff",
          7118 => x"58",
          7119 => x"ff",
          7120 => x"31",
          7121 => x"83",
          7122 => x"70",
          7123 => x"11",
          7124 => x"12",
          7125 => x"2b",
          7126 => x"31",
          7127 => x"ff",
          7128 => x"10",
          7129 => x"73",
          7130 => x"11",
          7131 => x"12",
          7132 => x"2b",
          7133 => x"2b",
          7134 => x"53",
          7135 => x"44",
          7136 => x"44",
          7137 => x"52",
          7138 => x"80",
          7139 => x"fd",
          7140 => x"33",
          7141 => x"71",
          7142 => x"70",
          7143 => x"19",
          7144 => x"12",
          7145 => x"2b",
          7146 => x"07",
          7147 => x"56",
          7148 => x"74",
          7149 => x"38",
          7150 => x"82",
          7151 => x"1b",
          7152 => x"2e",
          7153 => x"60",
          7154 => x"f9",
          7155 => x"58",
          7156 => x"87",
          7157 => x"18",
          7158 => x"24",
          7159 => x"76",
          7160 => x"81",
          7161 => x"8b",
          7162 => x"2b",
          7163 => x"70",
          7164 => x"33",
          7165 => x"71",
          7166 => x"47",
          7167 => x"53",
          7168 => x"80",
          7169 => x"ba",
          7170 => x"82",
          7171 => x"12",
          7172 => x"2b",
          7173 => x"07",
          7174 => x"11",
          7175 => x"33",
          7176 => x"71",
          7177 => x"7e",
          7178 => x"33",
          7179 => x"71",
          7180 => x"70",
          7181 => x"57",
          7182 => x"41",
          7183 => x"59",
          7184 => x"1d",
          7185 => x"1d",
          7186 => x"f4",
          7187 => x"84",
          7188 => x"12",
          7189 => x"2b",
          7190 => x"07",
          7191 => x"14",
          7192 => x"33",
          7193 => x"07",
          7194 => x"5f",
          7195 => x"40",
          7196 => x"77",
          7197 => x"7b",
          7198 => x"84",
          7199 => x"16",
          7200 => x"12",
          7201 => x"2b",
          7202 => x"ff",
          7203 => x"2a",
          7204 => x"59",
          7205 => x"79",
          7206 => x"84",
          7207 => x"70",
          7208 => x"33",
          7209 => x"71",
          7210 => x"83",
          7211 => x"05",
          7212 => x"15",
          7213 => x"2b",
          7214 => x"2a",
          7215 => x"5d",
          7216 => x"55",
          7217 => x"75",
          7218 => x"84",
          7219 => x"70",
          7220 => x"81",
          7221 => x"8b",
          7222 => x"2b",
          7223 => x"82",
          7224 => x"15",
          7225 => x"2b",
          7226 => x"2a",
          7227 => x"5d",
          7228 => x"55",
          7229 => x"34",
          7230 => x"34",
          7231 => x"08",
          7232 => x"11",
          7233 => x"33",
          7234 => x"07",
          7235 => x"56",
          7236 => x"42",
          7237 => x"7e",
          7238 => x"51",
          7239 => x"3f",
          7240 => x"08",
          7241 => x"61",
          7242 => x"70",
          7243 => x"06",
          7244 => x"7a",
          7245 => x"b6",
          7246 => x"73",
          7247 => x"0c",
          7248 => x"04",
          7249 => x"0b",
          7250 => x"0c",
          7251 => x"84",
          7252 => x"82",
          7253 => x"60",
          7254 => x"f4",
          7255 => x"a0",
          7256 => x"f4",
          7257 => x"7e",
          7258 => x"81",
          7259 => x"ba",
          7260 => x"60",
          7261 => x"81",
          7262 => x"34",
          7263 => x"08",
          7264 => x"1d",
          7265 => x"87",
          7266 => x"ba",
          7267 => x"ba",
          7268 => x"05",
          7269 => x"07",
          7270 => x"ff",
          7271 => x"2a",
          7272 => x"57",
          7273 => x"34",
          7274 => x"34",
          7275 => x"22",
          7276 => x"10",
          7277 => x"08",
          7278 => x"55",
          7279 => x"15",
          7280 => x"83",
          7281 => x"ba",
          7282 => x"7e",
          7283 => x"76",
          7284 => x"8c",
          7285 => x"7f",
          7286 => x"df",
          7287 => x"f4",
          7288 => x"bb",
          7289 => x"bb",
          7290 => x"3d",
          7291 => x"1c",
          7292 => x"08",
          7293 => x"71",
          7294 => x"7f",
          7295 => x"81",
          7296 => x"88",
          7297 => x"ff",
          7298 => x"88",
          7299 => x"5b",
          7300 => x"7b",
          7301 => x"1c",
          7302 => x"ba",
          7303 => x"7c",
          7304 => x"58",
          7305 => x"34",
          7306 => x"34",
          7307 => x"08",
          7308 => x"33",
          7309 => x"71",
          7310 => x"70",
          7311 => x"ff",
          7312 => x"05",
          7313 => x"ff",
          7314 => x"2a",
          7315 => x"57",
          7316 => x"63",
          7317 => x"34",
          7318 => x"06",
          7319 => x"83",
          7320 => x"ba",
          7321 => x"5b",
          7322 => x"60",
          7323 => x"61",
          7324 => x"08",
          7325 => x"51",
          7326 => x"7e",
          7327 => x"39",
          7328 => x"70",
          7329 => x"06",
          7330 => x"ac",
          7331 => x"ff",
          7332 => x"31",
          7333 => x"ff",
          7334 => x"33",
          7335 => x"71",
          7336 => x"70",
          7337 => x"1b",
          7338 => x"12",
          7339 => x"2b",
          7340 => x"07",
          7341 => x"54",
          7342 => x"54",
          7343 => x"f9",
          7344 => x"bc",
          7345 => x"24",
          7346 => x"80",
          7347 => x"8f",
          7348 => x"ff",
          7349 => x"61",
          7350 => x"dd",
          7351 => x"39",
          7352 => x"0b",
          7353 => x"0c",
          7354 => x"84",
          7355 => x"82",
          7356 => x"7e",
          7357 => x"f4",
          7358 => x"84",
          7359 => x"f4",
          7360 => x"7a",
          7361 => x"81",
          7362 => x"ba",
          7363 => x"7e",
          7364 => x"81",
          7365 => x"34",
          7366 => x"08",
          7367 => x"19",
          7368 => x"87",
          7369 => x"ba",
          7370 => x"ba",
          7371 => x"05",
          7372 => x"07",
          7373 => x"ff",
          7374 => x"2a",
          7375 => x"44",
          7376 => x"05",
          7377 => x"89",
          7378 => x"ba",
          7379 => x"10",
          7380 => x"ba",
          7381 => x"f8",
          7382 => x"7e",
          7383 => x"34",
          7384 => x"05",
          7385 => x"39",
          7386 => x"83",
          7387 => x"83",
          7388 => x"5b",
          7389 => x"fb",
          7390 => x"f2",
          7391 => x"2e",
          7392 => x"7e",
          7393 => x"3f",
          7394 => x"84",
          7395 => x"95",
          7396 => x"76",
          7397 => x"33",
          7398 => x"71",
          7399 => x"83",
          7400 => x"11",
          7401 => x"87",
          7402 => x"8b",
          7403 => x"2b",
          7404 => x"84",
          7405 => x"15",
          7406 => x"2b",
          7407 => x"2a",
          7408 => x"56",
          7409 => x"53",
          7410 => x"78",
          7411 => x"34",
          7412 => x"05",
          7413 => x"f4",
          7414 => x"84",
          7415 => x"12",
          7416 => x"2b",
          7417 => x"07",
          7418 => x"14",
          7419 => x"33",
          7420 => x"07",
          7421 => x"5b",
          7422 => x"5d",
          7423 => x"73",
          7424 => x"34",
          7425 => x"05",
          7426 => x"f4",
          7427 => x"33",
          7428 => x"71",
          7429 => x"81",
          7430 => x"70",
          7431 => x"5c",
          7432 => x"7d",
          7433 => x"1e",
          7434 => x"f4",
          7435 => x"82",
          7436 => x"12",
          7437 => x"2b",
          7438 => x"07",
          7439 => x"33",
          7440 => x"71",
          7441 => x"70",
          7442 => x"5c",
          7443 => x"57",
          7444 => x"7c",
          7445 => x"1d",
          7446 => x"f4",
          7447 => x"70",
          7448 => x"33",
          7449 => x"71",
          7450 => x"74",
          7451 => x"33",
          7452 => x"71",
          7453 => x"70",
          7454 => x"47",
          7455 => x"5c",
          7456 => x"82",
          7457 => x"83",
          7458 => x"ba",
          7459 => x"1f",
          7460 => x"83",
          7461 => x"88",
          7462 => x"57",
          7463 => x"83",
          7464 => x"58",
          7465 => x"84",
          7466 => x"bc",
          7467 => x"ba",
          7468 => x"84",
          7469 => x"ff",
          7470 => x"5f",
          7471 => x"84",
          7472 => x"84",
          7473 => x"a0",
          7474 => x"ba",
          7475 => x"80",
          7476 => x"52",
          7477 => x"51",
          7478 => x"3f",
          7479 => x"08",
          7480 => x"34",
          7481 => x"17",
          7482 => x"f4",
          7483 => x"84",
          7484 => x"0b",
          7485 => x"84",
          7486 => x"54",
          7487 => x"34",
          7488 => x"15",
          7489 => x"f4",
          7490 => x"f0",
          7491 => x"fe",
          7492 => x"70",
          7493 => x"06",
          7494 => x"45",
          7495 => x"61",
          7496 => x"60",
          7497 => x"84",
          7498 => x"70",
          7499 => x"84",
          7500 => x"05",
          7501 => x"5d",
          7502 => x"34",
          7503 => x"1c",
          7504 => x"e7",
          7505 => x"54",
          7506 => x"86",
          7507 => x"1a",
          7508 => x"2b",
          7509 => x"07",
          7510 => x"1c",
          7511 => x"33",
          7512 => x"07",
          7513 => x"5c",
          7514 => x"59",
          7515 => x"84",
          7516 => x"61",
          7517 => x"84",
          7518 => x"70",
          7519 => x"33",
          7520 => x"71",
          7521 => x"83",
          7522 => x"05",
          7523 => x"87",
          7524 => x"88",
          7525 => x"88",
          7526 => x"48",
          7527 => x"59",
          7528 => x"86",
          7529 => x"64",
          7530 => x"84",
          7531 => x"1d",
          7532 => x"12",
          7533 => x"2b",
          7534 => x"ff",
          7535 => x"2a",
          7536 => x"58",
          7537 => x"7f",
          7538 => x"84",
          7539 => x"70",
          7540 => x"81",
          7541 => x"8b",
          7542 => x"2b",
          7543 => x"70",
          7544 => x"33",
          7545 => x"07",
          7546 => x"8f",
          7547 => x"77",
          7548 => x"2a",
          7549 => x"5a",
          7550 => x"44",
          7551 => x"17",
          7552 => x"17",
          7553 => x"f4",
          7554 => x"70",
          7555 => x"33",
          7556 => x"71",
          7557 => x"74",
          7558 => x"81",
          7559 => x"88",
          7560 => x"ff",
          7561 => x"88",
          7562 => x"5e",
          7563 => x"41",
          7564 => x"34",
          7565 => x"05",
          7566 => x"ff",
          7567 => x"fa",
          7568 => x"15",
          7569 => x"33",
          7570 => x"71",
          7571 => x"79",
          7572 => x"33",
          7573 => x"71",
          7574 => x"70",
          7575 => x"5e",
          7576 => x"5d",
          7577 => x"34",
          7578 => x"34",
          7579 => x"08",
          7580 => x"11",
          7581 => x"33",
          7582 => x"71",
          7583 => x"74",
          7584 => x"33",
          7585 => x"71",
          7586 => x"70",
          7587 => x"56",
          7588 => x"42",
          7589 => x"60",
          7590 => x"75",
          7591 => x"34",
          7592 => x"08",
          7593 => x"81",
          7594 => x"88",
          7595 => x"ff",
          7596 => x"88",
          7597 => x"58",
          7598 => x"34",
          7599 => x"34",
          7600 => x"08",
          7601 => x"33",
          7602 => x"71",
          7603 => x"83",
          7604 => x"05",
          7605 => x"12",
          7606 => x"2b",
          7607 => x"2b",
          7608 => x"06",
          7609 => x"88",
          7610 => x"5f",
          7611 => x"42",
          7612 => x"82",
          7613 => x"83",
          7614 => x"ba",
          7615 => x"1f",
          7616 => x"12",
          7617 => x"2b",
          7618 => x"07",
          7619 => x"33",
          7620 => x"71",
          7621 => x"81",
          7622 => x"70",
          7623 => x"54",
          7624 => x"59",
          7625 => x"7c",
          7626 => x"1d",
          7627 => x"f4",
          7628 => x"82",
          7629 => x"12",
          7630 => x"2b",
          7631 => x"07",
          7632 => x"11",
          7633 => x"33",
          7634 => x"71",
          7635 => x"78",
          7636 => x"33",
          7637 => x"71",
          7638 => x"70",
          7639 => x"57",
          7640 => x"42",
          7641 => x"5a",
          7642 => x"84",
          7643 => x"85",
          7644 => x"ba",
          7645 => x"17",
          7646 => x"85",
          7647 => x"8b",
          7648 => x"2b",
          7649 => x"86",
          7650 => x"15",
          7651 => x"2b",
          7652 => x"2a",
          7653 => x"52",
          7654 => x"57",
          7655 => x"34",
          7656 => x"34",
          7657 => x"08",
          7658 => x"81",
          7659 => x"88",
          7660 => x"ff",
          7661 => x"88",
          7662 => x"5e",
          7663 => x"34",
          7664 => x"34",
          7665 => x"08",
          7666 => x"11",
          7667 => x"33",
          7668 => x"71",
          7669 => x"74",
          7670 => x"81",
          7671 => x"88",
          7672 => x"88",
          7673 => x"45",
          7674 => x"55",
          7675 => x"34",
          7676 => x"34",
          7677 => x"08",
          7678 => x"33",
          7679 => x"71",
          7680 => x"83",
          7681 => x"05",
          7682 => x"83",
          7683 => x"88",
          7684 => x"88",
          7685 => x"45",
          7686 => x"55",
          7687 => x"1a",
          7688 => x"1a",
          7689 => x"f4",
          7690 => x"82",
          7691 => x"12",
          7692 => x"2b",
          7693 => x"62",
          7694 => x"2b",
          7695 => x"5d",
          7696 => x"05",
          7697 => x"fb",
          7698 => x"f4",
          7699 => x"05",
          7700 => x"1c",
          7701 => x"ff",
          7702 => x"5f",
          7703 => x"86",
          7704 => x"1a",
          7705 => x"2b",
          7706 => x"07",
          7707 => x"1c",
          7708 => x"33",
          7709 => x"07",
          7710 => x"40",
          7711 => x"41",
          7712 => x"84",
          7713 => x"61",
          7714 => x"84",
          7715 => x"70",
          7716 => x"33",
          7717 => x"71",
          7718 => x"83",
          7719 => x"05",
          7720 => x"87",
          7721 => x"88",
          7722 => x"88",
          7723 => x"5f",
          7724 => x"41",
          7725 => x"86",
          7726 => x"64",
          7727 => x"84",
          7728 => x"1d",
          7729 => x"12",
          7730 => x"2b",
          7731 => x"ff",
          7732 => x"2a",
          7733 => x"55",
          7734 => x"7c",
          7735 => x"84",
          7736 => x"70",
          7737 => x"81",
          7738 => x"8b",
          7739 => x"2b",
          7740 => x"70",
          7741 => x"33",
          7742 => x"07",
          7743 => x"8f",
          7744 => x"77",
          7745 => x"2a",
          7746 => x"49",
          7747 => x"58",
          7748 => x"1e",
          7749 => x"1e",
          7750 => x"f4",
          7751 => x"70",
          7752 => x"33",
          7753 => x"71",
          7754 => x"74",
          7755 => x"81",
          7756 => x"88",
          7757 => x"ff",
          7758 => x"88",
          7759 => x"49",
          7760 => x"5e",
          7761 => x"34",
          7762 => x"34",
          7763 => x"ff",
          7764 => x"83",
          7765 => x"52",
          7766 => x"3f",
          7767 => x"08",
          7768 => x"84",
          7769 => x"93",
          7770 => x"73",
          7771 => x"84",
          7772 => x"b3",
          7773 => x"51",
          7774 => x"61",
          7775 => x"27",
          7776 => x"f0",
          7777 => x"3d",
          7778 => x"29",
          7779 => x"08",
          7780 => x"80",
          7781 => x"77",
          7782 => x"38",
          7783 => x"84",
          7784 => x"0d",
          7785 => x"e4",
          7786 => x"bb",
          7787 => x"84",
          7788 => x"80",
          7789 => x"77",
          7790 => x"84",
          7791 => x"51",
          7792 => x"3f",
          7793 => x"84",
          7794 => x"0d",
          7795 => x"f4",
          7796 => x"f4",
          7797 => x"0b",
          7798 => x"23",
          7799 => x"53",
          7800 => x"ff",
          7801 => x"b5",
          7802 => x"ba",
          7803 => x"76",
          7804 => x"0b",
          7805 => x"84",
          7806 => x"54",
          7807 => x"34",
          7808 => x"15",
          7809 => x"f4",
          7810 => x"86",
          7811 => x"0b",
          7812 => x"84",
          7813 => x"84",
          7814 => x"ff",
          7815 => x"80",
          7816 => x"ff",
          7817 => x"88",
          7818 => x"55",
          7819 => x"17",
          7820 => x"17",
          7821 => x"f0",
          7822 => x"10",
          7823 => x"f4",
          7824 => x"05",
          7825 => x"82",
          7826 => x"0b",
          7827 => x"77",
          7828 => x"2e",
          7829 => x"fe",
          7830 => x"3d",
          7831 => x"05",
          7832 => x"52",
          7833 => x"87",
          7834 => x"80",
          7835 => x"71",
          7836 => x"0c",
          7837 => x"04",
          7838 => x"02",
          7839 => x"52",
          7840 => x"81",
          7841 => x"71",
          7842 => x"3f",
          7843 => x"08",
          7844 => x"53",
          7845 => x"72",
          7846 => x"13",
          7847 => x"80",
          7848 => x"72",
          7849 => x"0c",
          7850 => x"04",
          7851 => x"7c",
          7852 => x"8c",
          7853 => x"33",
          7854 => x"59",
          7855 => x"74",
          7856 => x"84",
          7857 => x"33",
          7858 => x"06",
          7859 => x"73",
          7860 => x"58",
          7861 => x"c0",
          7862 => x"78",
          7863 => x"76",
          7864 => x"3f",
          7865 => x"08",
          7866 => x"55",
          7867 => x"a7",
          7868 => x"98",
          7869 => x"73",
          7870 => x"78",
          7871 => x"74",
          7872 => x"06",
          7873 => x"2e",
          7874 => x"54",
          7875 => x"84",
          7876 => x"8b",
          7877 => x"84",
          7878 => x"19",
          7879 => x"06",
          7880 => x"79",
          7881 => x"ac",
          7882 => x"f7",
          7883 => x"7e",
          7884 => x"05",
          7885 => x"5a",
          7886 => x"81",
          7887 => x"26",
          7888 => x"bb",
          7889 => x"54",
          7890 => x"54",
          7891 => x"bd",
          7892 => x"85",
          7893 => x"98",
          7894 => x"53",
          7895 => x"51",
          7896 => x"84",
          7897 => x"81",
          7898 => x"74",
          7899 => x"38",
          7900 => x"8c",
          7901 => x"e2",
          7902 => x"26",
          7903 => x"fc",
          7904 => x"54",
          7905 => x"83",
          7906 => x"73",
          7907 => x"bb",
          7908 => x"3d",
          7909 => x"80",
          7910 => x"70",
          7911 => x"5a",
          7912 => x"78",
          7913 => x"38",
          7914 => x"3d",
          7915 => x"84",
          7916 => x"33",
          7917 => x"9f",
          7918 => x"53",
          7919 => x"71",
          7920 => x"38",
          7921 => x"12",
          7922 => x"81",
          7923 => x"53",
          7924 => x"85",
          7925 => x"98",
          7926 => x"53",
          7927 => x"96",
          7928 => x"25",
          7929 => x"83",
          7930 => x"84",
          7931 => x"bb",
          7932 => x"3d",
          7933 => x"80",
          7934 => x"73",
          7935 => x"0c",
          7936 => x"04",
          7937 => x"0c",
          7938 => x"bb",
          7939 => x"3d",
          7940 => x"84",
          7941 => x"92",
          7942 => x"54",
          7943 => x"71",
          7944 => x"2a",
          7945 => x"51",
          7946 => x"8a",
          7947 => x"98",
          7948 => x"74",
          7949 => x"c0",
          7950 => x"51",
          7951 => x"81",
          7952 => x"c0",
          7953 => x"52",
          7954 => x"06",
          7955 => x"2e",
          7956 => x"71",
          7957 => x"54",
          7958 => x"ff",
          7959 => x"3d",
          7960 => x"80",
          7961 => x"33",
          7962 => x"57",
          7963 => x"09",
          7964 => x"38",
          7965 => x"75",
          7966 => x"87",
          7967 => x"80",
          7968 => x"33",
          7969 => x"3f",
          7970 => x"08",
          7971 => x"38",
          7972 => x"84",
          7973 => x"8c",
          7974 => x"81",
          7975 => x"08",
          7976 => x"70",
          7977 => x"33",
          7978 => x"ff",
          7979 => x"84",
          7980 => x"77",
          7981 => x"06",
          7982 => x"bb",
          7983 => x"19",
          7984 => x"08",
          7985 => x"08",
          7986 => x"08",
          7987 => x"08",
          7988 => x"5b",
          7989 => x"ff",
          7990 => x"18",
          7991 => x"82",
          7992 => x"06",
          7993 => x"81",
          7994 => x"53",
          7995 => x"18",
          7996 => x"b7",
          7997 => x"33",
          7998 => x"83",
          7999 => x"06",
          8000 => x"84",
          8001 => x"76",
          8002 => x"81",
          8003 => x"38",
          8004 => x"84",
          8005 => x"57",
          8006 => x"81",
          8007 => x"ff",
          8008 => x"f4",
          8009 => x"0b",
          8010 => x"34",
          8011 => x"84",
          8012 => x"80",
          8013 => x"80",
          8014 => x"19",
          8015 => x"0b",
          8016 => x"80",
          8017 => x"19",
          8018 => x"0b",
          8019 => x"34",
          8020 => x"84",
          8021 => x"80",
          8022 => x"9e",
          8023 => x"e1",
          8024 => x"19",
          8025 => x"08",
          8026 => x"a0",
          8027 => x"88",
          8028 => x"84",
          8029 => x"74",
          8030 => x"75",
          8031 => x"34",
          8032 => x"5b",
          8033 => x"19",
          8034 => x"08",
          8035 => x"a4",
          8036 => x"88",
          8037 => x"84",
          8038 => x"7a",
          8039 => x"75",
          8040 => x"34",
          8041 => x"55",
          8042 => x"19",
          8043 => x"08",
          8044 => x"b4",
          8045 => x"81",
          8046 => x"79",
          8047 => x"33",
          8048 => x"3f",
          8049 => x"34",
          8050 => x"52",
          8051 => x"51",
          8052 => x"84",
          8053 => x"80",
          8054 => x"38",
          8055 => x"f3",
          8056 => x"60",
          8057 => x"56",
          8058 => x"27",
          8059 => x"17",
          8060 => x"8c",
          8061 => x"77",
          8062 => x"0c",
          8063 => x"04",
          8064 => x"56",
          8065 => x"2e",
          8066 => x"74",
          8067 => x"a5",
          8068 => x"2e",
          8069 => x"dd",
          8070 => x"2a",
          8071 => x"2a",
          8072 => x"05",
          8073 => x"5b",
          8074 => x"79",
          8075 => x"83",
          8076 => x"7b",
          8077 => x"81",
          8078 => x"38",
          8079 => x"53",
          8080 => x"81",
          8081 => x"f8",
          8082 => x"bb",
          8083 => x"2e",
          8084 => x"59",
          8085 => x"b4",
          8086 => x"ff",
          8087 => x"83",
          8088 => x"b8",
          8089 => x"1c",
          8090 => x"a8",
          8091 => x"53",
          8092 => x"b4",
          8093 => x"2e",
          8094 => x"0b",
          8095 => x"71",
          8096 => x"74",
          8097 => x"81",
          8098 => x"38",
          8099 => x"53",
          8100 => x"81",
          8101 => x"f8",
          8102 => x"bb",
          8103 => x"2e",
          8104 => x"59",
          8105 => x"b4",
          8106 => x"fe",
          8107 => x"83",
          8108 => x"b8",
          8109 => x"88",
          8110 => x"78",
          8111 => x"84",
          8112 => x"59",
          8113 => x"fe",
          8114 => x"9f",
          8115 => x"bb",
          8116 => x"3d",
          8117 => x"88",
          8118 => x"08",
          8119 => x"17",
          8120 => x"b5",
          8121 => x"83",
          8122 => x"5c",
          8123 => x"7b",
          8124 => x"06",
          8125 => x"81",
          8126 => x"b8",
          8127 => x"17",
          8128 => x"a8",
          8129 => x"84",
          8130 => x"85",
          8131 => x"81",
          8132 => x"18",
          8133 => x"df",
          8134 => x"83",
          8135 => x"05",
          8136 => x"11",
          8137 => x"71",
          8138 => x"84",
          8139 => x"57",
          8140 => x"0d",
          8141 => x"2e",
          8142 => x"fd",
          8143 => x"87",
          8144 => x"08",
          8145 => x"17",
          8146 => x"b5",
          8147 => x"83",
          8148 => x"5c",
          8149 => x"7b",
          8150 => x"06",
          8151 => x"81",
          8152 => x"b8",
          8153 => x"17",
          8154 => x"c0",
          8155 => x"84",
          8156 => x"85",
          8157 => x"81",
          8158 => x"18",
          8159 => x"f7",
          8160 => x"2b",
          8161 => x"77",
          8162 => x"83",
          8163 => x"12",
          8164 => x"2b",
          8165 => x"07",
          8166 => x"70",
          8167 => x"2b",
          8168 => x"80",
          8169 => x"80",
          8170 => x"bb",
          8171 => x"5c",
          8172 => x"56",
          8173 => x"04",
          8174 => x"17",
          8175 => x"17",
          8176 => x"18",
          8177 => x"f6",
          8178 => x"5a",
          8179 => x"08",
          8180 => x"81",
          8181 => x"38",
          8182 => x"08",
          8183 => x"b4",
          8184 => x"18",
          8185 => x"bb",
          8186 => x"5e",
          8187 => x"08",
          8188 => x"38",
          8189 => x"55",
          8190 => x"09",
          8191 => x"f7",
          8192 => x"b4",
          8193 => x"18",
          8194 => x"7b",
          8195 => x"33",
          8196 => x"3f",
          8197 => x"df",
          8198 => x"b4",
          8199 => x"b8",
          8200 => x"81",
          8201 => x"5c",
          8202 => x"84",
          8203 => x"7b",
          8204 => x"06",
          8205 => x"84",
          8206 => x"83",
          8207 => x"17",
          8208 => x"08",
          8209 => x"a0",
          8210 => x"8b",
          8211 => x"33",
          8212 => x"2e",
          8213 => x"84",
          8214 => x"5b",
          8215 => x"81",
          8216 => x"08",
          8217 => x"70",
          8218 => x"33",
          8219 => x"bb",
          8220 => x"84",
          8221 => x"7b",
          8222 => x"06",
          8223 => x"84",
          8224 => x"83",
          8225 => x"17",
          8226 => x"08",
          8227 => x"84",
          8228 => x"7d",
          8229 => x"27",
          8230 => x"82",
          8231 => x"74",
          8232 => x"81",
          8233 => x"38",
          8234 => x"17",
          8235 => x"08",
          8236 => x"52",
          8237 => x"51",
          8238 => x"7a",
          8239 => x"39",
          8240 => x"17",
          8241 => x"17",
          8242 => x"18",
          8243 => x"f4",
          8244 => x"5a",
          8245 => x"08",
          8246 => x"81",
          8247 => x"38",
          8248 => x"08",
          8249 => x"b4",
          8250 => x"18",
          8251 => x"bb",
          8252 => x"55",
          8253 => x"08",
          8254 => x"38",
          8255 => x"55",
          8256 => x"09",
          8257 => x"84",
          8258 => x"b4",
          8259 => x"18",
          8260 => x"7d",
          8261 => x"33",
          8262 => x"3f",
          8263 => x"ec",
          8264 => x"b4",
          8265 => x"18",
          8266 => x"7b",
          8267 => x"33",
          8268 => x"3f",
          8269 => x"81",
          8270 => x"bb",
          8271 => x"39",
          8272 => x"60",
          8273 => x"57",
          8274 => x"81",
          8275 => x"38",
          8276 => x"08",
          8277 => x"78",
          8278 => x"78",
          8279 => x"74",
          8280 => x"80",
          8281 => x"2e",
          8282 => x"77",
          8283 => x"0c",
          8284 => x"04",
          8285 => x"a8",
          8286 => x"58",
          8287 => x"1a",
          8288 => x"76",
          8289 => x"b6",
          8290 => x"33",
          8291 => x"7c",
          8292 => x"81",
          8293 => x"38",
          8294 => x"53",
          8295 => x"81",
          8296 => x"f2",
          8297 => x"bb",
          8298 => x"2e",
          8299 => x"58",
          8300 => x"b4",
          8301 => x"58",
          8302 => x"38",
          8303 => x"fe",
          8304 => x"7b",
          8305 => x"06",
          8306 => x"b8",
          8307 => x"88",
          8308 => x"b9",
          8309 => x"0b",
          8310 => x"77",
          8311 => x"0c",
          8312 => x"04",
          8313 => x"09",
          8314 => x"ff",
          8315 => x"2a",
          8316 => x"05",
          8317 => x"b4",
          8318 => x"5c",
          8319 => x"85",
          8320 => x"19",
          8321 => x"5d",
          8322 => x"09",
          8323 => x"bd",
          8324 => x"77",
          8325 => x"52",
          8326 => x"51",
          8327 => x"84",
          8328 => x"80",
          8329 => x"ff",
          8330 => x"77",
          8331 => x"79",
          8332 => x"b7",
          8333 => x"2b",
          8334 => x"79",
          8335 => x"83",
          8336 => x"98",
          8337 => x"06",
          8338 => x"06",
          8339 => x"5e",
          8340 => x"34",
          8341 => x"56",
          8342 => x"34",
          8343 => x"5a",
          8344 => x"34",
          8345 => x"5b",
          8346 => x"34",
          8347 => x"1a",
          8348 => x"39",
          8349 => x"16",
          8350 => x"a8",
          8351 => x"b4",
          8352 => x"59",
          8353 => x"2e",
          8354 => x"0b",
          8355 => x"71",
          8356 => x"74",
          8357 => x"81",
          8358 => x"38",
          8359 => x"53",
          8360 => x"81",
          8361 => x"f0",
          8362 => x"bb",
          8363 => x"2e",
          8364 => x"58",
          8365 => x"b4",
          8366 => x"58",
          8367 => x"38",
          8368 => x"06",
          8369 => x"81",
          8370 => x"06",
          8371 => x"7a",
          8372 => x"2e",
          8373 => x"84",
          8374 => x"06",
          8375 => x"06",
          8376 => x"5a",
          8377 => x"81",
          8378 => x"34",
          8379 => x"a8",
          8380 => x"56",
          8381 => x"1a",
          8382 => x"74",
          8383 => x"dd",
          8384 => x"74",
          8385 => x"70",
          8386 => x"33",
          8387 => x"9b",
          8388 => x"84",
          8389 => x"7f",
          8390 => x"06",
          8391 => x"84",
          8392 => x"83",
          8393 => x"19",
          8394 => x"1b",
          8395 => x"1b",
          8396 => x"84",
          8397 => x"56",
          8398 => x"27",
          8399 => x"19",
          8400 => x"82",
          8401 => x"38",
          8402 => x"53",
          8403 => x"19",
          8404 => x"d8",
          8405 => x"84",
          8406 => x"85",
          8407 => x"81",
          8408 => x"1a",
          8409 => x"83",
          8410 => x"ff",
          8411 => x"05",
          8412 => x"56",
          8413 => x"38",
          8414 => x"76",
          8415 => x"06",
          8416 => x"07",
          8417 => x"76",
          8418 => x"83",
          8419 => x"cb",
          8420 => x"76",
          8421 => x"70",
          8422 => x"33",
          8423 => x"8b",
          8424 => x"84",
          8425 => x"7c",
          8426 => x"06",
          8427 => x"84",
          8428 => x"83",
          8429 => x"19",
          8430 => x"1b",
          8431 => x"1b",
          8432 => x"84",
          8433 => x"40",
          8434 => x"27",
          8435 => x"82",
          8436 => x"74",
          8437 => x"81",
          8438 => x"38",
          8439 => x"1e",
          8440 => x"81",
          8441 => x"ee",
          8442 => x"5a",
          8443 => x"81",
          8444 => x"b8",
          8445 => x"81",
          8446 => x"57",
          8447 => x"81",
          8448 => x"84",
          8449 => x"09",
          8450 => x"ae",
          8451 => x"84",
          8452 => x"34",
          8453 => x"70",
          8454 => x"31",
          8455 => x"84",
          8456 => x"5f",
          8457 => x"74",
          8458 => x"f0",
          8459 => x"33",
          8460 => x"2e",
          8461 => x"fc",
          8462 => x"54",
          8463 => x"76",
          8464 => x"33",
          8465 => x"3f",
          8466 => x"d0",
          8467 => x"76",
          8468 => x"70",
          8469 => x"33",
          8470 => x"cf",
          8471 => x"84",
          8472 => x"7c",
          8473 => x"06",
          8474 => x"84",
          8475 => x"83",
          8476 => x"19",
          8477 => x"1b",
          8478 => x"1b",
          8479 => x"84",
          8480 => x"40",
          8481 => x"27",
          8482 => x"82",
          8483 => x"74",
          8484 => x"81",
          8485 => x"38",
          8486 => x"1e",
          8487 => x"81",
          8488 => x"ed",
          8489 => x"5a",
          8490 => x"81",
          8491 => x"53",
          8492 => x"19",
          8493 => x"f3",
          8494 => x"fd",
          8495 => x"76",
          8496 => x"06",
          8497 => x"83",
          8498 => x"59",
          8499 => x"b8",
          8500 => x"88",
          8501 => x"b9",
          8502 => x"fa",
          8503 => x"fd",
          8504 => x"76",
          8505 => x"fc",
          8506 => x"b8",
          8507 => x"33",
          8508 => x"8f",
          8509 => x"f0",
          8510 => x"42",
          8511 => x"58",
          8512 => x"7d",
          8513 => x"75",
          8514 => x"7d",
          8515 => x"79",
          8516 => x"7d",
          8517 => x"7a",
          8518 => x"fa",
          8519 => x"3d",
          8520 => x"71",
          8521 => x"5a",
          8522 => x"38",
          8523 => x"57",
          8524 => x"80",
          8525 => x"9c",
          8526 => x"80",
          8527 => x"19",
          8528 => x"54",
          8529 => x"80",
          8530 => x"7b",
          8531 => x"38",
          8532 => x"16",
          8533 => x"08",
          8534 => x"38",
          8535 => x"77",
          8536 => x"38",
          8537 => x"51",
          8538 => x"84",
          8539 => x"80",
          8540 => x"38",
          8541 => x"bb",
          8542 => x"2e",
          8543 => x"bb",
          8544 => x"70",
          8545 => x"07",
          8546 => x"7b",
          8547 => x"55",
          8548 => x"aa",
          8549 => x"2e",
          8550 => x"ff",
          8551 => x"55",
          8552 => x"84",
          8553 => x"0d",
          8554 => x"ff",
          8555 => x"bb",
          8556 => x"ca",
          8557 => x"79",
          8558 => x"3f",
          8559 => x"84",
          8560 => x"27",
          8561 => x"bb",
          8562 => x"84",
          8563 => x"ff",
          8564 => x"9c",
          8565 => x"bb",
          8566 => x"c4",
          8567 => x"fe",
          8568 => x"1b",
          8569 => x"08",
          8570 => x"38",
          8571 => x"52",
          8572 => x"eb",
          8573 => x"84",
          8574 => x"81",
          8575 => x"38",
          8576 => x"08",
          8577 => x"70",
          8578 => x"25",
          8579 => x"84",
          8580 => x"54",
          8581 => x"55",
          8582 => x"38",
          8583 => x"08",
          8584 => x"38",
          8585 => x"54",
          8586 => x"fe",
          8587 => x"9c",
          8588 => x"fe",
          8589 => x"70",
          8590 => x"96",
          8591 => x"2e",
          8592 => x"ff",
          8593 => x"78",
          8594 => x"3f",
          8595 => x"08",
          8596 => x"08",
          8597 => x"bb",
          8598 => x"80",
          8599 => x"55",
          8600 => x"38",
          8601 => x"38",
          8602 => x"0c",
          8603 => x"fe",
          8604 => x"08",
          8605 => x"78",
          8606 => x"ff",
          8607 => x"0c",
          8608 => x"81",
          8609 => x"84",
          8610 => x"55",
          8611 => x"84",
          8612 => x"0d",
          8613 => x"84",
          8614 => x"8c",
          8615 => x"84",
          8616 => x"58",
          8617 => x"73",
          8618 => x"b8",
          8619 => x"7a",
          8620 => x"f5",
          8621 => x"bb",
          8622 => x"ff",
          8623 => x"bb",
          8624 => x"bb",
          8625 => x"3d",
          8626 => x"56",
          8627 => x"ff",
          8628 => x"55",
          8629 => x"f8",
          8630 => x"7c",
          8631 => x"55",
          8632 => x"80",
          8633 => x"df",
          8634 => x"06",
          8635 => x"d7",
          8636 => x"19",
          8637 => x"08",
          8638 => x"df",
          8639 => x"56",
          8640 => x"80",
          8641 => x"85",
          8642 => x"0b",
          8643 => x"5a",
          8644 => x"27",
          8645 => x"17",
          8646 => x"0c",
          8647 => x"0c",
          8648 => x"53",
          8649 => x"80",
          8650 => x"73",
          8651 => x"98",
          8652 => x"83",
          8653 => x"b8",
          8654 => x"0c",
          8655 => x"84",
          8656 => x"8a",
          8657 => x"82",
          8658 => x"84",
          8659 => x"0d",
          8660 => x"08",
          8661 => x"2e",
          8662 => x"8a",
          8663 => x"89",
          8664 => x"73",
          8665 => x"38",
          8666 => x"53",
          8667 => x"14",
          8668 => x"59",
          8669 => x"8d",
          8670 => x"22",
          8671 => x"b0",
          8672 => x"5a",
          8673 => x"19",
          8674 => x"39",
          8675 => x"51",
          8676 => x"84",
          8677 => x"55",
          8678 => x"08",
          8679 => x"38",
          8680 => x"bb",
          8681 => x"ff",
          8682 => x"17",
          8683 => x"bb",
          8684 => x"27",
          8685 => x"73",
          8686 => x"73",
          8687 => x"38",
          8688 => x"81",
          8689 => x"84",
          8690 => x"0d",
          8691 => x"0d",
          8692 => x"90",
          8693 => x"05",
          8694 => x"f0",
          8695 => x"27",
          8696 => x"0b",
          8697 => x"98",
          8698 => x"84",
          8699 => x"2e",
          8700 => x"83",
          8701 => x"7a",
          8702 => x"15",
          8703 => x"57",
          8704 => x"38",
          8705 => x"88",
          8706 => x"55",
          8707 => x"81",
          8708 => x"98",
          8709 => x"90",
          8710 => x"1b",
          8711 => x"18",
          8712 => x"75",
          8713 => x"0c",
          8714 => x"04",
          8715 => x"0c",
          8716 => x"ff",
          8717 => x"2a",
          8718 => x"da",
          8719 => x"76",
          8720 => x"3f",
          8721 => x"08",
          8722 => x"81",
          8723 => x"84",
          8724 => x"38",
          8725 => x"bb",
          8726 => x"2e",
          8727 => x"19",
          8728 => x"84",
          8729 => x"91",
          8730 => x"2e",
          8731 => x"94",
          8732 => x"76",
          8733 => x"3f",
          8734 => x"08",
          8735 => x"84",
          8736 => x"80",
          8737 => x"38",
          8738 => x"bb",
          8739 => x"2e",
          8740 => x"81",
          8741 => x"84",
          8742 => x"ff",
          8743 => x"bb",
          8744 => x"1a",
          8745 => x"7d",
          8746 => x"fe",
          8747 => x"08",
          8748 => x"56",
          8749 => x"78",
          8750 => x"8a",
          8751 => x"71",
          8752 => x"08",
          8753 => x"7b",
          8754 => x"b8",
          8755 => x"80",
          8756 => x"80",
          8757 => x"05",
          8758 => x"15",
          8759 => x"38",
          8760 => x"19",
          8761 => x"75",
          8762 => x"38",
          8763 => x"1c",
          8764 => x"81",
          8765 => x"e4",
          8766 => x"bb",
          8767 => x"e7",
          8768 => x"56",
          8769 => x"98",
          8770 => x"0b",
          8771 => x"0c",
          8772 => x"04",
          8773 => x"19",
          8774 => x"19",
          8775 => x"1a",
          8776 => x"e4",
          8777 => x"bb",
          8778 => x"f3",
          8779 => x"84",
          8780 => x"34",
          8781 => x"a8",
          8782 => x"55",
          8783 => x"08",
          8784 => x"38",
          8785 => x"5c",
          8786 => x"09",
          8787 => x"db",
          8788 => x"b4",
          8789 => x"1a",
          8790 => x"75",
          8791 => x"33",
          8792 => x"3f",
          8793 => x"8a",
          8794 => x"74",
          8795 => x"06",
          8796 => x"2e",
          8797 => x"a7",
          8798 => x"18",
          8799 => x"9c",
          8800 => x"05",
          8801 => x"58",
          8802 => x"fd",
          8803 => x"19",
          8804 => x"29",
          8805 => x"05",
          8806 => x"5c",
          8807 => x"81",
          8808 => x"84",
          8809 => x"0d",
          8810 => x"0d",
          8811 => x"5c",
          8812 => x"5a",
          8813 => x"70",
          8814 => x"58",
          8815 => x"80",
          8816 => x"38",
          8817 => x"75",
          8818 => x"b4",
          8819 => x"2e",
          8820 => x"83",
          8821 => x"58",
          8822 => x"2e",
          8823 => x"81",
          8824 => x"54",
          8825 => x"19",
          8826 => x"33",
          8827 => x"3f",
          8828 => x"08",
          8829 => x"38",
          8830 => x"57",
          8831 => x"0c",
          8832 => x"82",
          8833 => x"1c",
          8834 => x"58",
          8835 => x"2e",
          8836 => x"8b",
          8837 => x"06",
          8838 => x"06",
          8839 => x"86",
          8840 => x"81",
          8841 => x"30",
          8842 => x"70",
          8843 => x"25",
          8844 => x"07",
          8845 => x"57",
          8846 => x"38",
          8847 => x"06",
          8848 => x"88",
          8849 => x"38",
          8850 => x"81",
          8851 => x"ff",
          8852 => x"7b",
          8853 => x"3f",
          8854 => x"08",
          8855 => x"84",
          8856 => x"38",
          8857 => x"56",
          8858 => x"38",
          8859 => x"84",
          8860 => x"0d",
          8861 => x"b4",
          8862 => x"7e",
          8863 => x"33",
          8864 => x"3f",
          8865 => x"bb",
          8866 => x"2e",
          8867 => x"fe",
          8868 => x"bb",
          8869 => x"1a",
          8870 => x"08",
          8871 => x"31",
          8872 => x"08",
          8873 => x"a0",
          8874 => x"fe",
          8875 => x"19",
          8876 => x"82",
          8877 => x"06",
          8878 => x"81",
          8879 => x"08",
          8880 => x"05",
          8881 => x"81",
          8882 => x"e0",
          8883 => x"57",
          8884 => x"79",
          8885 => x"81",
          8886 => x"38",
          8887 => x"81",
          8888 => x"80",
          8889 => x"8d",
          8890 => x"81",
          8891 => x"90",
          8892 => x"ac",
          8893 => x"5e",
          8894 => x"2e",
          8895 => x"ff",
          8896 => x"fe",
          8897 => x"56",
          8898 => x"09",
          8899 => x"be",
          8900 => x"84",
          8901 => x"98",
          8902 => x"84",
          8903 => x"94",
          8904 => x"77",
          8905 => x"39",
          8906 => x"57",
          8907 => x"09",
          8908 => x"38",
          8909 => x"9b",
          8910 => x"1a",
          8911 => x"2b",
          8912 => x"41",
          8913 => x"38",
          8914 => x"81",
          8915 => x"29",
          8916 => x"5a",
          8917 => x"5b",
          8918 => x"17",
          8919 => x"81",
          8920 => x"33",
          8921 => x"07",
          8922 => x"7a",
          8923 => x"c5",
          8924 => x"fe",
          8925 => x"38",
          8926 => x"05",
          8927 => x"75",
          8928 => x"1a",
          8929 => x"57",
          8930 => x"cc",
          8931 => x"70",
          8932 => x"06",
          8933 => x"80",
          8934 => x"79",
          8935 => x"fe",
          8936 => x"10",
          8937 => x"80",
          8938 => x"1d",
          8939 => x"06",
          8940 => x"9d",
          8941 => x"ff",
          8942 => x"38",
          8943 => x"fe",
          8944 => x"a8",
          8945 => x"8b",
          8946 => x"2a",
          8947 => x"29",
          8948 => x"81",
          8949 => x"40",
          8950 => x"81",
          8951 => x"19",
          8952 => x"76",
          8953 => x"7e",
          8954 => x"38",
          8955 => x"1d",
          8956 => x"bb",
          8957 => x"3d",
          8958 => x"3d",
          8959 => x"08",
          8960 => x"52",
          8961 => x"cf",
          8962 => x"84",
          8963 => x"bb",
          8964 => x"80",
          8965 => x"70",
          8966 => x"0b",
          8967 => x"b8",
          8968 => x"1c",
          8969 => x"58",
          8970 => x"76",
          8971 => x"38",
          8972 => x"78",
          8973 => x"78",
          8974 => x"06",
          8975 => x"81",
          8976 => x"b8",
          8977 => x"1b",
          8978 => x"e0",
          8979 => x"84",
          8980 => x"85",
          8981 => x"81",
          8982 => x"1c",
          8983 => x"76",
          8984 => x"9c",
          8985 => x"33",
          8986 => x"80",
          8987 => x"38",
          8988 => x"bf",
          8989 => x"ff",
          8990 => x"77",
          8991 => x"76",
          8992 => x"80",
          8993 => x"83",
          8994 => x"55",
          8995 => x"81",
          8996 => x"80",
          8997 => x"8f",
          8998 => x"38",
          8999 => x"78",
          9000 => x"8b",
          9001 => x"2a",
          9002 => x"29",
          9003 => x"81",
          9004 => x"57",
          9005 => x"81",
          9006 => x"19",
          9007 => x"76",
          9008 => x"7f",
          9009 => x"38",
          9010 => x"81",
          9011 => x"a7",
          9012 => x"a0",
          9013 => x"78",
          9014 => x"5a",
          9015 => x"81",
          9016 => x"71",
          9017 => x"1a",
          9018 => x"40",
          9019 => x"81",
          9020 => x"80",
          9021 => x"81",
          9022 => x"0b",
          9023 => x"80",
          9024 => x"f5",
          9025 => x"bb",
          9026 => x"84",
          9027 => x"80",
          9028 => x"38",
          9029 => x"84",
          9030 => x"0d",
          9031 => x"b4",
          9032 => x"7d",
          9033 => x"33",
          9034 => x"3f",
          9035 => x"bb",
          9036 => x"2e",
          9037 => x"fe",
          9038 => x"bb",
          9039 => x"1c",
          9040 => x"08",
          9041 => x"31",
          9042 => x"08",
          9043 => x"a0",
          9044 => x"fd",
          9045 => x"1b",
          9046 => x"82",
          9047 => x"06",
          9048 => x"81",
          9049 => x"08",
          9050 => x"05",
          9051 => x"81",
          9052 => x"db",
          9053 => x"57",
          9054 => x"77",
          9055 => x"39",
          9056 => x"70",
          9057 => x"06",
          9058 => x"fe",
          9059 => x"86",
          9060 => x"5a",
          9061 => x"93",
          9062 => x"33",
          9063 => x"06",
          9064 => x"08",
          9065 => x"0c",
          9066 => x"76",
          9067 => x"38",
          9068 => x"74",
          9069 => x"7b",
          9070 => x"3f",
          9071 => x"08",
          9072 => x"84",
          9073 => x"fc",
          9074 => x"c8",
          9075 => x"2e",
          9076 => x"81",
          9077 => x"0b",
          9078 => x"fe",
          9079 => x"19",
          9080 => x"77",
          9081 => x"06",
          9082 => x"1b",
          9083 => x"33",
          9084 => x"71",
          9085 => x"59",
          9086 => x"ff",
          9087 => x"33",
          9088 => x"8d",
          9089 => x"5b",
          9090 => x"59",
          9091 => x"84",
          9092 => x"05",
          9093 => x"71",
          9094 => x"2b",
          9095 => x"57",
          9096 => x"80",
          9097 => x"81",
          9098 => x"84",
          9099 => x"81",
          9100 => x"84",
          9101 => x"7a",
          9102 => x"70",
          9103 => x"81",
          9104 => x"81",
          9105 => x"75",
          9106 => x"08",
          9107 => x"06",
          9108 => x"76",
          9109 => x"58",
          9110 => x"ff",
          9111 => x"33",
          9112 => x"81",
          9113 => x"75",
          9114 => x"38",
          9115 => x"8d",
          9116 => x"60",
          9117 => x"41",
          9118 => x"b4",
          9119 => x"70",
          9120 => x"5e",
          9121 => x"39",
          9122 => x"bb",
          9123 => x"3d",
          9124 => x"83",
          9125 => x"ff",
          9126 => x"ff",
          9127 => x"39",
          9128 => x"68",
          9129 => x"ab",
          9130 => x"a0",
          9131 => x"5d",
          9132 => x"74",
          9133 => x"74",
          9134 => x"70",
          9135 => x"5d",
          9136 => x"8e",
          9137 => x"70",
          9138 => x"22",
          9139 => x"74",
          9140 => x"3d",
          9141 => x"40",
          9142 => x"58",
          9143 => x"70",
          9144 => x"33",
          9145 => x"05",
          9146 => x"15",
          9147 => x"38",
          9148 => x"05",
          9149 => x"06",
          9150 => x"80",
          9151 => x"38",
          9152 => x"ab",
          9153 => x"0b",
          9154 => x"5b",
          9155 => x"7b",
          9156 => x"7a",
          9157 => x"55",
          9158 => x"05",
          9159 => x"70",
          9160 => x"34",
          9161 => x"74",
          9162 => x"7b",
          9163 => x"38",
          9164 => x"56",
          9165 => x"2e",
          9166 => x"82",
          9167 => x"8f",
          9168 => x"06",
          9169 => x"76",
          9170 => x"83",
          9171 => x"72",
          9172 => x"06",
          9173 => x"57",
          9174 => x"87",
          9175 => x"a0",
          9176 => x"ff",
          9177 => x"80",
          9178 => x"78",
          9179 => x"ca",
          9180 => x"84",
          9181 => x"05",
          9182 => x"b0",
          9183 => x"55",
          9184 => x"84",
          9185 => x"55",
          9186 => x"ff",
          9187 => x"78",
          9188 => x"59",
          9189 => x"38",
          9190 => x"80",
          9191 => x"76",
          9192 => x"80",
          9193 => x"38",
          9194 => x"74",
          9195 => x"38",
          9196 => x"75",
          9197 => x"a2",
          9198 => x"70",
          9199 => x"74",
          9200 => x"81",
          9201 => x"81",
          9202 => x"55",
          9203 => x"8e",
          9204 => x"78",
          9205 => x"81",
          9206 => x"57",
          9207 => x"77",
          9208 => x"27",
          9209 => x"7d",
          9210 => x"3f",
          9211 => x"08",
          9212 => x"1b",
          9213 => x"7b",
          9214 => x"38",
          9215 => x"80",
          9216 => x"e7",
          9217 => x"84",
          9218 => x"bb",
          9219 => x"2e",
          9220 => x"82",
          9221 => x"80",
          9222 => x"ab",
          9223 => x"08",
          9224 => x"80",
          9225 => x"57",
          9226 => x"2a",
          9227 => x"81",
          9228 => x"2e",
          9229 => x"52",
          9230 => x"fe",
          9231 => x"84",
          9232 => x"1b",
          9233 => x"7d",
          9234 => x"3f",
          9235 => x"08",
          9236 => x"84",
          9237 => x"38",
          9238 => x"08",
          9239 => x"59",
          9240 => x"56",
          9241 => x"18",
          9242 => x"85",
          9243 => x"18",
          9244 => x"77",
          9245 => x"06",
          9246 => x"81",
          9247 => x"b8",
          9248 => x"18",
          9249 => x"a4",
          9250 => x"84",
          9251 => x"85",
          9252 => x"81",
          9253 => x"19",
          9254 => x"76",
          9255 => x"1e",
          9256 => x"56",
          9257 => x"e5",
          9258 => x"38",
          9259 => x"80",
          9260 => x"56",
          9261 => x"2e",
          9262 => x"81",
          9263 => x"7b",
          9264 => x"38",
          9265 => x"51",
          9266 => x"84",
          9267 => x"56",
          9268 => x"08",
          9269 => x"88",
          9270 => x"75",
          9271 => x"89",
          9272 => x"75",
          9273 => x"ff",
          9274 => x"81",
          9275 => x"1e",
          9276 => x"1c",
          9277 => x"af",
          9278 => x"33",
          9279 => x"7f",
          9280 => x"81",
          9281 => x"b8",
          9282 => x"1c",
          9283 => x"9c",
          9284 => x"84",
          9285 => x"85",
          9286 => x"81",
          9287 => x"1d",
          9288 => x"75",
          9289 => x"a0",
          9290 => x"08",
          9291 => x"76",
          9292 => x"58",
          9293 => x"55",
          9294 => x"8b",
          9295 => x"08",
          9296 => x"55",
          9297 => x"05",
          9298 => x"70",
          9299 => x"34",
          9300 => x"74",
          9301 => x"1e",
          9302 => x"33",
          9303 => x"5a",
          9304 => x"34",
          9305 => x"1d",
          9306 => x"75",
          9307 => x"0c",
          9308 => x"04",
          9309 => x"70",
          9310 => x"07",
          9311 => x"74",
          9312 => x"74",
          9313 => x"7d",
          9314 => x"3f",
          9315 => x"08",
          9316 => x"84",
          9317 => x"fd",
          9318 => x"bd",
          9319 => x"b4",
          9320 => x"7c",
          9321 => x"33",
          9322 => x"3f",
          9323 => x"08",
          9324 => x"81",
          9325 => x"38",
          9326 => x"08",
          9327 => x"b4",
          9328 => x"19",
          9329 => x"74",
          9330 => x"27",
          9331 => x"18",
          9332 => x"82",
          9333 => x"38",
          9334 => x"08",
          9335 => x"39",
          9336 => x"90",
          9337 => x"31",
          9338 => x"51",
          9339 => x"84",
          9340 => x"58",
          9341 => x"08",
          9342 => x"79",
          9343 => x"08",
          9344 => x"57",
          9345 => x"75",
          9346 => x"05",
          9347 => x"05",
          9348 => x"76",
          9349 => x"ff",
          9350 => x"59",
          9351 => x"e4",
          9352 => x"ff",
          9353 => x"43",
          9354 => x"08",
          9355 => x"b4",
          9356 => x"2e",
          9357 => x"1c",
          9358 => x"76",
          9359 => x"06",
          9360 => x"81",
          9361 => x"b8",
          9362 => x"1c",
          9363 => x"dc",
          9364 => x"84",
          9365 => x"85",
          9366 => x"81",
          9367 => x"1d",
          9368 => x"75",
          9369 => x"8c",
          9370 => x"1f",
          9371 => x"ff",
          9372 => x"5f",
          9373 => x"34",
          9374 => x"1c",
          9375 => x"1c",
          9376 => x"1c",
          9377 => x"1c",
          9378 => x"29",
          9379 => x"77",
          9380 => x"76",
          9381 => x"2e",
          9382 => x"10",
          9383 => x"81",
          9384 => x"56",
          9385 => x"18",
          9386 => x"55",
          9387 => x"81",
          9388 => x"76",
          9389 => x"75",
          9390 => x"85",
          9391 => x"ff",
          9392 => x"58",
          9393 => x"cb",
          9394 => x"ff",
          9395 => x"b3",
          9396 => x"1f",
          9397 => x"58",
          9398 => x"81",
          9399 => x"7b",
          9400 => x"83",
          9401 => x"52",
          9402 => x"e1",
          9403 => x"84",
          9404 => x"bb",
          9405 => x"f1",
          9406 => x"05",
          9407 => x"a9",
          9408 => x"39",
          9409 => x"1c",
          9410 => x"1c",
          9411 => x"1d",
          9412 => x"d0",
          9413 => x"56",
          9414 => x"08",
          9415 => x"84",
          9416 => x"83",
          9417 => x"1c",
          9418 => x"08",
          9419 => x"84",
          9420 => x"60",
          9421 => x"27",
          9422 => x"82",
          9423 => x"61",
          9424 => x"81",
          9425 => x"38",
          9426 => x"1c",
          9427 => x"08",
          9428 => x"52",
          9429 => x"51",
          9430 => x"77",
          9431 => x"39",
          9432 => x"08",
          9433 => x"43",
          9434 => x"e5",
          9435 => x"06",
          9436 => x"fb",
          9437 => x"70",
          9438 => x"80",
          9439 => x"38",
          9440 => x"7c",
          9441 => x"5d",
          9442 => x"81",
          9443 => x"08",
          9444 => x"81",
          9445 => x"cf",
          9446 => x"bb",
          9447 => x"2e",
          9448 => x"bc",
          9449 => x"84",
          9450 => x"34",
          9451 => x"a8",
          9452 => x"55",
          9453 => x"08",
          9454 => x"82",
          9455 => x"7e",
          9456 => x"38",
          9457 => x"08",
          9458 => x"39",
          9459 => x"41",
          9460 => x"2e",
          9461 => x"fc",
          9462 => x"1a",
          9463 => x"39",
          9464 => x"56",
          9465 => x"fc",
          9466 => x"fd",
          9467 => x"b4",
          9468 => x"1d",
          9469 => x"61",
          9470 => x"33",
          9471 => x"3f",
          9472 => x"81",
          9473 => x"08",
          9474 => x"05",
          9475 => x"81",
          9476 => x"ce",
          9477 => x"e3",
          9478 => x"0d",
          9479 => x"08",
          9480 => x"80",
          9481 => x"34",
          9482 => x"80",
          9483 => x"38",
          9484 => x"ff",
          9485 => x"38",
          9486 => x"60",
          9487 => x"70",
          9488 => x"5b",
          9489 => x"78",
          9490 => x"77",
          9491 => x"70",
          9492 => x"5b",
          9493 => x"82",
          9494 => x"d0",
          9495 => x"83",
          9496 => x"58",
          9497 => x"ff",
          9498 => x"38",
          9499 => x"76",
          9500 => x"5d",
          9501 => x"79",
          9502 => x"30",
          9503 => x"70",
          9504 => x"5a",
          9505 => x"18",
          9506 => x"80",
          9507 => x"34",
          9508 => x"1f",
          9509 => x"9c",
          9510 => x"70",
          9511 => x"58",
          9512 => x"a0",
          9513 => x"74",
          9514 => x"bc",
          9515 => x"32",
          9516 => x"72",
          9517 => x"55",
          9518 => x"8b",
          9519 => x"72",
          9520 => x"38",
          9521 => x"81",
          9522 => x"81",
          9523 => x"77",
          9524 => x"59",
          9525 => x"58",
          9526 => x"ff",
          9527 => x"18",
          9528 => x"80",
          9529 => x"34",
          9530 => x"53",
          9531 => x"77",
          9532 => x"bf",
          9533 => x"34",
          9534 => x"17",
          9535 => x"80",
          9536 => x"34",
          9537 => x"8c",
          9538 => x"53",
          9539 => x"73",
          9540 => x"9c",
          9541 => x"8b",
          9542 => x"1e",
          9543 => x"08",
          9544 => x"11",
          9545 => x"33",
          9546 => x"71",
          9547 => x"81",
          9548 => x"72",
          9549 => x"75",
          9550 => x"64",
          9551 => x"16",
          9552 => x"33",
          9553 => x"07",
          9554 => x"40",
          9555 => x"55",
          9556 => x"23",
          9557 => x"98",
          9558 => x"88",
          9559 => x"54",
          9560 => x"23",
          9561 => x"04",
          9562 => x"fe",
          9563 => x"1d",
          9564 => x"ff",
          9565 => x"5b",
          9566 => x"52",
          9567 => x"74",
          9568 => x"90",
          9569 => x"bb",
          9570 => x"ff",
          9571 => x"81",
          9572 => x"ad",
          9573 => x"27",
          9574 => x"74",
          9575 => x"73",
          9576 => x"97",
          9577 => x"78",
          9578 => x"0b",
          9579 => x"56",
          9580 => x"75",
          9581 => x"5c",
          9582 => x"fd",
          9583 => x"ba",
          9584 => x"76",
          9585 => x"07",
          9586 => x"80",
          9587 => x"55",
          9588 => x"f9",
          9589 => x"34",
          9590 => x"58",
          9591 => x"1f",
          9592 => x"cd",
          9593 => x"89",
          9594 => x"57",
          9595 => x"2e",
          9596 => x"7c",
          9597 => x"57",
          9598 => x"14",
          9599 => x"11",
          9600 => x"99",
          9601 => x"9c",
          9602 => x"11",
          9603 => x"88",
          9604 => x"38",
          9605 => x"53",
          9606 => x"5e",
          9607 => x"8a",
          9608 => x"70",
          9609 => x"06",
          9610 => x"78",
          9611 => x"5a",
          9612 => x"81",
          9613 => x"71",
          9614 => x"5e",
          9615 => x"56",
          9616 => x"38",
          9617 => x"72",
          9618 => x"cc",
          9619 => x"30",
          9620 => x"70",
          9621 => x"53",
          9622 => x"fc",
          9623 => x"3d",
          9624 => x"08",
          9625 => x"5c",
          9626 => x"33",
          9627 => x"74",
          9628 => x"38",
          9629 => x"80",
          9630 => x"df",
          9631 => x"2e",
          9632 => x"98",
          9633 => x"1d",
          9634 => x"96",
          9635 => x"41",
          9636 => x"75",
          9637 => x"38",
          9638 => x"16",
          9639 => x"57",
          9640 => x"81",
          9641 => x"55",
          9642 => x"df",
          9643 => x"0c",
          9644 => x"81",
          9645 => x"ff",
          9646 => x"8b",
          9647 => x"18",
          9648 => x"23",
          9649 => x"73",
          9650 => x"06",
          9651 => x"70",
          9652 => x"27",
          9653 => x"07",
          9654 => x"55",
          9655 => x"38",
          9656 => x"2e",
          9657 => x"74",
          9658 => x"b2",
          9659 => x"a0",
          9660 => x"a0",
          9661 => x"ff",
          9662 => x"56",
          9663 => x"81",
          9664 => x"75",
          9665 => x"81",
          9666 => x"70",
          9667 => x"56",
          9668 => x"ee",
          9669 => x"ff",
          9670 => x"81",
          9671 => x"81",
          9672 => x"fd",
          9673 => x"18",
          9674 => x"23",
          9675 => x"70",
          9676 => x"52",
          9677 => x"57",
          9678 => x"fe",
          9679 => x"cb",
          9680 => x"80",
          9681 => x"30",
          9682 => x"73",
          9683 => x"58",
          9684 => x"2e",
          9685 => x"14",
          9686 => x"80",
          9687 => x"55",
          9688 => x"dd",
          9689 => x"dc",
          9690 => x"70",
          9691 => x"07",
          9692 => x"72",
          9693 => x"88",
          9694 => x"33",
          9695 => x"3d",
          9696 => x"74",
          9697 => x"90",
          9698 => x"83",
          9699 => x"51",
          9700 => x"3f",
          9701 => x"08",
          9702 => x"06",
          9703 => x"8d",
          9704 => x"73",
          9705 => x"0c",
          9706 => x"04",
          9707 => x"33",
          9708 => x"06",
          9709 => x"80",
          9710 => x"38",
          9711 => x"80",
          9712 => x"34",
          9713 => x"51",
          9714 => x"84",
          9715 => x"84",
          9716 => x"93",
          9717 => x"81",
          9718 => x"32",
          9719 => x"80",
          9720 => x"41",
          9721 => x"7d",
          9722 => x"38",
          9723 => x"80",
          9724 => x"55",
          9725 => x"af",
          9726 => x"72",
          9727 => x"70",
          9728 => x"25",
          9729 => x"54",
          9730 => x"38",
          9731 => x"9f",
          9732 => x"2b",
          9733 => x"2e",
          9734 => x"76",
          9735 => x"d1",
          9736 => x"59",
          9737 => x"a7",
          9738 => x"78",
          9739 => x"70",
          9740 => x"32",
          9741 => x"9f",
          9742 => x"56",
          9743 => x"7c",
          9744 => x"38",
          9745 => x"ff",
          9746 => x"dd",
          9747 => x"77",
          9748 => x"76",
          9749 => x"2e",
          9750 => x"80",
          9751 => x"83",
          9752 => x"72",
          9753 => x"56",
          9754 => x"82",
          9755 => x"83",
          9756 => x"53",
          9757 => x"82",
          9758 => x"80",
          9759 => x"77",
          9760 => x"70",
          9761 => x"78",
          9762 => x"38",
          9763 => x"fe",
          9764 => x"17",
          9765 => x"2e",
          9766 => x"14",
          9767 => x"54",
          9768 => x"09",
          9769 => x"38",
          9770 => x"1d",
          9771 => x"74",
          9772 => x"56",
          9773 => x"53",
          9774 => x"72",
          9775 => x"88",
          9776 => x"22",
          9777 => x"57",
          9778 => x"80",
          9779 => x"38",
          9780 => x"83",
          9781 => x"ae",
          9782 => x"70",
          9783 => x"5a",
          9784 => x"2e",
          9785 => x"72",
          9786 => x"72",
          9787 => x"26",
          9788 => x"59",
          9789 => x"70",
          9790 => x"07",
          9791 => x"7c",
          9792 => x"54",
          9793 => x"2e",
          9794 => x"7c",
          9795 => x"83",
          9796 => x"2e",
          9797 => x"83",
          9798 => x"77",
          9799 => x"76",
          9800 => x"8b",
          9801 => x"81",
          9802 => x"18",
          9803 => x"77",
          9804 => x"81",
          9805 => x"53",
          9806 => x"38",
          9807 => x"57",
          9808 => x"2e",
          9809 => x"7c",
          9810 => x"e3",
          9811 => x"06",
          9812 => x"2e",
          9813 => x"7d",
          9814 => x"74",
          9815 => x"e3",
          9816 => x"2a",
          9817 => x"75",
          9818 => x"81",
          9819 => x"80",
          9820 => x"79",
          9821 => x"7d",
          9822 => x"06",
          9823 => x"2e",
          9824 => x"88",
          9825 => x"ab",
          9826 => x"51",
          9827 => x"84",
          9828 => x"ab",
          9829 => x"54",
          9830 => x"08",
          9831 => x"ac",
          9832 => x"84",
          9833 => x"09",
          9834 => x"f7",
          9835 => x"2a",
          9836 => x"79",
          9837 => x"f0",
          9838 => x"2a",
          9839 => x"78",
          9840 => x"7b",
          9841 => x"56",
          9842 => x"16",
          9843 => x"57",
          9844 => x"81",
          9845 => x"79",
          9846 => x"40",
          9847 => x"7c",
          9848 => x"38",
          9849 => x"fd",
          9850 => x"83",
          9851 => x"8a",
          9852 => x"22",
          9853 => x"2e",
          9854 => x"fc",
          9855 => x"22",
          9856 => x"2e",
          9857 => x"fc",
          9858 => x"10",
          9859 => x"7b",
          9860 => x"a0",
          9861 => x"ae",
          9862 => x"26",
          9863 => x"54",
          9864 => x"81",
          9865 => x"81",
          9866 => x"73",
          9867 => x"79",
          9868 => x"77",
          9869 => x"7b",
          9870 => x"3f",
          9871 => x"08",
          9872 => x"56",
          9873 => x"84",
          9874 => x"38",
          9875 => x"81",
          9876 => x"fa",
          9877 => x"1c",
          9878 => x"2a",
          9879 => x"5d",
          9880 => x"83",
          9881 => x"1c",
          9882 => x"06",
          9883 => x"d3",
          9884 => x"d2",
          9885 => x"88",
          9886 => x"33",
          9887 => x"54",
          9888 => x"82",
          9889 => x"88",
          9890 => x"08",
          9891 => x"fe",
          9892 => x"22",
          9893 => x"2e",
          9894 => x"76",
          9895 => x"fb",
          9896 => x"ab",
          9897 => x"07",
          9898 => x"5a",
          9899 => x"7d",
          9900 => x"fc",
          9901 => x"06",
          9902 => x"8c",
          9903 => x"06",
          9904 => x"79",
          9905 => x"fd",
          9906 => x"0b",
          9907 => x"7c",
          9908 => x"81",
          9909 => x"38",
          9910 => x"80",
          9911 => x"34",
          9912 => x"bb",
          9913 => x"3d",
          9914 => x"80",
          9915 => x"38",
          9916 => x"27",
          9917 => x"ff",
          9918 => x"7b",
          9919 => x"38",
          9920 => x"7d",
          9921 => x"5c",
          9922 => x"39",
          9923 => x"5a",
          9924 => x"74",
          9925 => x"bd",
          9926 => x"84",
          9927 => x"ff",
          9928 => x"2a",
          9929 => x"55",
          9930 => x"c4",
          9931 => x"ff",
          9932 => x"94",
          9933 => x"54",
          9934 => x"26",
          9935 => x"74",
          9936 => x"85",
          9937 => x"ac",
          9938 => x"ac",
          9939 => x"ff",
          9940 => x"59",
          9941 => x"80",
          9942 => x"75",
          9943 => x"81",
          9944 => x"70",
          9945 => x"56",
          9946 => x"ee",
          9947 => x"ff",
          9948 => x"80",
          9949 => x"bf",
          9950 => x"99",
          9951 => x"7d",
          9952 => x"81",
          9953 => x"53",
          9954 => x"59",
          9955 => x"93",
          9956 => x"07",
          9957 => x"06",
          9958 => x"83",
          9959 => x"58",
          9960 => x"7b",
          9961 => x"59",
          9962 => x"81",
          9963 => x"16",
          9964 => x"39",
          9965 => x"b3",
          9966 => x"ac",
          9967 => x"ff",
          9968 => x"78",
          9969 => x"ae",
          9970 => x"7a",
          9971 => x"1d",
          9972 => x"5b",
          9973 => x"34",
          9974 => x"d2",
          9975 => x"14",
          9976 => x"15",
          9977 => x"2b",
          9978 => x"07",
          9979 => x"1f",
          9980 => x"fd",
          9981 => x"1b",
          9982 => x"88",
          9983 => x"72",
          9984 => x"1b",
          9985 => x"05",
          9986 => x"79",
          9987 => x"5b",
          9988 => x"79",
          9989 => x"1d",
          9990 => x"76",
          9991 => x"09",
          9992 => x"a3",
          9993 => x"39",
          9994 => x"81",
          9995 => x"f6",
          9996 => x"0b",
          9997 => x"0c",
          9998 => x"04",
          9999 => x"67",
         10000 => x"05",
         10001 => x"33",
         10002 => x"80",
         10003 => x"7e",
         10004 => x"5b",
         10005 => x"2e",
         10006 => x"79",
         10007 => x"5b",
         10008 => x"26",
         10009 => x"ba",
         10010 => x"38",
         10011 => x"75",
         10012 => x"c7",
         10013 => x"e0",
         10014 => x"76",
         10015 => x"38",
         10016 => x"84",
         10017 => x"70",
         10018 => x"8c",
         10019 => x"2e",
         10020 => x"76",
         10021 => x"81",
         10022 => x"33",
         10023 => x"80",
         10024 => x"81",
         10025 => x"ff",
         10026 => x"84",
         10027 => x"81",
         10028 => x"81",
         10029 => x"7c",
         10030 => x"96",
         10031 => x"34",
         10032 => x"84",
         10033 => x"33",
         10034 => x"81",
         10035 => x"33",
         10036 => x"a4",
         10037 => x"84",
         10038 => x"06",
         10039 => x"41",
         10040 => x"7f",
         10041 => x"78",
         10042 => x"38",
         10043 => x"81",
         10044 => x"58",
         10045 => x"38",
         10046 => x"83",
         10047 => x"0b",
         10048 => x"7a",
         10049 => x"81",
         10050 => x"b8",
         10051 => x"81",
         10052 => x"58",
         10053 => x"3f",
         10054 => x"08",
         10055 => x"38",
         10056 => x"59",
         10057 => x"0c",
         10058 => x"99",
         10059 => x"17",
         10060 => x"18",
         10061 => x"2b",
         10062 => x"83",
         10063 => x"d4",
         10064 => x"a5",
         10065 => x"26",
         10066 => x"ba",
         10067 => x"42",
         10068 => x"38",
         10069 => x"84",
         10070 => x"38",
         10071 => x"81",
         10072 => x"38",
         10073 => x"33",
         10074 => x"33",
         10075 => x"07",
         10076 => x"84",
         10077 => x"81",
         10078 => x"38",
         10079 => x"33",
         10080 => x"33",
         10081 => x"07",
         10082 => x"a4",
         10083 => x"17",
         10084 => x"82",
         10085 => x"90",
         10086 => x"2b",
         10087 => x"33",
         10088 => x"88",
         10089 => x"71",
         10090 => x"45",
         10091 => x"56",
         10092 => x"0c",
         10093 => x"33",
         10094 => x"80",
         10095 => x"ff",
         10096 => x"ff",
         10097 => x"59",
         10098 => x"81",
         10099 => x"38",
         10100 => x"06",
         10101 => x"80",
         10102 => x"5a",
         10103 => x"8a",
         10104 => x"59",
         10105 => x"87",
         10106 => x"18",
         10107 => x"61",
         10108 => x"80",
         10109 => x"80",
         10110 => x"71",
         10111 => x"56",
         10112 => x"18",
         10113 => x"8f",
         10114 => x"8d",
         10115 => x"98",
         10116 => x"17",
         10117 => x"18",
         10118 => x"2b",
         10119 => x"74",
         10120 => x"d8",
         10121 => x"33",
         10122 => x"71",
         10123 => x"88",
         10124 => x"14",
         10125 => x"07",
         10126 => x"33",
         10127 => x"44",
         10128 => x"42",
         10129 => x"17",
         10130 => x"18",
         10131 => x"2b",
         10132 => x"8d",
         10133 => x"2e",
         10134 => x"7d",
         10135 => x"2a",
         10136 => x"75",
         10137 => x"38",
         10138 => x"7a",
         10139 => x"ec",
         10140 => x"bb",
         10141 => x"84",
         10142 => x"80",
         10143 => x"38",
         10144 => x"08",
         10145 => x"ff",
         10146 => x"38",
         10147 => x"83",
         10148 => x"83",
         10149 => x"75",
         10150 => x"85",
         10151 => x"5d",
         10152 => x"9c",
         10153 => x"a4",
         10154 => x"1d",
         10155 => x"0c",
         10156 => x"1a",
         10157 => x"7c",
         10158 => x"87",
         10159 => x"22",
         10160 => x"7b",
         10161 => x"e0",
         10162 => x"ac",
         10163 => x"19",
         10164 => x"2e",
         10165 => x"10",
         10166 => x"2a",
         10167 => x"05",
         10168 => x"ff",
         10169 => x"59",
         10170 => x"a0",
         10171 => x"b8",
         10172 => x"94",
         10173 => x"0b",
         10174 => x"ff",
         10175 => x"18",
         10176 => x"2e",
         10177 => x"7c",
         10178 => x"e2",
         10179 => x"05",
         10180 => x"e2",
         10181 => x"86",
         10182 => x"e2",
         10183 => x"18",
         10184 => x"98",
         10185 => x"58",
         10186 => x"84",
         10187 => x"0d",
         10188 => x"84",
         10189 => x"97",
         10190 => x"76",
         10191 => x"70",
         10192 => x"57",
         10193 => x"89",
         10194 => x"82",
         10195 => x"ff",
         10196 => x"5d",
         10197 => x"2e",
         10198 => x"80",
         10199 => x"e6",
         10200 => x"5c",
         10201 => x"5a",
         10202 => x"81",
         10203 => x"79",
         10204 => x"5b",
         10205 => x"12",
         10206 => x"77",
         10207 => x"38",
         10208 => x"81",
         10209 => x"55",
         10210 => x"58",
         10211 => x"89",
         10212 => x"70",
         10213 => x"58",
         10214 => x"70",
         10215 => x"55",
         10216 => x"09",
         10217 => x"38",
         10218 => x"38",
         10219 => x"70",
         10220 => x"07",
         10221 => x"07",
         10222 => x"7a",
         10223 => x"98",
         10224 => x"84",
         10225 => x"83",
         10226 => x"98",
         10227 => x"f9",
         10228 => x"80",
         10229 => x"38",
         10230 => x"81",
         10231 => x"58",
         10232 => x"38",
         10233 => x"c0",
         10234 => x"33",
         10235 => x"81",
         10236 => x"81",
         10237 => x"81",
         10238 => x"eb",
         10239 => x"70",
         10240 => x"07",
         10241 => x"77",
         10242 => x"75",
         10243 => x"83",
         10244 => x"3d",
         10245 => x"83",
         10246 => x"16",
         10247 => x"5b",
         10248 => x"a5",
         10249 => x"16",
         10250 => x"17",
         10251 => x"2b",
         10252 => x"07",
         10253 => x"33",
         10254 => x"88",
         10255 => x"1b",
         10256 => x"52",
         10257 => x"40",
         10258 => x"70",
         10259 => x"0c",
         10260 => x"17",
         10261 => x"80",
         10262 => x"38",
         10263 => x"1d",
         10264 => x"70",
         10265 => x"71",
         10266 => x"71",
         10267 => x"f0",
         10268 => x"1c",
         10269 => x"43",
         10270 => x"08",
         10271 => x"7a",
         10272 => x"fb",
         10273 => x"83",
         10274 => x"0b",
         10275 => x"7a",
         10276 => x"7a",
         10277 => x"38",
         10278 => x"53",
         10279 => x"81",
         10280 => x"ff",
         10281 => x"84",
         10282 => x"76",
         10283 => x"ff",
         10284 => x"74",
         10285 => x"84",
         10286 => x"38",
         10287 => x"7f",
         10288 => x"2b",
         10289 => x"83",
         10290 => x"d4",
         10291 => x"81",
         10292 => x"80",
         10293 => x"33",
         10294 => x"81",
         10295 => x"b7",
         10296 => x"eb",
         10297 => x"70",
         10298 => x"07",
         10299 => x"7f",
         10300 => x"81",
         10301 => x"38",
         10302 => x"81",
         10303 => x"80",
         10304 => x"f9",
         10305 => x"58",
         10306 => x"09",
         10307 => x"38",
         10308 => x"76",
         10309 => x"38",
         10310 => x"f8",
         10311 => x"1a",
         10312 => x"5a",
         10313 => x"fe",
         10314 => x"a8",
         10315 => x"80",
         10316 => x"e6",
         10317 => x"58",
         10318 => x"05",
         10319 => x"70",
         10320 => x"33",
         10321 => x"ff",
         10322 => x"56",
         10323 => x"2e",
         10324 => x"75",
         10325 => x"38",
         10326 => x"8a",
         10327 => x"b8",
         10328 => x"7b",
         10329 => x"5d",
         10330 => x"81",
         10331 => x"71",
         10332 => x"1b",
         10333 => x"40",
         10334 => x"85",
         10335 => x"80",
         10336 => x"82",
         10337 => x"39",
         10338 => x"fa",
         10339 => x"84",
         10340 => x"97",
         10341 => x"75",
         10342 => x"2e",
         10343 => x"85",
         10344 => x"18",
         10345 => x"40",
         10346 => x"b7",
         10347 => x"84",
         10348 => x"97",
         10349 => x"83",
         10350 => x"18",
         10351 => x"5c",
         10352 => x"70",
         10353 => x"33",
         10354 => x"05",
         10355 => x"71",
         10356 => x"5b",
         10357 => x"77",
         10358 => x"d1",
         10359 => x"2e",
         10360 => x"0b",
         10361 => x"83",
         10362 => x"5a",
         10363 => x"81",
         10364 => x"7a",
         10365 => x"5c",
         10366 => x"31",
         10367 => x"58",
         10368 => x"80",
         10369 => x"38",
         10370 => x"e1",
         10371 => x"77",
         10372 => x"59",
         10373 => x"81",
         10374 => x"39",
         10375 => x"33",
         10376 => x"33",
         10377 => x"07",
         10378 => x"81",
         10379 => x"06",
         10380 => x"81",
         10381 => x"5a",
         10382 => x"78",
         10383 => x"83",
         10384 => x"7a",
         10385 => x"81",
         10386 => x"38",
         10387 => x"53",
         10388 => x"81",
         10389 => x"ff",
         10390 => x"84",
         10391 => x"80",
         10392 => x"ff",
         10393 => x"77",
         10394 => x"79",
         10395 => x"79",
         10396 => x"84",
         10397 => x"84",
         10398 => x"71",
         10399 => x"57",
         10400 => x"d4",
         10401 => x"81",
         10402 => x"38",
         10403 => x"11",
         10404 => x"33",
         10405 => x"71",
         10406 => x"81",
         10407 => x"72",
         10408 => x"75",
         10409 => x"5e",
         10410 => x"42",
         10411 => x"84",
         10412 => x"d2",
         10413 => x"06",
         10414 => x"84",
         10415 => x"11",
         10416 => x"33",
         10417 => x"71",
         10418 => x"81",
         10419 => x"72",
         10420 => x"75",
         10421 => x"47",
         10422 => x"5c",
         10423 => x"86",
         10424 => x"f2",
         10425 => x"06",
         10426 => x"84",
         10427 => x"11",
         10428 => x"33",
         10429 => x"71",
         10430 => x"81",
         10431 => x"72",
         10432 => x"75",
         10433 => x"94",
         10434 => x"84",
         10435 => x"11",
         10436 => x"33",
         10437 => x"71",
         10438 => x"81",
         10439 => x"72",
         10440 => x"75",
         10441 => x"62",
         10442 => x"59",
         10443 => x"5c",
         10444 => x"5b",
         10445 => x"77",
         10446 => x"dc",
         10447 => x"5d",
         10448 => x"dc",
         10449 => x"18",
         10450 => x"e4",
         10451 => x"0c",
         10452 => x"18",
         10453 => x"39",
         10454 => x"f8",
         10455 => x"7a",
         10456 => x"f2",
         10457 => x"54",
         10458 => x"53",
         10459 => x"53",
         10460 => x"52",
         10461 => x"b3",
         10462 => x"84",
         10463 => x"09",
         10464 => x"a4",
         10465 => x"84",
         10466 => x"34",
         10467 => x"a8",
         10468 => x"40",
         10469 => x"08",
         10470 => x"82",
         10471 => x"60",
         10472 => x"8d",
         10473 => x"84",
         10474 => x"a0",
         10475 => x"74",
         10476 => x"91",
         10477 => x"81",
         10478 => x"e6",
         10479 => x"58",
         10480 => x"80",
         10481 => x"80",
         10482 => x"71",
         10483 => x"5f",
         10484 => x"7d",
         10485 => x"88",
         10486 => x"61",
         10487 => x"80",
         10488 => x"11",
         10489 => x"33",
         10490 => x"71",
         10491 => x"81",
         10492 => x"72",
         10493 => x"75",
         10494 => x"ac",
         10495 => x"7d",
         10496 => x"43",
         10497 => x"40",
         10498 => x"75",
         10499 => x"2e",
         10500 => x"82",
         10501 => x"39",
         10502 => x"f2",
         10503 => x"3d",
         10504 => x"83",
         10505 => x"39",
         10506 => x"f5",
         10507 => x"bf",
         10508 => x"b4",
         10509 => x"18",
         10510 => x"78",
         10511 => x"33",
         10512 => x"e7",
         10513 => x"39",
         10514 => x"02",
         10515 => x"33",
         10516 => x"93",
         10517 => x"5d",
         10518 => x"40",
         10519 => x"80",
         10520 => x"70",
         10521 => x"33",
         10522 => x"55",
         10523 => x"2e",
         10524 => x"73",
         10525 => x"ba",
         10526 => x"38",
         10527 => x"33",
         10528 => x"24",
         10529 => x"73",
         10530 => x"e2",
         10531 => x"08",
         10532 => x"80",
         10533 => x"80",
         10534 => x"54",
         10535 => x"86",
         10536 => x"34",
         10537 => x"75",
         10538 => x"7c",
         10539 => x"38",
         10540 => x"3d",
         10541 => x"05",
         10542 => x"3f",
         10543 => x"08",
         10544 => x"bb",
         10545 => x"3d",
         10546 => x"0b",
         10547 => x"0c",
         10548 => x"04",
         10549 => x"11",
         10550 => x"06",
         10551 => x"73",
         10552 => x"38",
         10553 => x"81",
         10554 => x"05",
         10555 => x"79",
         10556 => x"38",
         10557 => x"83",
         10558 => x"5f",
         10559 => x"7e",
         10560 => x"70",
         10561 => x"33",
         10562 => x"05",
         10563 => x"9f",
         10564 => x"55",
         10565 => x"89",
         10566 => x"70",
         10567 => x"56",
         10568 => x"16",
         10569 => x"26",
         10570 => x"16",
         10571 => x"06",
         10572 => x"30",
         10573 => x"58",
         10574 => x"2e",
         10575 => x"85",
         10576 => x"be",
         10577 => x"32",
         10578 => x"72",
         10579 => x"79",
         10580 => x"54",
         10581 => x"92",
         10582 => x"84",
         10583 => x"83",
         10584 => x"99",
         10585 => x"fe",
         10586 => x"83",
         10587 => x"7a",
         10588 => x"54",
         10589 => x"e6",
         10590 => x"02",
         10591 => x"fb",
         10592 => x"5a",
         10593 => x"80",
         10594 => x"74",
         10595 => x"54",
         10596 => x"05",
         10597 => x"84",
         10598 => x"ed",
         10599 => x"bb",
         10600 => x"84",
         10601 => x"80",
         10602 => x"80",
         10603 => x"56",
         10604 => x"84",
         10605 => x"0d",
         10606 => x"6d",
         10607 => x"70",
         10608 => x"9a",
         10609 => x"84",
         10610 => x"bb",
         10611 => x"2e",
         10612 => x"78",
         10613 => x"7c",
         10614 => x"ca",
         10615 => x"2e",
         10616 => x"76",
         10617 => x"f2",
         10618 => x"07",
         10619 => x"bb",
         10620 => x"2a",
         10621 => x"77",
         10622 => x"d1",
         10623 => x"11",
         10624 => x"33",
         10625 => x"07",
         10626 => x"42",
         10627 => x"56",
         10628 => x"86",
         10629 => x"0b",
         10630 => x"80",
         10631 => x"34",
         10632 => x"17",
         10633 => x"0b",
         10634 => x"66",
         10635 => x"8b",
         10636 => x"67",
         10637 => x"0b",
         10638 => x"80",
         10639 => x"34",
         10640 => x"7c",
         10641 => x"d7",
         10642 => x"80",
         10643 => x"34",
         10644 => x"19",
         10645 => x"9e",
         10646 => x"0b",
         10647 => x"7e",
         10648 => x"83",
         10649 => x"80",
         10650 => x"38",
         10651 => x"08",
         10652 => x"59",
         10653 => x"81",
         10654 => x"38",
         10655 => x"7b",
         10656 => x"38",
         10657 => x"7a",
         10658 => x"39",
         10659 => x"05",
         10660 => x"2b",
         10661 => x"80",
         10662 => x"38",
         10663 => x"06",
         10664 => x"fe",
         10665 => x"fe",
         10666 => x"80",
         10667 => x"70",
         10668 => x"06",
         10669 => x"82",
         10670 => x"81",
         10671 => x"5d",
         10672 => x"89",
         10673 => x"06",
         10674 => x"95",
         10675 => x"2a",
         10676 => x"75",
         10677 => x"38",
         10678 => x"07",
         10679 => x"11",
         10680 => x"0c",
         10681 => x"0c",
         10682 => x"33",
         10683 => x"71",
         10684 => x"73",
         10685 => x"40",
         10686 => x"83",
         10687 => x"38",
         10688 => x"0c",
         10689 => x"11",
         10690 => x"33",
         10691 => x"71",
         10692 => x"81",
         10693 => x"72",
         10694 => x"75",
         10695 => x"60",
         10696 => x"43",
         10697 => x"41",
         10698 => x"56",
         10699 => x"84",
         10700 => x"90",
         10701 => x"0b",
         10702 => x"80",
         10703 => x"0c",
         10704 => x"1b",
         10705 => x"5c",
         10706 => x"57",
         10707 => x"70",
         10708 => x"34",
         10709 => x"74",
         10710 => x"85",
         10711 => x"59",
         10712 => x"fc",
         10713 => x"1a",
         10714 => x"80",
         10715 => x"38",
         10716 => x"0c",
         10717 => x"70",
         10718 => x"1c",
         10719 => x"5a",
         10720 => x"30",
         10721 => x"80",
         10722 => x"78",
         10723 => x"e7",
         10724 => x"76",
         10725 => x"7c",
         10726 => x"db",
         10727 => x"79",
         10728 => x"bb",
         10729 => x"84",
         10730 => x"bb",
         10731 => x"26",
         10732 => x"57",
         10733 => x"08",
         10734 => x"38",
         10735 => x"56",
         10736 => x"80",
         10737 => x"91",
         10738 => x"95",
         10739 => x"2a",
         10740 => x"74",
         10741 => x"99",
         10742 => x"80",
         10743 => x"ce",
         10744 => x"80",
         10745 => x"c6",
         10746 => x"80",
         10747 => x"be",
         10748 => x"7a",
         10749 => x"ff",
         10750 => x"16",
         10751 => x"33",
         10752 => x"71",
         10753 => x"7a",
         10754 => x"0c",
         10755 => x"11",
         10756 => x"33",
         10757 => x"71",
         10758 => x"81",
         10759 => x"72",
         10760 => x"75",
         10761 => x"62",
         10762 => x"45",
         10763 => x"55",
         10764 => x"58",
         10765 => x"1b",
         10766 => x"23",
         10767 => x"34",
         10768 => x"1b",
         10769 => x"9c",
         10770 => x"0b",
         10771 => x"a8",
         10772 => x"80",
         10773 => x"fd",
         10774 => x"51",
         10775 => x"84",
         10776 => x"79",
         10777 => x"57",
         10778 => x"38",
         10779 => x"74",
         10780 => x"ff",
         10781 => x"84",
         10782 => x"5d",
         10783 => x"08",
         10784 => x"cb",
         10785 => x"84",
         10786 => x"fb",
         10787 => x"bb",
         10788 => x"2e",
         10789 => x"80",
         10790 => x"75",
         10791 => x"a0",
         10792 => x"84",
         10793 => x"38",
         10794 => x"fe",
         10795 => x"08",
         10796 => x"76",
         10797 => x"38",
         10798 => x"17",
         10799 => x"33",
         10800 => x"74",
         10801 => x"7c",
         10802 => x"26",
         10803 => x"80",
         10804 => x"5f",
         10805 => x"b4",
         10806 => x"2e",
         10807 => x"16",
         10808 => x"7d",
         10809 => x"06",
         10810 => x"81",
         10811 => x"b8",
         10812 => x"16",
         10813 => x"a3",
         10814 => x"bb",
         10815 => x"2e",
         10816 => x"57",
         10817 => x"b4",
         10818 => x"56",
         10819 => x"90",
         10820 => x"7b",
         10821 => x"b5",
         10822 => x"0c",
         10823 => x"80",
         10824 => x"34",
         10825 => x"17",
         10826 => x"39",
         10827 => x"94",
         10828 => x"98",
         10829 => x"2b",
         10830 => x"5d",
         10831 => x"0b",
         10832 => x"80",
         10833 => x"34",
         10834 => x"17",
         10835 => x"0b",
         10836 => x"66",
         10837 => x"8b",
         10838 => x"67",
         10839 => x"0b",
         10840 => x"80",
         10841 => x"34",
         10842 => x"7c",
         10843 => x"81",
         10844 => x"38",
         10845 => x"77",
         10846 => x"76",
         10847 => x"75",
         10848 => x"59",
         10849 => x"f8",
         10850 => x"fe",
         10851 => x"08",
         10852 => x"59",
         10853 => x"27",
         10854 => x"8a",
         10855 => x"71",
         10856 => x"08",
         10857 => x"74",
         10858 => x"d8",
         10859 => x"2a",
         10860 => x"1c",
         10861 => x"54",
         10862 => x"52",
         10863 => x"51",
         10864 => x"3f",
         10865 => x"08",
         10866 => x"e2",
         10867 => x"80",
         10868 => x"da",
         10869 => x"b4",
         10870 => x"b8",
         10871 => x"81",
         10872 => x"58",
         10873 => x"3f",
         10874 => x"08",
         10875 => x"81",
         10876 => x"38",
         10877 => x"08",
         10878 => x"b4",
         10879 => x"17",
         10880 => x"bb",
         10881 => x"55",
         10882 => x"08",
         10883 => x"38",
         10884 => x"55",
         10885 => x"09",
         10886 => x"cf",
         10887 => x"b4",
         10888 => x"17",
         10889 => x"77",
         10890 => x"33",
         10891 => x"fb",
         10892 => x"fd",
         10893 => x"bb",
         10894 => x"80",
         10895 => x"ee",
         10896 => x"fd",
         10897 => x"3d",
         10898 => x"65",
         10899 => x"5b",
         10900 => x"0c",
         10901 => x"80",
         10902 => x"78",
         10903 => x"80",
         10904 => x"75",
         10905 => x"80",
         10906 => x"86",
         10907 => x"1a",
         10908 => x"7a",
         10909 => x"b4",
         10910 => x"74",
         10911 => x"76",
         10912 => x"91",
         10913 => x"74",
         10914 => x"90",
         10915 => x"06",
         10916 => x"76",
         10917 => x"c8",
         10918 => x"08",
         10919 => x"71",
         10920 => x"79",
         10921 => x"ca",
         10922 => x"2e",
         10923 => x"75",
         10924 => x"5c",
         10925 => x"38",
         10926 => x"22",
         10927 => x"89",
         10928 => x"58",
         10929 => x"75",
         10930 => x"88",
         10931 => x"81",
         10932 => x"c3",
         10933 => x"2e",
         10934 => x"74",
         10935 => x"7e",
         10936 => x"08",
         10937 => x"19",
         10938 => x"5c",
         10939 => x"27",
         10940 => x"8a",
         10941 => x"78",
         10942 => x"08",
         10943 => x"74",
         10944 => x"93",
         10945 => x"7a",
         10946 => x"57",
         10947 => x"80",
         10948 => x"1c",
         10949 => x"27",
         10950 => x"7c",
         10951 => x"54",
         10952 => x"52",
         10953 => x"51",
         10954 => x"3f",
         10955 => x"08",
         10956 => x"90",
         10957 => x"98",
         10958 => x"80",
         10959 => x"87",
         10960 => x"2b",
         10961 => x"31",
         10962 => x"7f",
         10963 => x"94",
         10964 => x"70",
         10965 => x"0c",
         10966 => x"fe",
         10967 => x"56",
         10968 => x"84",
         10969 => x"0d",
         10970 => x"bb",
         10971 => x"3d",
         10972 => x"5a",
         10973 => x"9c",
         10974 => x"75",
         10975 => x"c8",
         10976 => x"33",
         10977 => x"a8",
         10978 => x"5b",
         10979 => x"a3",
         10980 => x"75",
         10981 => x"81",
         10982 => x"ff",
         10983 => x"84",
         10984 => x"81",
         10985 => x"19",
         10986 => x"06",
         10987 => x"1a",
         10988 => x"81",
         10989 => x"7a",
         10990 => x"33",
         10991 => x"ec",
         10992 => x"84",
         10993 => x"38",
         10994 => x"0c",
         10995 => x"56",
         10996 => x"06",
         10997 => x"31",
         10998 => x"77",
         10999 => x"79",
         11000 => x"7a",
         11001 => x"57",
         11002 => x"80",
         11003 => x"38",
         11004 => x"05",
         11005 => x"70",
         11006 => x"34",
         11007 => x"75",
         11008 => x"c1",
         11009 => x"81",
         11010 => x"78",
         11011 => x"5a",
         11012 => x"56",
         11013 => x"fe",
         11014 => x"19",
         11015 => x"51",
         11016 => x"3f",
         11017 => x"08",
         11018 => x"39",
         11019 => x"51",
         11020 => x"3f",
         11021 => x"08",
         11022 => x"74",
         11023 => x"74",
         11024 => x"57",
         11025 => x"9c",
         11026 => x"31",
         11027 => x"27",
         11028 => x"84",
         11029 => x"29",
         11030 => x"58",
         11031 => x"70",
         11032 => x"33",
         11033 => x"05",
         11034 => x"15",
         11035 => x"2e",
         11036 => x"75",
         11037 => x"57",
         11038 => x"81",
         11039 => x"ff",
         11040 => x"da",
         11041 => x"39",
         11042 => x"1a",
         11043 => x"84",
         11044 => x"90",
         11045 => x"82",
         11046 => x"34",
         11047 => x"bb",
         11048 => x"3d",
         11049 => x"3d",
         11050 => x"66",
         11051 => x"5c",
         11052 => x"0c",
         11053 => x"80",
         11054 => x"78",
         11055 => x"80",
         11056 => x"75",
         11057 => x"80",
         11058 => x"86",
         11059 => x"1a",
         11060 => x"79",
         11061 => x"a8",
         11062 => x"74",
         11063 => x"76",
         11064 => x"91",
         11065 => x"74",
         11066 => x"90",
         11067 => x"81",
         11068 => x"58",
         11069 => x"76",
         11070 => x"a9",
         11071 => x"08",
         11072 => x"57",
         11073 => x"84",
         11074 => x"5b",
         11075 => x"82",
         11076 => x"83",
         11077 => x"7c",
         11078 => x"7f",
         11079 => x"ff",
         11080 => x"2a",
         11081 => x"7c",
         11082 => x"82",
         11083 => x"19",
         11084 => x"80",
         11085 => x"38",
         11086 => x"83",
         11087 => x"ff",
         11088 => x"38",
         11089 => x"0c",
         11090 => x"85",
         11091 => x"1a",
         11092 => x"90",
         11093 => x"98",
         11094 => x"80",
         11095 => x"f9",
         11096 => x"08",
         11097 => x"19",
         11098 => x"5d",
         11099 => x"27",
         11100 => x"8a",
         11101 => x"78",
         11102 => x"08",
         11103 => x"74",
         11104 => x"a6",
         11105 => x"7b",
         11106 => x"5c",
         11107 => x"81",
         11108 => x"1d",
         11109 => x"27",
         11110 => x"7d",
         11111 => x"54",
         11112 => x"52",
         11113 => x"51",
         11114 => x"3f",
         11115 => x"08",
         11116 => x"9c",
         11117 => x"31",
         11118 => x"27",
         11119 => x"80",
         11120 => x"77",
         11121 => x"05",
         11122 => x"75",
         11123 => x"57",
         11124 => x"81",
         11125 => x"ff",
         11126 => x"ef",
         11127 => x"33",
         11128 => x"5d",
         11129 => x"34",
         11130 => x"58",
         11131 => x"7f",
         11132 => x"0c",
         11133 => x"1b",
         11134 => x"71",
         11135 => x"8c",
         11136 => x"5a",
         11137 => x"74",
         11138 => x"38",
         11139 => x"8c",
         11140 => x"fd",
         11141 => x"19",
         11142 => x"80",
         11143 => x"7a",
         11144 => x"80",
         11145 => x"bb",
         11146 => x"3d",
         11147 => x"84",
         11148 => x"91",
         11149 => x"9c",
         11150 => x"2e",
         11151 => x"19",
         11152 => x"8c",
         11153 => x"9b",
         11154 => x"7b",
         11155 => x"52",
         11156 => x"51",
         11157 => x"3f",
         11158 => x"08",
         11159 => x"94",
         11160 => x"7b",
         11161 => x"76",
         11162 => x"84",
         11163 => x"59",
         11164 => x"27",
         11165 => x"58",
         11166 => x"a8",
         11167 => x"56",
         11168 => x"2e",
         11169 => x"70",
         11170 => x"33",
         11171 => x"05",
         11172 => x"16",
         11173 => x"38",
         11174 => x"ff",
         11175 => x"79",
         11176 => x"fe",
         11177 => x"19",
         11178 => x"51",
         11179 => x"3f",
         11180 => x"08",
         11181 => x"84",
         11182 => x"38",
         11183 => x"58",
         11184 => x"76",
         11185 => x"ff",
         11186 => x"84",
         11187 => x"55",
         11188 => x"08",
         11189 => x"e4",
         11190 => x"9c",
         11191 => x"a8",
         11192 => x"18",
         11193 => x"98",
         11194 => x"bb",
         11195 => x"38",
         11196 => x"80",
         11197 => x"75",
         11198 => x"7f",
         11199 => x"39",
         11200 => x"51",
         11201 => x"3f",
         11202 => x"08",
         11203 => x"74",
         11204 => x"74",
         11205 => x"57",
         11206 => x"81",
         11207 => x"34",
         11208 => x"bb",
         11209 => x"3d",
         11210 => x"0b",
         11211 => x"82",
         11212 => x"84",
         11213 => x"0d",
         11214 => x"0d",
         11215 => x"57",
         11216 => x"9f",
         11217 => x"56",
         11218 => x"97",
         11219 => x"55",
         11220 => x"8f",
         11221 => x"22",
         11222 => x"5a",
         11223 => x"2e",
         11224 => x"80",
         11225 => x"76",
         11226 => x"ee",
         11227 => x"33",
         11228 => x"81",
         11229 => x"7a",
         11230 => x"de",
         11231 => x"2b",
         11232 => x"24",
         11233 => x"7b",
         11234 => x"58",
         11235 => x"08",
         11236 => x"38",
         11237 => x"17",
         11238 => x"5c",
         11239 => x"2e",
         11240 => x"81",
         11241 => x"54",
         11242 => x"16",
         11243 => x"33",
         11244 => x"f8",
         11245 => x"84",
         11246 => x"85",
         11247 => x"81",
         11248 => x"17",
         11249 => x"78",
         11250 => x"a4",
         11251 => x"11",
         11252 => x"56",
         11253 => x"18",
         11254 => x"88",
         11255 => x"83",
         11256 => x"5d",
         11257 => x"9a",
         11258 => x"88",
         11259 => x"9b",
         11260 => x"17",
         11261 => x"19",
         11262 => x"74",
         11263 => x"c8",
         11264 => x"08",
         11265 => x"34",
         11266 => x"5b",
         11267 => x"34",
         11268 => x"56",
         11269 => x"34",
         11270 => x"59",
         11271 => x"34",
         11272 => x"80",
         11273 => x"34",
         11274 => x"18",
         11275 => x"0b",
         11276 => x"80",
         11277 => x"34",
         11278 => x"18",
         11279 => x"81",
         11280 => x"34",
         11281 => x"98",
         11282 => x"bb",
         11283 => x"19",
         11284 => x"06",
         11285 => x"90",
         11286 => x"55",
         11287 => x"84",
         11288 => x"0d",
         11289 => x"b4",
         11290 => x"b8",
         11291 => x"81",
         11292 => x"5b",
         11293 => x"3f",
         11294 => x"bb",
         11295 => x"2e",
         11296 => x"fe",
         11297 => x"bb",
         11298 => x"17",
         11299 => x"08",
         11300 => x"31",
         11301 => x"08",
         11302 => x"a0",
         11303 => x"fe",
         11304 => x"16",
         11305 => x"82",
         11306 => x"06",
         11307 => x"81",
         11308 => x"08",
         11309 => x"05",
         11310 => x"81",
         11311 => x"ff",
         11312 => x"79",
         11313 => x"39",
         11314 => x"55",
         11315 => x"34",
         11316 => x"56",
         11317 => x"34",
         11318 => x"55",
         11319 => x"74",
         11320 => x"7a",
         11321 => x"74",
         11322 => x"75",
         11323 => x"74",
         11324 => x"78",
         11325 => x"80",
         11326 => x"0b",
         11327 => x"a1",
         11328 => x"34",
         11329 => x"99",
         11330 => x"0b",
         11331 => x"80",
         11332 => x"34",
         11333 => x"0b",
         11334 => x"7b",
         11335 => x"be",
         11336 => x"84",
         11337 => x"33",
         11338 => x"5b",
         11339 => x"19",
         11340 => x"39",
         11341 => x"51",
         11342 => x"3f",
         11343 => x"08",
         11344 => x"74",
         11345 => x"74",
         11346 => x"57",
         11347 => x"81",
         11348 => x"08",
         11349 => x"52",
         11350 => x"33",
         11351 => x"93",
         11352 => x"55",
         11353 => x"08",
         11354 => x"90",
         11355 => x"ff",
         11356 => x"90",
         11357 => x"a0",
         11358 => x"56",
         11359 => x"77",
         11360 => x"06",
         11361 => x"fc",
         11362 => x"3d",
         11363 => x"52",
         11364 => x"3f",
         11365 => x"08",
         11366 => x"84",
         11367 => x"89",
         11368 => x"2e",
         11369 => x"08",
         11370 => x"2e",
         11371 => x"33",
         11372 => x"2e",
         11373 => x"13",
         11374 => x"22",
         11375 => x"77",
         11376 => x"80",
         11377 => x"75",
         11378 => x"38",
         11379 => x"73",
         11380 => x"0c",
         11381 => x"04",
         11382 => x"51",
         11383 => x"3f",
         11384 => x"08",
         11385 => x"72",
         11386 => x"75",
         11387 => x"d5",
         11388 => x"0d",
         11389 => x"5b",
         11390 => x"80",
         11391 => x"75",
         11392 => x"57",
         11393 => x"26",
         11394 => x"ba",
         11395 => x"70",
         11396 => x"ba",
         11397 => x"84",
         11398 => x"51",
         11399 => x"90",
         11400 => x"e2",
         11401 => x"0b",
         11402 => x"0c",
         11403 => x"04",
         11404 => x"bb",
         11405 => x"3d",
         11406 => x"33",
         11407 => x"81",
         11408 => x"53",
         11409 => x"26",
         11410 => x"19",
         11411 => x"06",
         11412 => x"54",
         11413 => x"80",
         11414 => x"0b",
         11415 => x"5b",
         11416 => x"79",
         11417 => x"70",
         11418 => x"33",
         11419 => x"05",
         11420 => x"9f",
         11421 => x"52",
         11422 => x"89",
         11423 => x"70",
         11424 => x"53",
         11425 => x"13",
         11426 => x"26",
         11427 => x"13",
         11428 => x"06",
         11429 => x"30",
         11430 => x"55",
         11431 => x"2e",
         11432 => x"85",
         11433 => x"be",
         11434 => x"32",
         11435 => x"72",
         11436 => x"76",
         11437 => x"52",
         11438 => x"92",
         11439 => x"84",
         11440 => x"83",
         11441 => x"99",
         11442 => x"fe",
         11443 => x"83",
         11444 => x"77",
         11445 => x"fe",
         11446 => x"3d",
         11447 => x"98",
         11448 => x"52",
         11449 => x"d2",
         11450 => x"bb",
         11451 => x"84",
         11452 => x"80",
         11453 => x"74",
         11454 => x"0c",
         11455 => x"04",
         11456 => x"52",
         11457 => x"05",
         11458 => x"3f",
         11459 => x"08",
         11460 => x"84",
         11461 => x"38",
         11462 => x"05",
         11463 => x"2b",
         11464 => x"77",
         11465 => x"38",
         11466 => x"33",
         11467 => x"81",
         11468 => x"75",
         11469 => x"38",
         11470 => x"11",
         11471 => x"33",
         11472 => x"07",
         11473 => x"5a",
         11474 => x"79",
         11475 => x"38",
         11476 => x"0c",
         11477 => x"84",
         11478 => x"0d",
         11479 => x"84",
         11480 => x"09",
         11481 => x"8f",
         11482 => x"84",
         11483 => x"98",
         11484 => x"95",
         11485 => x"17",
         11486 => x"2b",
         11487 => x"07",
         11488 => x"1b",
         11489 => x"cc",
         11490 => x"98",
         11491 => x"74",
         11492 => x"0c",
         11493 => x"04",
         11494 => x"0d",
         11495 => x"08",
         11496 => x"08",
         11497 => x"7c",
         11498 => x"80",
         11499 => x"b4",
         11500 => x"e5",
         11501 => x"84",
         11502 => x"84",
         11503 => x"bb",
         11504 => x"c8",
         11505 => x"d9",
         11506 => x"61",
         11507 => x"80",
         11508 => x"58",
         11509 => x"08",
         11510 => x"80",
         11511 => x"38",
         11512 => x"98",
         11513 => x"a0",
         11514 => x"ff",
         11515 => x"84",
         11516 => x"59",
         11517 => x"08",
         11518 => x"60",
         11519 => x"08",
         11520 => x"16",
         11521 => x"b1",
         11522 => x"84",
         11523 => x"33",
         11524 => x"83",
         11525 => x"54",
         11526 => x"16",
         11527 => x"33",
         11528 => x"88",
         11529 => x"84",
         11530 => x"85",
         11531 => x"81",
         11532 => x"17",
         11533 => x"d4",
         11534 => x"3d",
         11535 => x"33",
         11536 => x"71",
         11537 => x"63",
         11538 => x"40",
         11539 => x"78",
         11540 => x"da",
         11541 => x"db",
         11542 => x"52",
         11543 => x"a4",
         11544 => x"bb",
         11545 => x"84",
         11546 => x"82",
         11547 => x"52",
         11548 => x"aa",
         11549 => x"bb",
         11550 => x"84",
         11551 => x"bb",
         11552 => x"3d",
         11553 => x"33",
         11554 => x"71",
         11555 => x"63",
         11556 => x"58",
         11557 => x"7d",
         11558 => x"fd",
         11559 => x"2e",
         11560 => x"bb",
         11561 => x"7a",
         11562 => x"a1",
         11563 => x"84",
         11564 => x"bb",
         11565 => x"2e",
         11566 => x"78",
         11567 => x"d8",
         11568 => x"c8",
         11569 => x"3d",
         11570 => x"52",
         11571 => x"be",
         11572 => x"7f",
         11573 => x"5b",
         11574 => x"2e",
         11575 => x"1f",
         11576 => x"81",
         11577 => x"5f",
         11578 => x"f5",
         11579 => x"56",
         11580 => x"81",
         11581 => x"80",
         11582 => x"7e",
         11583 => x"56",
         11584 => x"e6",
         11585 => x"ff",
         11586 => x"59",
         11587 => x"75",
         11588 => x"76",
         11589 => x"18",
         11590 => x"08",
         11591 => x"af",
         11592 => x"da",
         11593 => x"79",
         11594 => x"77",
         11595 => x"8a",
         11596 => x"84",
         11597 => x"70",
         11598 => x"e6",
         11599 => x"08",
         11600 => x"59",
         11601 => x"7e",
         11602 => x"38",
         11603 => x"17",
         11604 => x"5f",
         11605 => x"38",
         11606 => x"7a",
         11607 => x"38",
         11608 => x"7a",
         11609 => x"76",
         11610 => x"33",
         11611 => x"05",
         11612 => x"17",
         11613 => x"26",
         11614 => x"7c",
         11615 => x"5e",
         11616 => x"2e",
         11617 => x"81",
         11618 => x"59",
         11619 => x"78",
         11620 => x"0c",
         11621 => x"0d",
         11622 => x"33",
         11623 => x"71",
         11624 => x"90",
         11625 => x"07",
         11626 => x"fd",
         11627 => x"16",
         11628 => x"33",
         11629 => x"71",
         11630 => x"79",
         11631 => x"3d",
         11632 => x"80",
         11633 => x"ff",
         11634 => x"84",
         11635 => x"59",
         11636 => x"08",
         11637 => x"96",
         11638 => x"39",
         11639 => x"16",
         11640 => x"16",
         11641 => x"17",
         11642 => x"ff",
         11643 => x"81",
         11644 => x"84",
         11645 => x"38",
         11646 => x"08",
         11647 => x"b4",
         11648 => x"17",
         11649 => x"bb",
         11650 => x"55",
         11651 => x"08",
         11652 => x"38",
         11653 => x"55",
         11654 => x"09",
         11655 => x"f6",
         11656 => x"b4",
         11657 => x"17",
         11658 => x"7d",
         11659 => x"33",
         11660 => x"f7",
         11661 => x"fb",
         11662 => x"18",
         11663 => x"08",
         11664 => x"af",
         11665 => x"0b",
         11666 => x"33",
         11667 => x"83",
         11668 => x"70",
         11669 => x"43",
         11670 => x"5a",
         11671 => x"09",
         11672 => x"e8",
         11673 => x"39",
         11674 => x"08",
         11675 => x"59",
         11676 => x"7c",
         11677 => x"5e",
         11678 => x"27",
         11679 => x"80",
         11680 => x"18",
         11681 => x"5a",
         11682 => x"70",
         11683 => x"34",
         11684 => x"d4",
         11685 => x"39",
         11686 => x"7c",
         11687 => x"bb",
         11688 => x"e4",
         11689 => x"f5",
         11690 => x"7f",
         11691 => x"58",
         11692 => x"9f",
         11693 => x"56",
         11694 => x"97",
         11695 => x"55",
         11696 => x"8f",
         11697 => x"22",
         11698 => x"5b",
         11699 => x"2e",
         11700 => x"80",
         11701 => x"77",
         11702 => x"fb",
         11703 => x"33",
         11704 => x"f3",
         11705 => x"08",
         11706 => x"26",
         11707 => x"94",
         11708 => x"80",
         11709 => x"2e",
         11710 => x"7b",
         11711 => x"70",
         11712 => x"5c",
         11713 => x"2e",
         11714 => x"77",
         11715 => x"51",
         11716 => x"3f",
         11717 => x"08",
         11718 => x"54",
         11719 => x"55",
         11720 => x"3f",
         11721 => x"08",
         11722 => x"da",
         11723 => x"76",
         11724 => x"19",
         11725 => x"31",
         11726 => x"58",
         11727 => x"80",
         11728 => x"38",
         11729 => x"80",
         11730 => x"78",
         11731 => x"08",
         11732 => x"0c",
         11733 => x"70",
         11734 => x"06",
         11735 => x"7a",
         11736 => x"cc",
         11737 => x"76",
         11738 => x"b2",
         11739 => x"84",
         11740 => x"bb",
         11741 => x"2e",
         11742 => x"ff",
         11743 => x"38",
         11744 => x"83",
         11745 => x"55",
         11746 => x"08",
         11747 => x"38",
         11748 => x"0c",
         11749 => x"84",
         11750 => x"59",
         11751 => x"19",
         11752 => x"78",
         11753 => x"58",
         11754 => x"a9",
         11755 => x"17",
         11756 => x"fe",
         11757 => x"58",
         11758 => x"82",
         11759 => x"18",
         11760 => x"29",
         11761 => x"05",
         11762 => x"11",
         11763 => x"7a",
         11764 => x"b3",
         11765 => x"08",
         11766 => x"08",
         11767 => x"27",
         11768 => x"8c",
         11769 => x"17",
         11770 => x"07",
         11771 => x"18",
         11772 => x"ff",
         11773 => x"80",
         11774 => x"38",
         11775 => x"56",
         11776 => x"81",
         11777 => x"17",
         11778 => x"2b",
         11779 => x"56",
         11780 => x"25",
         11781 => x"54",
         11782 => x"52",
         11783 => x"33",
         11784 => x"86",
         11785 => x"bb",
         11786 => x"38",
         11787 => x"80",
         11788 => x"74",
         11789 => x"81",
         11790 => x"77",
         11791 => x"11",
         11792 => x"ff",
         11793 => x"84",
         11794 => x"80",
         11795 => x"38",
         11796 => x"18",
         11797 => x"74",
         11798 => x"0c",
         11799 => x"04",
         11800 => x"70",
         11801 => x"06",
         11802 => x"fd",
         11803 => x"94",
         11804 => x"59",
         11805 => x"7a",
         11806 => x"06",
         11807 => x"79",
         11808 => x"fe",
         11809 => x"0b",
         11810 => x"88",
         11811 => x"75",
         11812 => x"c7",
         11813 => x"18",
         11814 => x"2e",
         11815 => x"fd",
         11816 => x"9c",
         11817 => x"0b",
         11818 => x"0c",
         11819 => x"04",
         11820 => x"51",
         11821 => x"3f",
         11822 => x"08",
         11823 => x"39",
         11824 => x"51",
         11825 => x"3f",
         11826 => x"08",
         11827 => x"74",
         11828 => x"74",
         11829 => x"58",
         11830 => x"75",
         11831 => x"ff",
         11832 => x"84",
         11833 => x"56",
         11834 => x"08",
         11835 => x"38",
         11836 => x"08",
         11837 => x"d8",
         11838 => x"84",
         11839 => x"0c",
         11840 => x"0c",
         11841 => x"82",
         11842 => x"34",
         11843 => x"bb",
         11844 => x"3d",
         11845 => x"3d",
         11846 => x"89",
         11847 => x"2e",
         11848 => x"53",
         11849 => x"05",
         11850 => x"84",
         11851 => x"8c",
         11852 => x"84",
         11853 => x"bb",
         11854 => x"2e",
         11855 => x"76",
         11856 => x"73",
         11857 => x"0c",
         11858 => x"04",
         11859 => x"7d",
         11860 => x"ff",
         11861 => x"84",
         11862 => x"55",
         11863 => x"08",
         11864 => x"ab",
         11865 => x"98",
         11866 => x"80",
         11867 => x"38",
         11868 => x"70",
         11869 => x"06",
         11870 => x"80",
         11871 => x"38",
         11872 => x"9b",
         11873 => x"12",
         11874 => x"2b",
         11875 => x"33",
         11876 => x"55",
         11877 => x"2e",
         11878 => x"88",
         11879 => x"58",
         11880 => x"84",
         11881 => x"52",
         11882 => x"9a",
         11883 => x"bb",
         11884 => x"74",
         11885 => x"38",
         11886 => x"ff",
         11887 => x"76",
         11888 => x"39",
         11889 => x"76",
         11890 => x"39",
         11891 => x"94",
         11892 => x"98",
         11893 => x"2b",
         11894 => x"88",
         11895 => x"5a",
         11896 => x"fa",
         11897 => x"55",
         11898 => x"80",
         11899 => x"74",
         11900 => x"80",
         11901 => x"72",
         11902 => x"80",
         11903 => x"86",
         11904 => x"16",
         11905 => x"71",
         11906 => x"38",
         11907 => x"57",
         11908 => x"73",
         11909 => x"84",
         11910 => x"88",
         11911 => x"81",
         11912 => x"ff",
         11913 => x"84",
         11914 => x"81",
         11915 => x"dc",
         11916 => x"08",
         11917 => x"39",
         11918 => x"7a",
         11919 => x"89",
         11920 => x"2e",
         11921 => x"08",
         11922 => x"2e",
         11923 => x"33",
         11924 => x"2e",
         11925 => x"14",
         11926 => x"22",
         11927 => x"78",
         11928 => x"38",
         11929 => x"59",
         11930 => x"80",
         11931 => x"80",
         11932 => x"38",
         11933 => x"51",
         11934 => x"3f",
         11935 => x"08",
         11936 => x"84",
         11937 => x"b5",
         11938 => x"84",
         11939 => x"76",
         11940 => x"ff",
         11941 => x"72",
         11942 => x"ff",
         11943 => x"84",
         11944 => x"84",
         11945 => x"70",
         11946 => x"2c",
         11947 => x"08",
         11948 => x"54",
         11949 => x"84",
         11950 => x"0d",
         11951 => x"53",
         11952 => x"ff",
         11953 => x"72",
         11954 => x"ff",
         11955 => x"84",
         11956 => x"84",
         11957 => x"70",
         11958 => x"2c",
         11959 => x"08",
         11960 => x"54",
         11961 => x"52",
         11962 => x"97",
         11963 => x"bb",
         11964 => x"bb",
         11965 => x"3d",
         11966 => x"14",
         11967 => x"fe",
         11968 => x"bb",
         11969 => x"06",
         11970 => x"d8",
         11971 => x"08",
         11972 => x"d2",
         11973 => x"0d",
         11974 => x"53",
         11975 => x"53",
         11976 => x"56",
         11977 => x"84",
         11978 => x"55",
         11979 => x"08",
         11980 => x"38",
         11981 => x"84",
         11982 => x"0d",
         11983 => x"75",
         11984 => x"9a",
         11985 => x"84",
         11986 => x"bb",
         11987 => x"38",
         11988 => x"05",
         11989 => x"2b",
         11990 => x"74",
         11991 => x"76",
         11992 => x"38",
         11993 => x"51",
         11994 => x"3f",
         11995 => x"84",
         11996 => x"0d",
         11997 => x"84",
         11998 => x"95",
         11999 => x"ed",
         12000 => x"68",
         12001 => x"53",
         12002 => x"05",
         12003 => x"51",
         12004 => x"84",
         12005 => x"5a",
         12006 => x"08",
         12007 => x"75",
         12008 => x"9c",
         12009 => x"11",
         12010 => x"59",
         12011 => x"75",
         12012 => x"38",
         12013 => x"79",
         12014 => x"0c",
         12015 => x"04",
         12016 => x"08",
         12017 => x"5b",
         12018 => x"82",
         12019 => x"a8",
         12020 => x"bb",
         12021 => x"5d",
         12022 => x"c1",
         12023 => x"1d",
         12024 => x"56",
         12025 => x"76",
         12026 => x"38",
         12027 => x"78",
         12028 => x"81",
         12029 => x"54",
         12030 => x"17",
         12031 => x"33",
         12032 => x"a8",
         12033 => x"84",
         12034 => x"85",
         12035 => x"81",
         12036 => x"18",
         12037 => x"5b",
         12038 => x"cc",
         12039 => x"5e",
         12040 => x"82",
         12041 => x"17",
         12042 => x"11",
         12043 => x"33",
         12044 => x"71",
         12045 => x"81",
         12046 => x"72",
         12047 => x"75",
         12048 => x"ff",
         12049 => x"06",
         12050 => x"70",
         12051 => x"05",
         12052 => x"83",
         12053 => x"ff",
         12054 => x"43",
         12055 => x"53",
         12056 => x"56",
         12057 => x"38",
         12058 => x"7a",
         12059 => x"84",
         12060 => x"07",
         12061 => x"18",
         12062 => x"bb",
         12063 => x"3d",
         12064 => x"54",
         12065 => x"53",
         12066 => x"53",
         12067 => x"52",
         12068 => x"97",
         12069 => x"84",
         12070 => x"fe",
         12071 => x"bb",
         12072 => x"18",
         12073 => x"08",
         12074 => x"31",
         12075 => x"08",
         12076 => x"a0",
         12077 => x"fe",
         12078 => x"17",
         12079 => x"82",
         12080 => x"06",
         12081 => x"81",
         12082 => x"08",
         12083 => x"05",
         12084 => x"81",
         12085 => x"fe",
         12086 => x"77",
         12087 => x"39",
         12088 => x"92",
         12089 => x"75",
         12090 => x"ff",
         12091 => x"84",
         12092 => x"ff",
         12093 => x"38",
         12094 => x"08",
         12095 => x"f7",
         12096 => x"84",
         12097 => x"84",
         12098 => x"07",
         12099 => x"05",
         12100 => x"5a",
         12101 => x"9c",
         12102 => x"26",
         12103 => x"7f",
         12104 => x"18",
         12105 => x"33",
         12106 => x"77",
         12107 => x"fe",
         12108 => x"17",
         12109 => x"11",
         12110 => x"71",
         12111 => x"70",
         12112 => x"25",
         12113 => x"83",
         12114 => x"1f",
         12115 => x"59",
         12116 => x"78",
         12117 => x"fe",
         12118 => x"5a",
         12119 => x"81",
         12120 => x"7a",
         12121 => x"94",
         12122 => x"17",
         12123 => x"58",
         12124 => x"34",
         12125 => x"82",
         12126 => x"e7",
         12127 => x"0d",
         12128 => x"57",
         12129 => x"9f",
         12130 => x"56",
         12131 => x"97",
         12132 => x"55",
         12133 => x"8f",
         12134 => x"22",
         12135 => x"5a",
         12136 => x"2e",
         12137 => x"80",
         12138 => x"76",
         12139 => x"91",
         12140 => x"76",
         12141 => x"90",
         12142 => x"81",
         12143 => x"56",
         12144 => x"74",
         12145 => x"eb",
         12146 => x"08",
         12147 => x"19",
         12148 => x"dd",
         12149 => x"fb",
         12150 => x"08",
         12151 => x"55",
         12152 => x"89",
         12153 => x"08",
         12154 => x"d8",
         12155 => x"80",
         12156 => x"0c",
         12157 => x"8c",
         12158 => x"80",
         12159 => x"74",
         12160 => x"76",
         12161 => x"98",
         12162 => x"80",
         12163 => x"81",
         12164 => x"08",
         12165 => x"52",
         12166 => x"33",
         12167 => x"fa",
         12168 => x"bb",
         12169 => x"2e",
         12170 => x"81",
         12171 => x"19",
         12172 => x"75",
         12173 => x"0c",
         12174 => x"04",
         12175 => x"79",
         12176 => x"38",
         12177 => x"51",
         12178 => x"3f",
         12179 => x"08",
         12180 => x"84",
         12181 => x"80",
         12182 => x"bb",
         12183 => x"2e",
         12184 => x"84",
         12185 => x"ff",
         12186 => x"38",
         12187 => x"52",
         12188 => x"85",
         12189 => x"bb",
         12190 => x"d8",
         12191 => x"08",
         12192 => x"19",
         12193 => x"59",
         12194 => x"ff",
         12195 => x"16",
         12196 => x"84",
         12197 => x"07",
         12198 => x"18",
         12199 => x"78",
         12200 => x"a0",
         12201 => x"81",
         12202 => x"fe",
         12203 => x"84",
         12204 => x"81",
         12205 => x"fd",
         12206 => x"78",
         12207 => x"fd",
         12208 => x"0b",
         12209 => x"5a",
         12210 => x"80",
         12211 => x"0c",
         12212 => x"98",
         12213 => x"77",
         12214 => x"83",
         12215 => x"84",
         12216 => x"81",
         12217 => x"bb",
         12218 => x"2e",
         12219 => x"76",
         12220 => x"7a",
         12221 => x"84",
         12222 => x"08",
         12223 => x"38",
         12224 => x"08",
         12225 => x"79",
         12226 => x"55",
         12227 => x"bb",
         12228 => x"81",
         12229 => x"bb",
         12230 => x"18",
         12231 => x"96",
         12232 => x"2e",
         12233 => x"53",
         12234 => x"51",
         12235 => x"3f",
         12236 => x"08",
         12237 => x"84",
         12238 => x"38",
         12239 => x"51",
         12240 => x"3f",
         12241 => x"08",
         12242 => x"84",
         12243 => x"80",
         12244 => x"bb",
         12245 => x"2e",
         12246 => x"84",
         12247 => x"ff",
         12248 => x"38",
         12249 => x"52",
         12250 => x"83",
         12251 => x"bb",
         12252 => x"f6",
         12253 => x"08",
         12254 => x"19",
         12255 => x"59",
         12256 => x"90",
         12257 => x"94",
         12258 => x"17",
         12259 => x"55",
         12260 => x"34",
         12261 => x"7a",
         12262 => x"38",
         12263 => x"57",
         12264 => x"59",
         12265 => x"81",
         12266 => x"39",
         12267 => x"19",
         12268 => x"fc",
         12269 => x"57",
         12270 => x"18",
         12271 => x"06",
         12272 => x"19",
         12273 => x"fc",
         12274 => x"0b",
         12275 => x"5a",
         12276 => x"39",
         12277 => x"08",
         12278 => x"5a",
         12279 => x"39",
         12280 => x"19",
         12281 => x"fd",
         12282 => x"bb",
         12283 => x"ff",
         12284 => x"57",
         12285 => x"db",
         12286 => x"53",
         12287 => x"9c",
         12288 => x"3d",
         12289 => x"b4",
         12290 => x"84",
         12291 => x"bb",
         12292 => x"2e",
         12293 => x"84",
         12294 => x"a7",
         12295 => x"7d",
         12296 => x"08",
         12297 => x"70",
         12298 => x"ac",
         12299 => x"bb",
         12300 => x"84",
         12301 => x"de",
         12302 => x"93",
         12303 => x"85",
         12304 => x"59",
         12305 => x"77",
         12306 => x"98",
         12307 => x"7b",
         12308 => x"02",
         12309 => x"33",
         12310 => x"5d",
         12311 => x"7b",
         12312 => x"7d",
         12313 => x"9b",
         12314 => x"12",
         12315 => x"2b",
         12316 => x"41",
         12317 => x"58",
         12318 => x"80",
         12319 => x"84",
         12320 => x"57",
         12321 => x"80",
         12322 => x"56",
         12323 => x"7b",
         12324 => x"38",
         12325 => x"41",
         12326 => x"08",
         12327 => x"70",
         12328 => x"8c",
         12329 => x"bb",
         12330 => x"84",
         12331 => x"fe",
         12332 => x"bb",
         12333 => x"74",
         12334 => x"ed",
         12335 => x"84",
         12336 => x"bb",
         12337 => x"38",
         12338 => x"bb",
         12339 => x"3d",
         12340 => x"16",
         12341 => x"33",
         12342 => x"71",
         12343 => x"7d",
         12344 => x"5d",
         12345 => x"84",
         12346 => x"84",
         12347 => x"84",
         12348 => x"fe",
         12349 => x"08",
         12350 => x"08",
         12351 => x"74",
         12352 => x"d3",
         12353 => x"78",
         12354 => x"cb",
         12355 => x"84",
         12356 => x"bb",
         12357 => x"2e",
         12358 => x"30",
         12359 => x"80",
         12360 => x"7a",
         12361 => x"38",
         12362 => x"95",
         12363 => x"08",
         12364 => x"7b",
         12365 => x"9c",
         12366 => x"26",
         12367 => x"82",
         12368 => x"d2",
         12369 => x"fe",
         12370 => x"84",
         12371 => x"84",
         12372 => x"a7",
         12373 => x"b8",
         12374 => x"19",
         12375 => x"5a",
         12376 => x"76",
         12377 => x"38",
         12378 => x"7a",
         12379 => x"7a",
         12380 => x"06",
         12381 => x"81",
         12382 => x"b8",
         12383 => x"17",
         12384 => x"f2",
         12385 => x"bb",
         12386 => x"2e",
         12387 => x"56",
         12388 => x"b4",
         12389 => x"56",
         12390 => x"9c",
         12391 => x"e5",
         12392 => x"0b",
         12393 => x"90",
         12394 => x"27",
         12395 => x"80",
         12396 => x"ff",
         12397 => x"84",
         12398 => x"56",
         12399 => x"08",
         12400 => x"96",
         12401 => x"2e",
         12402 => x"fe",
         12403 => x"56",
         12404 => x"81",
         12405 => x"08",
         12406 => x"81",
         12407 => x"fe",
         12408 => x"81",
         12409 => x"84",
         12410 => x"09",
         12411 => x"a6",
         12412 => x"84",
         12413 => x"34",
         12414 => x"a8",
         12415 => x"84",
         12416 => x"59",
         12417 => x"18",
         12418 => x"eb",
         12419 => x"33",
         12420 => x"2e",
         12421 => x"fe",
         12422 => x"54",
         12423 => x"a0",
         12424 => x"53",
         12425 => x"17",
         12426 => x"f1",
         12427 => x"58",
         12428 => x"79",
         12429 => x"27",
         12430 => x"74",
         12431 => x"fe",
         12432 => x"84",
         12433 => x"5a",
         12434 => x"08",
         12435 => x"cb",
         12436 => x"84",
         12437 => x"fd",
         12438 => x"bb",
         12439 => x"2e",
         12440 => x"80",
         12441 => x"76",
         12442 => x"d4",
         12443 => x"84",
         12444 => x"9c",
         12445 => x"11",
         12446 => x"58",
         12447 => x"7b",
         12448 => x"38",
         12449 => x"18",
         12450 => x"33",
         12451 => x"7b",
         12452 => x"79",
         12453 => x"26",
         12454 => x"80",
         12455 => x"39",
         12456 => x"f7",
         12457 => x"84",
         12458 => x"95",
         12459 => x"fd",
         12460 => x"3d",
         12461 => x"9f",
         12462 => x"05",
         12463 => x"51",
         12464 => x"3f",
         12465 => x"08",
         12466 => x"84",
         12467 => x"8a",
         12468 => x"bb",
         12469 => x"3d",
         12470 => x"43",
         12471 => x"3d",
         12472 => x"ff",
         12473 => x"84",
         12474 => x"56",
         12475 => x"08",
         12476 => x"0b",
         12477 => x"0c",
         12478 => x"04",
         12479 => x"08",
         12480 => x"81",
         12481 => x"02",
         12482 => x"33",
         12483 => x"81",
         12484 => x"86",
         12485 => x"b9",
         12486 => x"74",
         12487 => x"70",
         12488 => x"83",
         12489 => x"bb",
         12490 => x"57",
         12491 => x"84",
         12492 => x"87",
         12493 => x"84",
         12494 => x"80",
         12495 => x"bb",
         12496 => x"2e",
         12497 => x"75",
         12498 => x"7d",
         12499 => x"08",
         12500 => x"5d",
         12501 => x"80",
         12502 => x"19",
         12503 => x"fe",
         12504 => x"80",
         12505 => x"27",
         12506 => x"17",
         12507 => x"29",
         12508 => x"05",
         12509 => x"b4",
         12510 => x"17",
         12511 => x"79",
         12512 => x"76",
         12513 => x"58",
         12514 => x"55",
         12515 => x"74",
         12516 => x"22",
         12517 => x"27",
         12518 => x"81",
         12519 => x"53",
         12520 => x"17",
         12521 => x"ef",
         12522 => x"bb",
         12523 => x"df",
         12524 => x"58",
         12525 => x"56",
         12526 => x"81",
         12527 => x"08",
         12528 => x"70",
         12529 => x"33",
         12530 => x"ee",
         12531 => x"56",
         12532 => x"08",
         12533 => x"bb",
         12534 => x"18",
         12535 => x"08",
         12536 => x"31",
         12537 => x"18",
         12538 => x"ee",
         12539 => x"33",
         12540 => x"2e",
         12541 => x"fe",
         12542 => x"54",
         12543 => x"a0",
         12544 => x"53",
         12545 => x"17",
         12546 => x"ee",
         12547 => x"ca",
         12548 => x"7b",
         12549 => x"55",
         12550 => x"fd",
         12551 => x"9c",
         12552 => x"fd",
         12553 => x"52",
         12554 => x"f3",
         12555 => x"bb",
         12556 => x"84",
         12557 => x"80",
         12558 => x"38",
         12559 => x"08",
         12560 => x"8d",
         12561 => x"84",
         12562 => x"fd",
         12563 => x"53",
         12564 => x"51",
         12565 => x"3f",
         12566 => x"08",
         12567 => x"9c",
         12568 => x"11",
         12569 => x"5a",
         12570 => x"7b",
         12571 => x"81",
         12572 => x"0c",
         12573 => x"81",
         12574 => x"84",
         12575 => x"55",
         12576 => x"ff",
         12577 => x"84",
         12578 => x"9f",
         12579 => x"8a",
         12580 => x"74",
         12581 => x"06",
         12582 => x"76",
         12583 => x"81",
         12584 => x"38",
         12585 => x"1f",
         12586 => x"75",
         12587 => x"57",
         12588 => x"56",
         12589 => x"7d",
         12590 => x"b8",
         12591 => x"58",
         12592 => x"c3",
         12593 => x"59",
         12594 => x"1a",
         12595 => x"cf",
         12596 => x"0b",
         12597 => x"34",
         12598 => x"80",
         12599 => x"7d",
         12600 => x"ff",
         12601 => x"77",
         12602 => x"34",
         12603 => x"5b",
         12604 => x"17",
         12605 => x"55",
         12606 => x"81",
         12607 => x"59",
         12608 => x"d8",
         12609 => x"57",
         12610 => x"70",
         12611 => x"33",
         12612 => x"05",
         12613 => x"16",
         12614 => x"38",
         12615 => x"0b",
         12616 => x"34",
         12617 => x"83",
         12618 => x"5b",
         12619 => x"80",
         12620 => x"78",
         12621 => x"7a",
         12622 => x"34",
         12623 => x"74",
         12624 => x"f0",
         12625 => x"81",
         12626 => x"34",
         12627 => x"92",
         12628 => x"bb",
         12629 => x"84",
         12630 => x"fd",
         12631 => x"56",
         12632 => x"08",
         12633 => x"84",
         12634 => x"97",
         12635 => x"0b",
         12636 => x"80",
         12637 => x"17",
         12638 => x"58",
         12639 => x"18",
         12640 => x"2a",
         12641 => x"18",
         12642 => x"5a",
         12643 => x"80",
         12644 => x"55",
         12645 => x"16",
         12646 => x"81",
         12647 => x"34",
         12648 => x"ed",
         12649 => x"bb",
         12650 => x"75",
         12651 => x"0c",
         12652 => x"04",
         12653 => x"55",
         12654 => x"17",
         12655 => x"2a",
         12656 => x"ed",
         12657 => x"fd",
         12658 => x"2a",
         12659 => x"cc",
         12660 => x"88",
         12661 => x"80",
         12662 => x"7d",
         12663 => x"80",
         12664 => x"1b",
         12665 => x"fe",
         12666 => x"90",
         12667 => x"94",
         12668 => x"88",
         12669 => x"95",
         12670 => x"55",
         12671 => x"16",
         12672 => x"81",
         12673 => x"34",
         12674 => x"ec",
         12675 => x"bb",
         12676 => x"ff",
         12677 => x"3d",
         12678 => x"b4",
         12679 => x"59",
         12680 => x"80",
         12681 => x"79",
         12682 => x"5b",
         12683 => x"26",
         12684 => x"ba",
         12685 => x"38",
         12686 => x"75",
         12687 => x"af",
         12688 => x"b1",
         12689 => x"05",
         12690 => x"51",
         12691 => x"3f",
         12692 => x"08",
         12693 => x"84",
         12694 => x"8a",
         12695 => x"bb",
         12696 => x"3d",
         12697 => x"a6",
         12698 => x"3d",
         12699 => x"3d",
         12700 => x"ff",
         12701 => x"84",
         12702 => x"56",
         12703 => x"08",
         12704 => x"81",
         12705 => x"81",
         12706 => x"86",
         12707 => x"38",
         12708 => x"3d",
         12709 => x"58",
         12710 => x"70",
         12711 => x"33",
         12712 => x"05",
         12713 => x"15",
         12714 => x"38",
         12715 => x"b0",
         12716 => x"58",
         12717 => x"81",
         12718 => x"77",
         12719 => x"59",
         12720 => x"55",
         12721 => x"b3",
         12722 => x"77",
         12723 => x"8e",
         12724 => x"84",
         12725 => x"bb",
         12726 => x"d8",
         12727 => x"3d",
         12728 => x"cb",
         12729 => x"84",
         12730 => x"b1",
         12731 => x"76",
         12732 => x"70",
         12733 => x"57",
         12734 => x"89",
         12735 => x"82",
         12736 => x"ff",
         12737 => x"5d",
         12738 => x"2e",
         12739 => x"80",
         12740 => x"e6",
         12741 => x"72",
         12742 => x"5f",
         12743 => x"81",
         12744 => x"79",
         12745 => x"5b",
         12746 => x"12",
         12747 => x"77",
         12748 => x"38",
         12749 => x"81",
         12750 => x"55",
         12751 => x"58",
         12752 => x"89",
         12753 => x"70",
         12754 => x"58",
         12755 => x"70",
         12756 => x"55",
         12757 => x"09",
         12758 => x"38",
         12759 => x"38",
         12760 => x"70",
         12761 => x"07",
         12762 => x"07",
         12763 => x"7a",
         12764 => x"38",
         12765 => x"1e",
         12766 => x"83",
         12767 => x"38",
         12768 => x"5a",
         12769 => x"39",
         12770 => x"fd",
         12771 => x"7f",
         12772 => x"b1",
         12773 => x"05",
         12774 => x"51",
         12775 => x"3f",
         12776 => x"08",
         12777 => x"84",
         12778 => x"38",
         12779 => x"6c",
         12780 => x"2e",
         12781 => x"fe",
         12782 => x"51",
         12783 => x"3f",
         12784 => x"08",
         12785 => x"84",
         12786 => x"38",
         12787 => x"0b",
         12788 => x"88",
         12789 => x"05",
         12790 => x"75",
         12791 => x"57",
         12792 => x"81",
         12793 => x"ff",
         12794 => x"ef",
         12795 => x"cb",
         12796 => x"19",
         12797 => x"33",
         12798 => x"81",
         12799 => x"7e",
         12800 => x"a0",
         12801 => x"8b",
         12802 => x"5d",
         12803 => x"1e",
         12804 => x"33",
         12805 => x"81",
         12806 => x"75",
         12807 => x"c5",
         12808 => x"08",
         12809 => x"bd",
         12810 => x"19",
         12811 => x"33",
         12812 => x"07",
         12813 => x"58",
         12814 => x"83",
         12815 => x"38",
         12816 => x"18",
         12817 => x"5e",
         12818 => x"27",
         12819 => x"8a",
         12820 => x"71",
         12821 => x"08",
         12822 => x"75",
         12823 => x"b5",
         12824 => x"5d",
         12825 => x"08",
         12826 => x"38",
         12827 => x"5f",
         12828 => x"38",
         12829 => x"53",
         12830 => x"81",
         12831 => x"fe",
         12832 => x"84",
         12833 => x"80",
         12834 => x"ff",
         12835 => x"77",
         12836 => x"7f",
         12837 => x"d8",
         12838 => x"7b",
         12839 => x"81",
         12840 => x"79",
         12841 => x"81",
         12842 => x"6a",
         12843 => x"ff",
         12844 => x"7b",
         12845 => x"34",
         12846 => x"58",
         12847 => x"18",
         12848 => x"5b",
         12849 => x"09",
         12850 => x"38",
         12851 => x"5e",
         12852 => x"18",
         12853 => x"2a",
         12854 => x"ed",
         12855 => x"57",
         12856 => x"18",
         12857 => x"aa",
         12858 => x"3d",
         12859 => x"56",
         12860 => x"95",
         12861 => x"78",
         12862 => x"db",
         12863 => x"84",
         12864 => x"bb",
         12865 => x"f5",
         12866 => x"5c",
         12867 => x"57",
         12868 => x"16",
         12869 => x"b4",
         12870 => x"33",
         12871 => x"7e",
         12872 => x"81",
         12873 => x"38",
         12874 => x"53",
         12875 => x"81",
         12876 => x"fe",
         12877 => x"84",
         12878 => x"80",
         12879 => x"ff",
         12880 => x"76",
         12881 => x"77",
         12882 => x"38",
         12883 => x"5a",
         12884 => x"81",
         12885 => x"34",
         12886 => x"7b",
         12887 => x"80",
         12888 => x"fe",
         12889 => x"84",
         12890 => x"55",
         12891 => x"08",
         12892 => x"98",
         12893 => x"74",
         12894 => x"e1",
         12895 => x"74",
         12896 => x"7f",
         12897 => x"d6",
         12898 => x"84",
         12899 => x"84",
         12900 => x"0d",
         12901 => x"84",
         12902 => x"b1",
         12903 => x"95",
         12904 => x"19",
         12905 => x"2b",
         12906 => x"07",
         12907 => x"56",
         12908 => x"39",
         12909 => x"08",
         12910 => x"fe",
         12911 => x"84",
         12912 => x"fe",
         12913 => x"84",
         12914 => x"b1",
         12915 => x"81",
         12916 => x"08",
         12917 => x"81",
         12918 => x"fe",
         12919 => x"81",
         12920 => x"84",
         12921 => x"09",
         12922 => x"db",
         12923 => x"84",
         12924 => x"34",
         12925 => x"a8",
         12926 => x"84",
         12927 => x"59",
         12928 => x"17",
         12929 => x"a0",
         12930 => x"33",
         12931 => x"2e",
         12932 => x"fe",
         12933 => x"54",
         12934 => x"a0",
         12935 => x"53",
         12936 => x"16",
         12937 => x"e2",
         12938 => x"58",
         12939 => x"81",
         12940 => x"08",
         12941 => x"70",
         12942 => x"33",
         12943 => x"e1",
         12944 => x"5c",
         12945 => x"08",
         12946 => x"84",
         12947 => x"83",
         12948 => x"17",
         12949 => x"08",
         12950 => x"84",
         12951 => x"74",
         12952 => x"27",
         12953 => x"82",
         12954 => x"7c",
         12955 => x"81",
         12956 => x"38",
         12957 => x"17",
         12958 => x"08",
         12959 => x"52",
         12960 => x"51",
         12961 => x"3f",
         12962 => x"e8",
         12963 => x"0d",
         12964 => x"05",
         12965 => x"05",
         12966 => x"33",
         12967 => x"53",
         12968 => x"05",
         12969 => x"51",
         12970 => x"3f",
         12971 => x"08",
         12972 => x"84",
         12973 => x"8a",
         12974 => x"bb",
         12975 => x"3d",
         12976 => x"5a",
         12977 => x"3d",
         12978 => x"ff",
         12979 => x"84",
         12980 => x"56",
         12981 => x"08",
         12982 => x"80",
         12983 => x"81",
         12984 => x"86",
         12985 => x"38",
         12986 => x"61",
         12987 => x"12",
         12988 => x"7a",
         12989 => x"51",
         12990 => x"73",
         12991 => x"78",
         12992 => x"83",
         12993 => x"51",
         12994 => x"3f",
         12995 => x"08",
         12996 => x"0c",
         12997 => x"04",
         12998 => x"67",
         12999 => x"96",
         13000 => x"52",
         13001 => x"ff",
         13002 => x"84",
         13003 => x"55",
         13004 => x"08",
         13005 => x"38",
         13006 => x"84",
         13007 => x"0d",
         13008 => x"66",
         13009 => x"d0",
         13010 => x"96",
         13011 => x"bb",
         13012 => x"84",
         13013 => x"e0",
         13014 => x"cf",
         13015 => x"a0",
         13016 => x"55",
         13017 => x"60",
         13018 => x"86",
         13019 => x"90",
         13020 => x"59",
         13021 => x"17",
         13022 => x"2a",
         13023 => x"17",
         13024 => x"2a",
         13025 => x"17",
         13026 => x"2a",
         13027 => x"17",
         13028 => x"81",
         13029 => x"34",
         13030 => x"e1",
         13031 => x"bb",
         13032 => x"bb",
         13033 => x"3d",
         13034 => x"3d",
         13035 => x"5d",
         13036 => x"9a",
         13037 => x"52",
         13038 => x"ff",
         13039 => x"84",
         13040 => x"84",
         13041 => x"30",
         13042 => x"84",
         13043 => x"25",
         13044 => x"7a",
         13045 => x"38",
         13046 => x"06",
         13047 => x"81",
         13048 => x"30",
         13049 => x"80",
         13050 => x"7b",
         13051 => x"8c",
         13052 => x"76",
         13053 => x"78",
         13054 => x"80",
         13055 => x"11",
         13056 => x"80",
         13057 => x"08",
         13058 => x"f6",
         13059 => x"33",
         13060 => x"74",
         13061 => x"81",
         13062 => x"38",
         13063 => x"53",
         13064 => x"81",
         13065 => x"fe",
         13066 => x"84",
         13067 => x"80",
         13068 => x"ff",
         13069 => x"76",
         13070 => x"78",
         13071 => x"38",
         13072 => x"56",
         13073 => x"56",
         13074 => x"8b",
         13075 => x"56",
         13076 => x"83",
         13077 => x"75",
         13078 => x"83",
         13079 => x"12",
         13080 => x"2b",
         13081 => x"07",
         13082 => x"70",
         13083 => x"2b",
         13084 => x"07",
         13085 => x"5d",
         13086 => x"56",
         13087 => x"84",
         13088 => x"0d",
         13089 => x"80",
         13090 => x"8e",
         13091 => x"55",
         13092 => x"3f",
         13093 => x"08",
         13094 => x"84",
         13095 => x"81",
         13096 => x"84",
         13097 => x"06",
         13098 => x"80",
         13099 => x"57",
         13100 => x"77",
         13101 => x"08",
         13102 => x"70",
         13103 => x"33",
         13104 => x"dc",
         13105 => x"59",
         13106 => x"08",
         13107 => x"81",
         13108 => x"38",
         13109 => x"08",
         13110 => x"b4",
         13111 => x"17",
         13112 => x"bb",
         13113 => x"55",
         13114 => x"08",
         13115 => x"38",
         13116 => x"55",
         13117 => x"09",
         13118 => x"a0",
         13119 => x"b4",
         13120 => x"17",
         13121 => x"7a",
         13122 => x"33",
         13123 => x"9b",
         13124 => x"81",
         13125 => x"b8",
         13126 => x"16",
         13127 => x"db",
         13128 => x"bb",
         13129 => x"2e",
         13130 => x"fe",
         13131 => x"52",
         13132 => x"f8",
         13133 => x"bb",
         13134 => x"84",
         13135 => x"fe",
         13136 => x"bb",
         13137 => x"bb",
         13138 => x"5c",
         13139 => x"18",
         13140 => x"1b",
         13141 => x"75",
         13142 => x"81",
         13143 => x"78",
         13144 => x"8b",
         13145 => x"58",
         13146 => x"77",
         13147 => x"f2",
         13148 => x"7b",
         13149 => x"5c",
         13150 => x"a0",
         13151 => x"fc",
         13152 => x"57",
         13153 => x"e1",
         13154 => x"53",
         13155 => x"b4",
         13156 => x"3d",
         13157 => x"a4",
         13158 => x"84",
         13159 => x"bb",
         13160 => x"a6",
         13161 => x"5d",
         13162 => x"55",
         13163 => x"81",
         13164 => x"ff",
         13165 => x"f4",
         13166 => x"3d",
         13167 => x"70",
         13168 => x"5b",
         13169 => x"9f",
         13170 => x"b7",
         13171 => x"90",
         13172 => x"75",
         13173 => x"81",
         13174 => x"74",
         13175 => x"75",
         13176 => x"83",
         13177 => x"81",
         13178 => x"51",
         13179 => x"83",
         13180 => x"bb",
         13181 => x"9f",
         13182 => x"bb",
         13183 => x"ff",
         13184 => x"76",
         13185 => x"e0",
         13186 => x"94",
         13187 => x"94",
         13188 => x"ff",
         13189 => x"58",
         13190 => x"81",
         13191 => x"56",
         13192 => x"99",
         13193 => x"70",
         13194 => x"ff",
         13195 => x"58",
         13196 => x"89",
         13197 => x"2e",
         13198 => x"e9",
         13199 => x"ff",
         13200 => x"81",
         13201 => x"ff",
         13202 => x"f8",
         13203 => x"26",
         13204 => x"81",
         13205 => x"8f",
         13206 => x"2a",
         13207 => x"70",
         13208 => x"34",
         13209 => x"76",
         13210 => x"05",
         13211 => x"1a",
         13212 => x"70",
         13213 => x"ff",
         13214 => x"58",
         13215 => x"26",
         13216 => x"8f",
         13217 => x"86",
         13218 => x"e5",
         13219 => x"79",
         13220 => x"38",
         13221 => x"56",
         13222 => x"33",
         13223 => x"a0",
         13224 => x"06",
         13225 => x"1a",
         13226 => x"38",
         13227 => x"47",
         13228 => x"3d",
         13229 => x"fe",
         13230 => x"84",
         13231 => x"55",
         13232 => x"08",
         13233 => x"38",
         13234 => x"84",
         13235 => x"a1",
         13236 => x"83",
         13237 => x"51",
         13238 => x"84",
         13239 => x"83",
         13240 => x"55",
         13241 => x"38",
         13242 => x"84",
         13243 => x"a1",
         13244 => x"83",
         13245 => x"56",
         13246 => x"81",
         13247 => x"fe",
         13248 => x"84",
         13249 => x"55",
         13250 => x"08",
         13251 => x"79",
         13252 => x"c4",
         13253 => x"7e",
         13254 => x"76",
         13255 => x"58",
         13256 => x"81",
         13257 => x"ff",
         13258 => x"ef",
         13259 => x"81",
         13260 => x"34",
         13261 => x"da",
         13262 => x"bb",
         13263 => x"74",
         13264 => x"39",
         13265 => x"fe",
         13266 => x"56",
         13267 => x"84",
         13268 => x"84",
         13269 => x"06",
         13270 => x"80",
         13271 => x"2e",
         13272 => x"75",
         13273 => x"76",
         13274 => x"ee",
         13275 => x"bb",
         13276 => x"84",
         13277 => x"75",
         13278 => x"06",
         13279 => x"84",
         13280 => x"b8",
         13281 => x"98",
         13282 => x"80",
         13283 => x"08",
         13284 => x"38",
         13285 => x"55",
         13286 => x"09",
         13287 => x"d7",
         13288 => x"76",
         13289 => x"52",
         13290 => x"51",
         13291 => x"3f",
         13292 => x"08",
         13293 => x"38",
         13294 => x"59",
         13295 => x"0c",
         13296 => x"be",
         13297 => x"17",
         13298 => x"57",
         13299 => x"81",
         13300 => x"9e",
         13301 => x"70",
         13302 => x"07",
         13303 => x"80",
         13304 => x"38",
         13305 => x"79",
         13306 => x"38",
         13307 => x"51",
         13308 => x"3f",
         13309 => x"08",
         13310 => x"84",
         13311 => x"ff",
         13312 => x"55",
         13313 => x"fd",
         13314 => x"55",
         13315 => x"38",
         13316 => x"55",
         13317 => x"81",
         13318 => x"ff",
         13319 => x"f4",
         13320 => x"88",
         13321 => x"34",
         13322 => x"59",
         13323 => x"70",
         13324 => x"33",
         13325 => x"05",
         13326 => x"15",
         13327 => x"2e",
         13328 => x"76",
         13329 => x"58",
         13330 => x"81",
         13331 => x"ff",
         13332 => x"da",
         13333 => x"39",
         13334 => x"7a",
         13335 => x"81",
         13336 => x"34",
         13337 => x"d7",
         13338 => x"bb",
         13339 => x"fd",
         13340 => x"57",
         13341 => x"81",
         13342 => x"08",
         13343 => x"81",
         13344 => x"fe",
         13345 => x"84",
         13346 => x"79",
         13347 => x"06",
         13348 => x"84",
         13349 => x"83",
         13350 => x"18",
         13351 => x"08",
         13352 => x"a0",
         13353 => x"8a",
         13354 => x"33",
         13355 => x"2e",
         13356 => x"bb",
         13357 => x"fd",
         13358 => x"5a",
         13359 => x"51",
         13360 => x"3f",
         13361 => x"08",
         13362 => x"84",
         13363 => x"fd",
         13364 => x"ae",
         13365 => x"58",
         13366 => x"2e",
         13367 => x"fe",
         13368 => x"54",
         13369 => x"a0",
         13370 => x"53",
         13371 => x"18",
         13372 => x"d4",
         13373 => x"a9",
         13374 => x"0d",
         13375 => x"88",
         13376 => x"05",
         13377 => x"57",
         13378 => x"80",
         13379 => x"76",
         13380 => x"80",
         13381 => x"74",
         13382 => x"80",
         13383 => x"86",
         13384 => x"18",
         13385 => x"78",
         13386 => x"c2",
         13387 => x"73",
         13388 => x"a5",
         13389 => x"33",
         13390 => x"9d",
         13391 => x"2e",
         13392 => x"8c",
         13393 => x"9c",
         13394 => x"33",
         13395 => x"81",
         13396 => x"74",
         13397 => x"8c",
         13398 => x"11",
         13399 => x"2b",
         13400 => x"54",
         13401 => x"fd",
         13402 => x"ff",
         13403 => x"70",
         13404 => x"07",
         13405 => x"bb",
         13406 => x"90",
         13407 => x"42",
         13408 => x"58",
         13409 => x"88",
         13410 => x"08",
         13411 => x"38",
         13412 => x"78",
         13413 => x"59",
         13414 => x"51",
         13415 => x"3f",
         13416 => x"55",
         13417 => x"08",
         13418 => x"38",
         13419 => x"bb",
         13420 => x"2e",
         13421 => x"84",
         13422 => x"ff",
         13423 => x"38",
         13424 => x"08",
         13425 => x"81",
         13426 => x"7d",
         13427 => x"74",
         13428 => x"81",
         13429 => x"87",
         13430 => x"73",
         13431 => x"0c",
         13432 => x"04",
         13433 => x"bb",
         13434 => x"3d",
         13435 => x"15",
         13436 => x"d0",
         13437 => x"bb",
         13438 => x"06",
         13439 => x"ad",
         13440 => x"08",
         13441 => x"a7",
         13442 => x"2e",
         13443 => x"7a",
         13444 => x"7c",
         13445 => x"38",
         13446 => x"74",
         13447 => x"e6",
         13448 => x"77",
         13449 => x"fe",
         13450 => x"84",
         13451 => x"56",
         13452 => x"08",
         13453 => x"77",
         13454 => x"17",
         13455 => x"74",
         13456 => x"7e",
         13457 => x"55",
         13458 => x"ff",
         13459 => x"88",
         13460 => x"8c",
         13461 => x"17",
         13462 => x"07",
         13463 => x"18",
         13464 => x"08",
         13465 => x"16",
         13466 => x"76",
         13467 => x"e9",
         13468 => x"31",
         13469 => x"84",
         13470 => x"07",
         13471 => x"16",
         13472 => x"fe",
         13473 => x"54",
         13474 => x"74",
         13475 => x"fe",
         13476 => x"54",
         13477 => x"81",
         13478 => x"39",
         13479 => x"ff",
         13480 => x"bb",
         13481 => x"3d",
         13482 => x"08",
         13483 => x"02",
         13484 => x"87",
         13485 => x"42",
         13486 => x"a2",
         13487 => x"5f",
         13488 => x"80",
         13489 => x"38",
         13490 => x"05",
         13491 => x"9f",
         13492 => x"75",
         13493 => x"9b",
         13494 => x"38",
         13495 => x"85",
         13496 => x"e2",
         13497 => x"80",
         13498 => x"e5",
         13499 => x"10",
         13500 => x"05",
         13501 => x"5a",
         13502 => x"84",
         13503 => x"34",
         13504 => x"ba",
         13505 => x"84",
         13506 => x"33",
         13507 => x"81",
         13508 => x"fe",
         13509 => x"84",
         13510 => x"81",
         13511 => x"81",
         13512 => x"83",
         13513 => x"ab",
         13514 => x"2a",
         13515 => x"8a",
         13516 => x"9f",
         13517 => x"fc",
         13518 => x"52",
         13519 => x"d0",
         13520 => x"bb",
         13521 => x"98",
         13522 => x"74",
         13523 => x"90",
         13524 => x"80",
         13525 => x"88",
         13526 => x"75",
         13527 => x"83",
         13528 => x"80",
         13529 => x"84",
         13530 => x"83",
         13531 => x"81",
         13532 => x"83",
         13533 => x"1f",
         13534 => x"74",
         13535 => x"7e",
         13536 => x"3d",
         13537 => x"70",
         13538 => x"59",
         13539 => x"60",
         13540 => x"ab",
         13541 => x"70",
         13542 => x"07",
         13543 => x"57",
         13544 => x"38",
         13545 => x"84",
         13546 => x"54",
         13547 => x"52",
         13548 => x"cd",
         13549 => x"57",
         13550 => x"08",
         13551 => x"60",
         13552 => x"33",
         13553 => x"05",
         13554 => x"2b",
         13555 => x"8e",
         13556 => x"d4",
         13557 => x"81",
         13558 => x"38",
         13559 => x"61",
         13560 => x"11",
         13561 => x"62",
         13562 => x"e7",
         13563 => x"18",
         13564 => x"82",
         13565 => x"90",
         13566 => x"2b",
         13567 => x"33",
         13568 => x"88",
         13569 => x"71",
         13570 => x"1f",
         13571 => x"82",
         13572 => x"90",
         13573 => x"2b",
         13574 => x"33",
         13575 => x"88",
         13576 => x"71",
         13577 => x"3d",
         13578 => x"3d",
         13579 => x"0c",
         13580 => x"45",
         13581 => x"5a",
         13582 => x"8e",
         13583 => x"79",
         13584 => x"38",
         13585 => x"81",
         13586 => x"87",
         13587 => x"2a",
         13588 => x"45",
         13589 => x"2e",
         13590 => x"61",
         13591 => x"64",
         13592 => x"38",
         13593 => x"47",
         13594 => x"38",
         13595 => x"30",
         13596 => x"7a",
         13597 => x"2e",
         13598 => x"7a",
         13599 => x"8c",
         13600 => x"0b",
         13601 => x"22",
         13602 => x"80",
         13603 => x"74",
         13604 => x"38",
         13605 => x"56",
         13606 => x"17",
         13607 => x"57",
         13608 => x"2e",
         13609 => x"75",
         13610 => x"77",
         13611 => x"fc",
         13612 => x"84",
         13613 => x"10",
         13614 => x"84",
         13615 => x"9f",
         13616 => x"38",
         13617 => x"bb",
         13618 => x"84",
         13619 => x"05",
         13620 => x"2a",
         13621 => x"4c",
         13622 => x"15",
         13623 => x"81",
         13624 => x"7b",
         13625 => x"68",
         13626 => x"ff",
         13627 => x"06",
         13628 => x"4e",
         13629 => x"83",
         13630 => x"38",
         13631 => x"77",
         13632 => x"70",
         13633 => x"57",
         13634 => x"82",
         13635 => x"7c",
         13636 => x"78",
         13637 => x"31",
         13638 => x"ff",
         13639 => x"bb",
         13640 => x"62",
         13641 => x"f6",
         13642 => x"2e",
         13643 => x"82",
         13644 => x"ff",
         13645 => x"bb",
         13646 => x"82",
         13647 => x"89",
         13648 => x"18",
         13649 => x"c0",
         13650 => x"38",
         13651 => x"a3",
         13652 => x"76",
         13653 => x"0c",
         13654 => x"84",
         13655 => x"04",
         13656 => x"fe",
         13657 => x"84",
         13658 => x"9f",
         13659 => x"bb",
         13660 => x"7c",
         13661 => x"70",
         13662 => x"57",
         13663 => x"89",
         13664 => x"82",
         13665 => x"ff",
         13666 => x"5d",
         13667 => x"2e",
         13668 => x"80",
         13669 => x"f4",
         13670 => x"08",
         13671 => x"7a",
         13672 => x"5c",
         13673 => x"81",
         13674 => x"ff",
         13675 => x"59",
         13676 => x"26",
         13677 => x"17",
         13678 => x"06",
         13679 => x"9f",
         13680 => x"99",
         13681 => x"e0",
         13682 => x"ff",
         13683 => x"76",
         13684 => x"2a",
         13685 => x"78",
         13686 => x"06",
         13687 => x"ff",
         13688 => x"7a",
         13689 => x"70",
         13690 => x"2a",
         13691 => x"4a",
         13692 => x"2e",
         13693 => x"81",
         13694 => x"5f",
         13695 => x"25",
         13696 => x"7f",
         13697 => x"39",
         13698 => x"05",
         13699 => x"79",
         13700 => x"96",
         13701 => x"84",
         13702 => x"fe",
         13703 => x"83",
         13704 => x"84",
         13705 => x"40",
         13706 => x"38",
         13707 => x"55",
         13708 => x"75",
         13709 => x"38",
         13710 => x"59",
         13711 => x"81",
         13712 => x"39",
         13713 => x"ff",
         13714 => x"7a",
         13715 => x"56",
         13716 => x"61",
         13717 => x"93",
         13718 => x"2e",
         13719 => x"82",
         13720 => x"4a",
         13721 => x"8b",
         13722 => x"84",
         13723 => x"26",
         13724 => x"8b",
         13725 => x"5b",
         13726 => x"27",
         13727 => x"8e",
         13728 => x"bb",
         13729 => x"3d",
         13730 => x"90",
         13731 => x"55",
         13732 => x"86",
         13733 => x"f5",
         13734 => x"38",
         13735 => x"5b",
         13736 => x"fd",
         13737 => x"80",
         13738 => x"80",
         13739 => x"05",
         13740 => x"15",
         13741 => x"38",
         13742 => x"e6",
         13743 => x"55",
         13744 => x"05",
         13745 => x"70",
         13746 => x"34",
         13747 => x"74",
         13748 => x"8b",
         13749 => x"65",
         13750 => x"8c",
         13751 => x"61",
         13752 => x"7b",
         13753 => x"06",
         13754 => x"8e",
         13755 => x"88",
         13756 => x"61",
         13757 => x"81",
         13758 => x"34",
         13759 => x"70",
         13760 => x"80",
         13761 => x"34",
         13762 => x"82",
         13763 => x"61",
         13764 => x"6c",
         13765 => x"ff",
         13766 => x"ad",
         13767 => x"ff",
         13768 => x"74",
         13769 => x"34",
         13770 => x"4c",
         13771 => x"05",
         13772 => x"95",
         13773 => x"61",
         13774 => x"80",
         13775 => x"34",
         13776 => x"05",
         13777 => x"9b",
         13778 => x"61",
         13779 => x"7e",
         13780 => x"67",
         13781 => x"34",
         13782 => x"4c",
         13783 => x"05",
         13784 => x"2a",
         13785 => x"0c",
         13786 => x"08",
         13787 => x"34",
         13788 => x"85",
         13789 => x"61",
         13790 => x"80",
         13791 => x"34",
         13792 => x"05",
         13793 => x"61",
         13794 => x"7c",
         13795 => x"06",
         13796 => x"96",
         13797 => x"88",
         13798 => x"61",
         13799 => x"ff",
         13800 => x"05",
         13801 => x"a6",
         13802 => x"61",
         13803 => x"e6",
         13804 => x"55",
         13805 => x"05",
         13806 => x"70",
         13807 => x"34",
         13808 => x"74",
         13809 => x"83",
         13810 => x"80",
         13811 => x"60",
         13812 => x"4b",
         13813 => x"34",
         13814 => x"53",
         13815 => x"51",
         13816 => x"3f",
         13817 => x"bb",
         13818 => x"e7",
         13819 => x"5c",
         13820 => x"87",
         13821 => x"61",
         13822 => x"76",
         13823 => x"58",
         13824 => x"55",
         13825 => x"63",
         13826 => x"62",
         13827 => x"c0",
         13828 => x"ff",
         13829 => x"81",
         13830 => x"f8",
         13831 => x"34",
         13832 => x"7c",
         13833 => x"64",
         13834 => x"46",
         13835 => x"2a",
         13836 => x"70",
         13837 => x"34",
         13838 => x"56",
         13839 => x"7c",
         13840 => x"76",
         13841 => x"38",
         13842 => x"54",
         13843 => x"52",
         13844 => x"c5",
         13845 => x"bb",
         13846 => x"e6",
         13847 => x"61",
         13848 => x"76",
         13849 => x"58",
         13850 => x"55",
         13851 => x"78",
         13852 => x"31",
         13853 => x"c9",
         13854 => x"05",
         13855 => x"2e",
         13856 => x"77",
         13857 => x"2e",
         13858 => x"56",
         13859 => x"66",
         13860 => x"75",
         13861 => x"7a",
         13862 => x"79",
         13863 => x"8b",
         13864 => x"84",
         13865 => x"38",
         13866 => x"76",
         13867 => x"75",
         13868 => x"58",
         13869 => x"93",
         13870 => x"6c",
         13871 => x"26",
         13872 => x"58",
         13873 => x"83",
         13874 => x"7d",
         13875 => x"61",
         13876 => x"06",
         13877 => x"b3",
         13878 => x"61",
         13879 => x"75",
         13880 => x"57",
         13881 => x"59",
         13882 => x"80",
         13883 => x"ff",
         13884 => x"60",
         13885 => x"47",
         13886 => x"81",
         13887 => x"34",
         13888 => x"05",
         13889 => x"83",
         13890 => x"67",
         13891 => x"6c",
         13892 => x"c1",
         13893 => x"51",
         13894 => x"3f",
         13895 => x"05",
         13896 => x"84",
         13897 => x"bf",
         13898 => x"67",
         13899 => x"84",
         13900 => x"67",
         13901 => x"7e",
         13902 => x"05",
         13903 => x"83",
         13904 => x"6b",
         13905 => x"05",
         13906 => x"90",
         13907 => x"c9",
         13908 => x"61",
         13909 => x"34",
         13910 => x"45",
         13911 => x"cb",
         13912 => x"90",
         13913 => x"61",
         13914 => x"34",
         13915 => x"5f",
         13916 => x"cd",
         13917 => x"54",
         13918 => x"52",
         13919 => x"c3",
         13920 => x"57",
         13921 => x"08",
         13922 => x"80",
         13923 => x"79",
         13924 => x"96",
         13925 => x"84",
         13926 => x"f7",
         13927 => x"bb",
         13928 => x"bb",
         13929 => x"3d",
         13930 => x"90",
         13931 => x"55",
         13932 => x"74",
         13933 => x"45",
         13934 => x"39",
         13935 => x"78",
         13936 => x"81",
         13937 => x"b8",
         13938 => x"74",
         13939 => x"38",
         13940 => x"98",
         13941 => x"b8",
         13942 => x"82",
         13943 => x"57",
         13944 => x"80",
         13945 => x"76",
         13946 => x"38",
         13947 => x"51",
         13948 => x"3f",
         13949 => x"08",
         13950 => x"87",
         13951 => x"2a",
         13952 => x"5c",
         13953 => x"bb",
         13954 => x"80",
         13955 => x"47",
         13956 => x"0a",
         13957 => x"cb",
         13958 => x"f8",
         13959 => x"bb",
         13960 => x"ff",
         13961 => x"e6",
         13962 => x"d3",
         13963 => x"2a",
         13964 => x"bf",
         13965 => x"f8",
         13966 => x"81",
         13967 => x"80",
         13968 => x"38",
         13969 => x"ab",
         13970 => x"a0",
         13971 => x"88",
         13972 => x"61",
         13973 => x"75",
         13974 => x"7a",
         13975 => x"34",
         13976 => x"57",
         13977 => x"05",
         13978 => x"39",
         13979 => x"c3",
         13980 => x"61",
         13981 => x"34",
         13982 => x"c5",
         13983 => x"cc",
         13984 => x"05",
         13985 => x"a4",
         13986 => x"88",
         13987 => x"61",
         13988 => x"7c",
         13989 => x"78",
         13990 => x"34",
         13991 => x"56",
         13992 => x"05",
         13993 => x"ac",
         13994 => x"61",
         13995 => x"80",
         13996 => x"34",
         13997 => x"05",
         13998 => x"b0",
         13999 => x"61",
         14000 => x"86",
         14001 => x"34",
         14002 => x"05",
         14003 => x"61",
         14004 => x"34",
         14005 => x"c2",
         14006 => x"61",
         14007 => x"83",
         14008 => x"57",
         14009 => x"81",
         14010 => x"76",
         14011 => x"58",
         14012 => x"55",
         14013 => x"f9",
         14014 => x"70",
         14015 => x"33",
         14016 => x"05",
         14017 => x"15",
         14018 => x"38",
         14019 => x"81",
         14020 => x"60",
         14021 => x"fe",
         14022 => x"81",
         14023 => x"84",
         14024 => x"38",
         14025 => x"61",
         14026 => x"62",
         14027 => x"34",
         14028 => x"bb",
         14029 => x"60",
         14030 => x"fe",
         14031 => x"fc",
         14032 => x"0b",
         14033 => x"0c",
         14034 => x"84",
         14035 => x"04",
         14036 => x"7b",
         14037 => x"70",
         14038 => x"34",
         14039 => x"81",
         14040 => x"ff",
         14041 => x"61",
         14042 => x"ff",
         14043 => x"34",
         14044 => x"05",
         14045 => x"87",
         14046 => x"61",
         14047 => x"ff",
         14048 => x"34",
         14049 => x"05",
         14050 => x"34",
         14051 => x"b1",
         14052 => x"86",
         14053 => x"52",
         14054 => x"bf",
         14055 => x"80",
         14056 => x"80",
         14057 => x"05",
         14058 => x"17",
         14059 => x"38",
         14060 => x"d2",
         14061 => x"05",
         14062 => x"55",
         14063 => x"70",
         14064 => x"34",
         14065 => x"70",
         14066 => x"34",
         14067 => x"34",
         14068 => x"83",
         14069 => x"80",
         14070 => x"e5",
         14071 => x"c1",
         14072 => x"05",
         14073 => x"61",
         14074 => x"34",
         14075 => x"5b",
         14076 => x"e8",
         14077 => x"88",
         14078 => x"61",
         14079 => x"34",
         14080 => x"56",
         14081 => x"ea",
         14082 => x"98",
         14083 => x"61",
         14084 => x"34",
         14085 => x"ec",
         14086 => x"61",
         14087 => x"34",
         14088 => x"ee",
         14089 => x"61",
         14090 => x"34",
         14091 => x"34",
         14092 => x"34",
         14093 => x"1f",
         14094 => x"79",
         14095 => x"eb",
         14096 => x"81",
         14097 => x"52",
         14098 => x"bd",
         14099 => x"61",
         14100 => x"a6",
         14101 => x"0d",
         14102 => x"5b",
         14103 => x"ff",
         14104 => x"57",
         14105 => x"b8",
         14106 => x"59",
         14107 => x"05",
         14108 => x"78",
         14109 => x"ff",
         14110 => x"7b",
         14111 => x"81",
         14112 => x"8d",
         14113 => x"74",
         14114 => x"38",
         14115 => x"81",
         14116 => x"81",
         14117 => x"8a",
         14118 => x"77",
         14119 => x"38",
         14120 => x"7a",
         14121 => x"38",
         14122 => x"84",
         14123 => x"8e",
         14124 => x"f7",
         14125 => x"02",
         14126 => x"05",
         14127 => x"77",
         14128 => x"d5",
         14129 => x"08",
         14130 => x"24",
         14131 => x"17",
         14132 => x"8c",
         14133 => x"77",
         14134 => x"16",
         14135 => x"24",
         14136 => x"84",
         14137 => x"19",
         14138 => x"8b",
         14139 => x"8b",
         14140 => x"54",
         14141 => x"17",
         14142 => x"51",
         14143 => x"3f",
         14144 => x"70",
         14145 => x"07",
         14146 => x"30",
         14147 => x"81",
         14148 => x"0c",
         14149 => x"d3",
         14150 => x"76",
         14151 => x"3f",
         14152 => x"e3",
         14153 => x"80",
         14154 => x"8d",
         14155 => x"80",
         14156 => x"55",
         14157 => x"81",
         14158 => x"ff",
         14159 => x"f4",
         14160 => x"08",
         14161 => x"8a",
         14162 => x"38",
         14163 => x"76",
         14164 => x"38",
         14165 => x"8c",
         14166 => x"77",
         14167 => x"16",
         14168 => x"24",
         14169 => x"84",
         14170 => x"19",
         14171 => x"7c",
         14172 => x"24",
         14173 => x"3d",
         14174 => x"55",
         14175 => x"05",
         14176 => x"51",
         14177 => x"3f",
         14178 => x"08",
         14179 => x"7a",
         14180 => x"ff",
         14181 => x"84",
         14182 => x"0d",
         14183 => x"ff",
         14184 => x"75",
         14185 => x"52",
         14186 => x"ff",
         14187 => x"74",
         14188 => x"30",
         14189 => x"9f",
         14190 => x"52",
         14191 => x"ff",
         14192 => x"52",
         14193 => x"eb",
         14194 => x"39",
         14195 => x"84",
         14196 => x"0d",
         14197 => x"0d",
         14198 => x"05",
         14199 => x"52",
         14200 => x"72",
         14201 => x"90",
         14202 => x"ff",
         14203 => x"71",
         14204 => x"0c",
         14205 => x"04",
         14206 => x"73",
         14207 => x"83",
         14208 => x"81",
         14209 => x"73",
         14210 => x"38",
         14211 => x"22",
         14212 => x"2e",
         14213 => x"12",
         14214 => x"ff",
         14215 => x"71",
         14216 => x"8d",
         14217 => x"83",
         14218 => x"70",
         14219 => x"e1",
         14220 => x"12",
         14221 => x"06",
         14222 => x"0c",
         14223 => x"0d",
         14224 => x"0d",
         14225 => x"22",
         14226 => x"96",
         14227 => x"51",
         14228 => x"80",
         14229 => x"38",
         14230 => x"84",
         14231 => x"84",
         14232 => x"71",
         14233 => x"09",
         14234 => x"38",
         14235 => x"26",
         14236 => x"10",
         14237 => x"05",
         14238 => x"bb",
         14239 => x"84",
         14240 => x"fb",
         14241 => x"51",
         14242 => x"ff",
         14243 => x"38",
         14244 => x"ff",
         14245 => x"c8",
         14246 => x"9f",
         14247 => x"d9",
         14248 => x"82",
         14249 => x"75",
         14250 => x"80",
         14251 => x"26",
         14252 => x"53",
         14253 => x"38",
         14254 => x"05",
         14255 => x"71",
         14256 => x"56",
         14257 => x"70",
         14258 => x"70",
         14259 => x"38",
         14260 => x"73",
         14261 => x"70",
         14262 => x"22",
         14263 => x"70",
         14264 => x"79",
         14265 => x"55",
         14266 => x"2e",
         14267 => x"51",
         14268 => x"84",
         14269 => x"0d",
         14270 => x"bc",
         14271 => x"39",
         14272 => x"ea",
         14273 => x"10",
         14274 => x"05",
         14275 => x"04",
         14276 => x"70",
         14277 => x"06",
         14278 => x"51",
         14279 => x"b0",
         14280 => x"ff",
         14281 => x"51",
         14282 => x"16",
         14283 => x"ff",
         14284 => x"e6",
         14285 => x"70",
         14286 => x"06",
         14287 => x"39",
         14288 => x"83",
         14289 => x"57",
         14290 => x"e0",
         14291 => x"ff",
         14292 => x"51",
         14293 => x"16",
         14294 => x"ff",
         14295 => x"ff",
         14296 => x"73",
         14297 => x"76",
         14298 => x"83",
         14299 => x"58",
         14300 => x"a6",
         14301 => x"31",
         14302 => x"70",
         14303 => x"fe",
         14304 => x"00",
         14305 => x"ff",
         14306 => x"ff",
         14307 => x"00",
         14308 => x"ff",
         14309 => x"19",
         14310 => x"19",
         14311 => x"19",
         14312 => x"19",
         14313 => x"19",
         14314 => x"19",
         14315 => x"19",
         14316 => x"19",
         14317 => x"19",
         14318 => x"19",
         14319 => x"19",
         14320 => x"19",
         14321 => x"19",
         14322 => x"18",
         14323 => x"18",
         14324 => x"18",
         14325 => x"18",
         14326 => x"18",
         14327 => x"18",
         14328 => x"18",
         14329 => x"1e",
         14330 => x"1f",
         14331 => x"1f",
         14332 => x"1f",
         14333 => x"1f",
         14334 => x"1f",
         14335 => x"1f",
         14336 => x"1f",
         14337 => x"1f",
         14338 => x"1f",
         14339 => x"1f",
         14340 => x"1f",
         14341 => x"1f",
         14342 => x"1f",
         14343 => x"1f",
         14344 => x"1f",
         14345 => x"1f",
         14346 => x"1f",
         14347 => x"1f",
         14348 => x"1f",
         14349 => x"1f",
         14350 => x"1f",
         14351 => x"1f",
         14352 => x"1f",
         14353 => x"1f",
         14354 => x"1f",
         14355 => x"1f",
         14356 => x"1f",
         14357 => x"1f",
         14358 => x"1f",
         14359 => x"1f",
         14360 => x"1f",
         14361 => x"1f",
         14362 => x"1f",
         14363 => x"1f",
         14364 => x"1f",
         14365 => x"1f",
         14366 => x"1f",
         14367 => x"1f",
         14368 => x"1f",
         14369 => x"1f",
         14370 => x"1f",
         14371 => x"1f",
         14372 => x"24",
         14373 => x"1f",
         14374 => x"1f",
         14375 => x"1f",
         14376 => x"1f",
         14377 => x"1f",
         14378 => x"1f",
         14379 => x"1f",
         14380 => x"1f",
         14381 => x"1f",
         14382 => x"1f",
         14383 => x"1f",
         14384 => x"1f",
         14385 => x"1f",
         14386 => x"1f",
         14387 => x"1f",
         14388 => x"1f",
         14389 => x"24",
         14390 => x"23",
         14391 => x"1f",
         14392 => x"22",
         14393 => x"24",
         14394 => x"23",
         14395 => x"22",
         14396 => x"21",
         14397 => x"1f",
         14398 => x"1f",
         14399 => x"1f",
         14400 => x"1f",
         14401 => x"1f",
         14402 => x"1f",
         14403 => x"1f",
         14404 => x"1f",
         14405 => x"1f",
         14406 => x"1f",
         14407 => x"1f",
         14408 => x"1f",
         14409 => x"1f",
         14410 => x"1f",
         14411 => x"1f",
         14412 => x"1f",
         14413 => x"1f",
         14414 => x"1f",
         14415 => x"1f",
         14416 => x"1f",
         14417 => x"1f",
         14418 => x"1f",
         14419 => x"1f",
         14420 => x"1f",
         14421 => x"1f",
         14422 => x"1f",
         14423 => x"1f",
         14424 => x"1f",
         14425 => x"1f",
         14426 => x"1f",
         14427 => x"1f",
         14428 => x"1f",
         14429 => x"1f",
         14430 => x"1f",
         14431 => x"1f",
         14432 => x"1f",
         14433 => x"1f",
         14434 => x"1f",
         14435 => x"1f",
         14436 => x"1f",
         14437 => x"1f",
         14438 => x"1f",
         14439 => x"1f",
         14440 => x"1f",
         14441 => x"1f",
         14442 => x"1f",
         14443 => x"1f",
         14444 => x"1f",
         14445 => x"1f",
         14446 => x"1f",
         14447 => x"1f",
         14448 => x"1f",
         14449 => x"21",
         14450 => x"21",
         14451 => x"1f",
         14452 => x"1f",
         14453 => x"1f",
         14454 => x"1f",
         14455 => x"1f",
         14456 => x"1f",
         14457 => x"1f",
         14458 => x"1f",
         14459 => x"21",
         14460 => x"21",
         14461 => x"1f",
         14462 => x"21",
         14463 => x"1f",
         14464 => x"21",
         14465 => x"21",
         14466 => x"21",
         14467 => x"32",
         14468 => x"32",
         14469 => x"32",
         14470 => x"32",
         14471 => x"32",
         14472 => x"32",
         14473 => x"3c",
         14474 => x"3a",
         14475 => x"39",
         14476 => x"36",
         14477 => x"3b",
         14478 => x"34",
         14479 => x"37",
         14480 => x"36",
         14481 => x"3a",
         14482 => x"36",
         14483 => x"37",
         14484 => x"39",
         14485 => x"34",
         14486 => x"39",
         14487 => x"38",
         14488 => x"37",
         14489 => x"34",
         14490 => x"34",
         14491 => x"37",
         14492 => x"36",
         14493 => x"36",
         14494 => x"36",
         14495 => x"47",
         14496 => x"47",
         14497 => x"47",
         14498 => x"47",
         14499 => x"47",
         14500 => x"47",
         14501 => x"47",
         14502 => x"48",
         14503 => x"48",
         14504 => x"48",
         14505 => x"48",
         14506 => x"48",
         14507 => x"48",
         14508 => x"48",
         14509 => x"48",
         14510 => x"48",
         14511 => x"48",
         14512 => x"48",
         14513 => x"48",
         14514 => x"48",
         14515 => x"48",
         14516 => x"48",
         14517 => x"48",
         14518 => x"48",
         14519 => x"48",
         14520 => x"48",
         14521 => x"48",
         14522 => x"48",
         14523 => x"48",
         14524 => x"48",
         14525 => x"48",
         14526 => x"48",
         14527 => x"48",
         14528 => x"48",
         14529 => x"48",
         14530 => x"48",
         14531 => x"48",
         14532 => x"49",
         14533 => x"49",
         14534 => x"49",
         14535 => x"49",
         14536 => x"48",
         14537 => x"48",
         14538 => x"48",
         14539 => x"48",
         14540 => x"48",
         14541 => x"48",
         14542 => x"48",
         14543 => x"49",
         14544 => x"48",
         14545 => x"48",
         14546 => x"48",
         14547 => x"48",
         14548 => x"48",
         14549 => x"48",
         14550 => x"48",
         14551 => x"48",
         14552 => x"54",
         14553 => x"56",
         14554 => x"56",
         14555 => x"55",
         14556 => x"55",
         14557 => x"55",
         14558 => x"54",
         14559 => x"56",
         14560 => x"53",
         14561 => x"56",
         14562 => x"58",
         14563 => x"53",
         14564 => x"53",
         14565 => x"53",
         14566 => x"53",
         14567 => x"53",
         14568 => x"53",
         14569 => x"56",
         14570 => x"58",
         14571 => x"57",
         14572 => x"53",
         14573 => x"53",
         14574 => x"53",
         14575 => x"53",
         14576 => x"53",
         14577 => x"53",
         14578 => x"53",
         14579 => x"53",
         14580 => x"53",
         14581 => x"53",
         14582 => x"53",
         14583 => x"53",
         14584 => x"53",
         14585 => x"53",
         14586 => x"53",
         14587 => x"53",
         14588 => x"53",
         14589 => x"53",
         14590 => x"53",
         14591 => x"55",
         14592 => x"53",
         14593 => x"53",
         14594 => x"53",
         14595 => x"55",
         14596 => x"54",
         14597 => x"54",
         14598 => x"53",
         14599 => x"53",
         14600 => x"53",
         14601 => x"53",
         14602 => x"54",
         14603 => x"53",
         14604 => x"54",
         14605 => x"5a",
         14606 => x"59",
         14607 => x"59",
         14608 => x"59",
         14609 => x"59",
         14610 => x"59",
         14611 => x"59",
         14612 => x"59",
         14613 => x"59",
         14614 => x"59",
         14615 => x"59",
         14616 => x"59",
         14617 => x"59",
         14618 => x"59",
         14619 => x"59",
         14620 => x"59",
         14621 => x"59",
         14622 => x"59",
         14623 => x"59",
         14624 => x"59",
         14625 => x"59",
         14626 => x"59",
         14627 => x"59",
         14628 => x"59",
         14629 => x"59",
         14630 => x"59",
         14631 => x"59",
         14632 => x"59",
         14633 => x"59",
         14634 => x"59",
         14635 => x"5a",
         14636 => x"5a",
         14637 => x"5a",
         14638 => x"5a",
         14639 => x"5a",
         14640 => x"5b",
         14641 => x"5b",
         14642 => x"5b",
         14643 => x"59",
         14644 => x"5b",
         14645 => x"5b",
         14646 => x"5b",
         14647 => x"5a",
         14648 => x"5a",
         14649 => x"5a",
         14650 => x"5a",
         14651 => x"5a",
         14652 => x"5a",
         14653 => x"59",
         14654 => x"5a",
         14655 => x"64",
         14656 => x"62",
         14657 => x"62",
         14658 => x"62",
         14659 => x"62",
         14660 => x"62",
         14661 => x"62",
         14662 => x"62",
         14663 => x"62",
         14664 => x"62",
         14665 => x"62",
         14666 => x"62",
         14667 => x"62",
         14668 => x"62",
         14669 => x"5f",
         14670 => x"62",
         14671 => x"62",
         14672 => x"62",
         14673 => x"62",
         14674 => x"62",
         14675 => x"62",
         14676 => x"64",
         14677 => x"62",
         14678 => x"62",
         14679 => x"64",
         14680 => x"62",
         14681 => x"64",
         14682 => x"5f",
         14683 => x"64",
         14684 => x"df",
         14685 => x"df",
         14686 => x"df",
         14687 => x"df",
         14688 => x"df",
         14689 => x"df",
         14690 => x"df",
         14691 => x"df",
         14692 => x"df",
         14693 => x"0e",
         14694 => x"0b",
         14695 => x"0b",
         14696 => x"0f",
         14697 => x"0b",
         14698 => x"0b",
         14699 => x"0b",
         14700 => x"0b",
         14701 => x"0b",
         14702 => x"0b",
         14703 => x"0b",
         14704 => x"0d",
         14705 => x"0b",
         14706 => x"0f",
         14707 => x"0f",
         14708 => x"0b",
         14709 => x"0b",
         14710 => x"0b",
         14711 => x"0b",
         14712 => x"0b",
         14713 => x"0b",
         14714 => x"0b",
         14715 => x"0b",
         14716 => x"0b",
         14717 => x"0b",
         14718 => x"0b",
         14719 => x"0b",
         14720 => x"0b",
         14721 => x"0b",
         14722 => x"0b",
         14723 => x"0b",
         14724 => x"0b",
         14725 => x"0b",
         14726 => x"0b",
         14727 => x"0b",
         14728 => x"0b",
         14729 => x"0b",
         14730 => x"0b",
         14731 => x"0b",
         14732 => x"0b",
         14733 => x"0b",
         14734 => x"0b",
         14735 => x"0b",
         14736 => x"0b",
         14737 => x"0b",
         14738 => x"0b",
         14739 => x"0b",
         14740 => x"0b",
         14741 => x"0b",
         14742 => x"0b",
         14743 => x"0b",
         14744 => x"0f",
         14745 => x"0b",
         14746 => x"0b",
         14747 => x"0b",
         14748 => x"0b",
         14749 => x"0e",
         14750 => x"0b",
         14751 => x"0b",
         14752 => x"0b",
         14753 => x"0b",
         14754 => x"0b",
         14755 => x"0b",
         14756 => x"0b",
         14757 => x"0b",
         14758 => x"0b",
         14759 => x"0b",
         14760 => x"0e",
         14761 => x"0e",
         14762 => x"0e",
         14763 => x"0e",
         14764 => x"0e",
         14765 => x"0b",
         14766 => x"0e",
         14767 => x"0b",
         14768 => x"0b",
         14769 => x"0e",
         14770 => x"0b",
         14771 => x"0b",
         14772 => x"0c",
         14773 => x"0e",
         14774 => x"0b",
         14775 => x"0b",
         14776 => x"0f",
         14777 => x"0b",
         14778 => x"0c",
         14779 => x"0b",
         14780 => x"0b",
         14781 => x"0e",
         14782 => x"6e",
         14783 => x"00",
         14784 => x"6f",
         14785 => x"00",
         14786 => x"6e",
         14787 => x"00",
         14788 => x"6f",
         14789 => x"00",
         14790 => x"78",
         14791 => x"00",
         14792 => x"6c",
         14793 => x"00",
         14794 => x"6f",
         14795 => x"00",
         14796 => x"69",
         14797 => x"00",
         14798 => x"75",
         14799 => x"00",
         14800 => x"62",
         14801 => x"68",
         14802 => x"77",
         14803 => x"64",
         14804 => x"65",
         14805 => x"64",
         14806 => x"65",
         14807 => x"6c",
         14808 => x"00",
         14809 => x"70",
         14810 => x"73",
         14811 => x"74",
         14812 => x"73",
         14813 => x"00",
         14814 => x"66",
         14815 => x"00",
         14816 => x"73",
         14817 => x"00",
         14818 => x"73",
         14819 => x"30",
         14820 => x"61",
         14821 => x"00",
         14822 => x"61",
         14823 => x"00",
         14824 => x"6c",
         14825 => x"00",
         14826 => x"00",
         14827 => x"6b",
         14828 => x"6e",
         14829 => x"72",
         14830 => x"00",
         14831 => x"72",
         14832 => x"74",
         14833 => x"20",
         14834 => x"6f",
         14835 => x"63",
         14836 => x"00",
         14837 => x"6f",
         14838 => x"6e",
         14839 => x"70",
         14840 => x"66",
         14841 => x"73",
         14842 => x"00",
         14843 => x"73",
         14844 => x"69",
         14845 => x"6e",
         14846 => x"65",
         14847 => x"79",
         14848 => x"00",
         14849 => x"6c",
         14850 => x"73",
         14851 => x"63",
         14852 => x"2e",
         14853 => x"6d",
         14854 => x"74",
         14855 => x"70",
         14856 => x"74",
         14857 => x"20",
         14858 => x"63",
         14859 => x"65",
         14860 => x"00",
         14861 => x"72",
         14862 => x"20",
         14863 => x"72",
         14864 => x"2e",
         14865 => x"20",
         14866 => x"70",
         14867 => x"62",
         14868 => x"66",
         14869 => x"73",
         14870 => x"65",
         14871 => x"6f",
         14872 => x"20",
         14873 => x"64",
         14874 => x"2e",
         14875 => x"73",
         14876 => x"6f",
         14877 => x"6e",
         14878 => x"65",
         14879 => x"00",
         14880 => x"69",
         14881 => x"6e",
         14882 => x"65",
         14883 => x"73",
         14884 => x"76",
         14885 => x"64",
         14886 => x"00",
         14887 => x"20",
         14888 => x"77",
         14889 => x"65",
         14890 => x"6f",
         14891 => x"74",
         14892 => x"00",
         14893 => x"6c",
         14894 => x"61",
         14895 => x"65",
         14896 => x"76",
         14897 => x"64",
         14898 => x"00",
         14899 => x"6c",
         14900 => x"6c",
         14901 => x"64",
         14902 => x"78",
         14903 => x"73",
         14904 => x"00",
         14905 => x"63",
         14906 => x"20",
         14907 => x"69",
         14908 => x"00",
         14909 => x"76",
         14910 => x"64",
         14911 => x"6c",
         14912 => x"6d",
         14913 => x"00",
         14914 => x"20",
         14915 => x"68",
         14916 => x"75",
         14917 => x"00",
         14918 => x"20",
         14919 => x"65",
         14920 => x"75",
         14921 => x"00",
         14922 => x"73",
         14923 => x"6f",
         14924 => x"65",
         14925 => x"2e",
         14926 => x"74",
         14927 => x"61",
         14928 => x"72",
         14929 => x"2e",
         14930 => x"73",
         14931 => x"72",
         14932 => x"00",
         14933 => x"63",
         14934 => x"73",
         14935 => x"00",
         14936 => x"6c",
         14937 => x"79",
         14938 => x"20",
         14939 => x"61",
         14940 => x"6c",
         14941 => x"79",
         14942 => x"2f",
         14943 => x"2e",
         14944 => x"00",
         14945 => x"61",
         14946 => x"00",
         14947 => x"38",
         14948 => x"00",
         14949 => x"20",
         14950 => x"32",
         14951 => x"00",
         14952 => x"00",
         14953 => x"00",
         14954 => x"00",
         14955 => x"34",
         14956 => x"00",
         14957 => x"20",
         14958 => x"20",
         14959 => x"00",
         14960 => x"53",
         14961 => x"20",
         14962 => x"28",
         14963 => x"2f",
         14964 => x"32",
         14965 => x"00",
         14966 => x"2e",
         14967 => x"00",
         14968 => x"50",
         14969 => x"72",
         14970 => x"25",
         14971 => x"29",
         14972 => x"20",
         14973 => x"2a",
         14974 => x"00",
         14975 => x"3a",
         14976 => x"20",
         14977 => x"73",
         14978 => x"64",
         14979 => x"73",
         14980 => x"20",
         14981 => x"20",
         14982 => x"20",
         14983 => x"20",
         14984 => x"6c",
         14985 => x"00",
         14986 => x"20",
         14987 => x"70",
         14988 => x"64",
         14989 => x"73",
         14990 => x"20",
         14991 => x"20",
         14992 => x"20",
         14993 => x"20",
         14994 => x"6c",
         14995 => x"00",
         14996 => x"55",
         14997 => x"74",
         14998 => x"75",
         14999 => x"48",
         15000 => x"6c",
         15001 => x"00",
         15002 => x"52",
         15003 => x"54",
         15004 => x"6e",
         15005 => x"72",
         15006 => x"00",
         15007 => x"52",
         15008 => x"52",
         15009 => x"6e",
         15010 => x"72",
         15011 => x"00",
         15012 => x"52",
         15013 => x"54",
         15014 => x"6e",
         15015 => x"72",
         15016 => x"00",
         15017 => x"52",
         15018 => x"52",
         15019 => x"6e",
         15020 => x"72",
         15021 => x"00",
         15022 => x"43",
         15023 => x"57",
         15024 => x"6e",
         15025 => x"72",
         15026 => x"00",
         15027 => x"43",
         15028 => x"52",
         15029 => x"6e",
         15030 => x"72",
         15031 => x"00",
         15032 => x"32",
         15033 => x"74",
         15034 => x"75",
         15035 => x"00",
         15036 => x"6d",
         15037 => x"69",
         15038 => x"72",
         15039 => x"74",
         15040 => x"74",
         15041 => x"67",
         15042 => x"20",
         15043 => x"65",
         15044 => x"2e",
         15045 => x"61",
         15046 => x"6e",
         15047 => x"69",
         15048 => x"2e",
         15049 => x"00",
         15050 => x"74",
         15051 => x"65",
         15052 => x"61",
         15053 => x"00",
         15054 => x"53",
         15055 => x"75",
         15056 => x"74",
         15057 => x"69",
         15058 => x"20",
         15059 => x"69",
         15060 => x"69",
         15061 => x"73",
         15062 => x"64",
         15063 => x"72",
         15064 => x"2c",
         15065 => x"65",
         15066 => x"20",
         15067 => x"74",
         15068 => x"6e",
         15069 => x"6c",
         15070 => x"00",
         15071 => x"00",
         15072 => x"3a",
         15073 => x"00",
         15074 => x"00",
         15075 => x"64",
         15076 => x"6d",
         15077 => x"64",
         15078 => x"00",
         15079 => x"55",
         15080 => x"6e",
         15081 => x"3a",
         15082 => x"5c",
         15083 => x"25",
         15084 => x"00",
         15085 => x"6c",
         15086 => x"65",
         15087 => x"74",
         15088 => x"2e",
         15089 => x"00",
         15090 => x"73",
         15091 => x"74",
         15092 => x"20",
         15093 => x"6c",
         15094 => x"74",
         15095 => x"2e",
         15096 => x"00",
         15097 => x"6c",
         15098 => x"67",
         15099 => x"64",
         15100 => x"20",
         15101 => x"6c",
         15102 => x"2e",
         15103 => x"00",
         15104 => x"6c",
         15105 => x"65",
         15106 => x"6e",
         15107 => x"63",
         15108 => x"20",
         15109 => x"29",
         15110 => x"00",
         15111 => x"65",
         15112 => x"69",
         15113 => x"63",
         15114 => x"20",
         15115 => x"30",
         15116 => x"20",
         15117 => x"0a",
         15118 => x"38",
         15119 => x"25",
         15120 => x"58",
         15121 => x"00",
         15122 => x"38",
         15123 => x"25",
         15124 => x"2d",
         15125 => x"6d",
         15126 => x"69",
         15127 => x"2e",
         15128 => x"00",
         15129 => x"38",
         15130 => x"25",
         15131 => x"29",
         15132 => x"30",
         15133 => x"28",
         15134 => x"78",
         15135 => x"00",
         15136 => x"70",
         15137 => x"67",
         15138 => x"00",
         15139 => x"38",
         15140 => x"25",
         15141 => x"2d",
         15142 => x"65",
         15143 => x"6e",
         15144 => x"2e",
         15145 => x"00",
         15146 => x"6d",
         15147 => x"65",
         15148 => x"79",
         15149 => x"6f",
         15150 => x"65",
         15151 => x"00",
         15152 => x"3a",
         15153 => x"5c",
         15154 => x"00",
         15155 => x"6d",
         15156 => x"20",
         15157 => x"61",
         15158 => x"65",
         15159 => x"63",
         15160 => x"6f",
         15161 => x"72",
         15162 => x"73",
         15163 => x"6f",
         15164 => x"6e",
         15165 => x"00",
         15166 => x"3f",
         15167 => x"2f",
         15168 => x"25",
         15169 => x"64",
         15170 => x"3a",
         15171 => x"25",
         15172 => x"0a",
         15173 => x"43",
         15174 => x"6e",
         15175 => x"75",
         15176 => x"69",
         15177 => x"00",
         15178 => x"44",
         15179 => x"63",
         15180 => x"69",
         15181 => x"65",
         15182 => x"74",
         15183 => x"00",
         15184 => x"64",
         15185 => x"73",
         15186 => x"00",
         15187 => x"20",
         15188 => x"55",
         15189 => x"73",
         15190 => x"56",
         15191 => x"6f",
         15192 => x"64",
         15193 => x"73",
         15194 => x"20",
         15195 => x"58",
         15196 => x"00",
         15197 => x"20",
         15198 => x"55",
         15199 => x"6d",
         15200 => x"20",
         15201 => x"72",
         15202 => x"64",
         15203 => x"73",
         15204 => x"20",
         15205 => x"58",
         15206 => x"00",
         15207 => x"20",
         15208 => x"61",
         15209 => x"53",
         15210 => x"74",
         15211 => x"64",
         15212 => x"73",
         15213 => x"20",
         15214 => x"20",
         15215 => x"58",
         15216 => x"00",
         15217 => x"73",
         15218 => x"00",
         15219 => x"20",
         15220 => x"55",
         15221 => x"20",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"20",
         15226 => x"20",
         15227 => x"58",
         15228 => x"00",
         15229 => x"20",
         15230 => x"73",
         15231 => x"20",
         15232 => x"63",
         15233 => x"72",
         15234 => x"20",
         15235 => x"20",
         15236 => x"20",
         15237 => x"25",
         15238 => x"4d",
         15239 => x"00",
         15240 => x"20",
         15241 => x"73",
         15242 => x"6e",
         15243 => x"44",
         15244 => x"20",
         15245 => x"63",
         15246 => x"72",
         15247 => x"20",
         15248 => x"25",
         15249 => x"4d",
         15250 => x"00",
         15251 => x"20",
         15252 => x"52",
         15253 => x"43",
         15254 => x"6b",
         15255 => x"65",
         15256 => x"20",
         15257 => x"20",
         15258 => x"20",
         15259 => x"25",
         15260 => x"4d",
         15261 => x"00",
         15262 => x"20",
         15263 => x"49",
         15264 => x"20",
         15265 => x"32",
         15266 => x"20",
         15267 => x"43",
         15268 => x"00",
         15269 => x"20",
         15270 => x"20",
         15271 => x"00",
         15272 => x"20",
         15273 => x"53",
         15274 => x"4e",
         15275 => x"55",
         15276 => x"00",
         15277 => x"20",
         15278 => x"54",
         15279 => x"54",
         15280 => x"28",
         15281 => x"6e",
         15282 => x"73",
         15283 => x"32",
         15284 => x"0a",
         15285 => x"20",
         15286 => x"4d",
         15287 => x"20",
         15288 => x"28",
         15289 => x"65",
         15290 => x"20",
         15291 => x"32",
         15292 => x"0a",
         15293 => x"20",
         15294 => x"20",
         15295 => x"44",
         15296 => x"28",
         15297 => x"69",
         15298 => x"20",
         15299 => x"32",
         15300 => x"0a",
         15301 => x"20",
         15302 => x"4d",
         15303 => x"20",
         15304 => x"28",
         15305 => x"58",
         15306 => x"38",
         15307 => x"0a",
         15308 => x"20",
         15309 => x"41",
         15310 => x"20",
         15311 => x"28",
         15312 => x"58",
         15313 => x"38",
         15314 => x"0a",
         15315 => x"20",
         15316 => x"53",
         15317 => x"52",
         15318 => x"28",
         15319 => x"58",
         15320 => x"38",
         15321 => x"0a",
         15322 => x"20",
         15323 => x"52",
         15324 => x"20",
         15325 => x"28",
         15326 => x"58",
         15327 => x"38",
         15328 => x"0a",
         15329 => x"20",
         15330 => x"20",
         15331 => x"41",
         15332 => x"28",
         15333 => x"58",
         15334 => x"38",
         15335 => x"0a",
         15336 => x"66",
         15337 => x"20",
         15338 => x"20",
         15339 => x"66",
         15340 => x"00",
         15341 => x"6b",
         15342 => x"6e",
         15343 => x"4f",
         15344 => x"00",
         15345 => x"61",
         15346 => x"00",
         15347 => x"64",
         15348 => x"00",
         15349 => x"65",
         15350 => x"00",
         15351 => x"4f",
         15352 => x"f1",
         15353 => x"00",
         15354 => x"00",
         15355 => x"f1",
         15356 => x"00",
         15357 => x"00",
         15358 => x"f1",
         15359 => x"00",
         15360 => x"00",
         15361 => x"f1",
         15362 => x"00",
         15363 => x"00",
         15364 => x"f1",
         15365 => x"00",
         15366 => x"00",
         15367 => x"f1",
         15368 => x"00",
         15369 => x"00",
         15370 => x"f1",
         15371 => x"00",
         15372 => x"00",
         15373 => x"f1",
         15374 => x"00",
         15375 => x"00",
         15376 => x"f1",
         15377 => x"00",
         15378 => x"00",
         15379 => x"f1",
         15380 => x"00",
         15381 => x"00",
         15382 => x"f1",
         15383 => x"00",
         15384 => x"00",
         15385 => x"f1",
         15386 => x"00",
         15387 => x"00",
         15388 => x"f1",
         15389 => x"00",
         15390 => x"00",
         15391 => x"f1",
         15392 => x"00",
         15393 => x"00",
         15394 => x"f1",
         15395 => x"00",
         15396 => x"00",
         15397 => x"f1",
         15398 => x"00",
         15399 => x"00",
         15400 => x"f0",
         15401 => x"00",
         15402 => x"00",
         15403 => x"f0",
         15404 => x"00",
         15405 => x"00",
         15406 => x"f0",
         15407 => x"00",
         15408 => x"00",
         15409 => x"f0",
         15410 => x"00",
         15411 => x"00",
         15412 => x"f0",
         15413 => x"00",
         15414 => x"00",
         15415 => x"f0",
         15416 => x"00",
         15417 => x"00",
         15418 => x"44",
         15419 => x"43",
         15420 => x"42",
         15421 => x"41",
         15422 => x"36",
         15423 => x"35",
         15424 => x"34",
         15425 => x"46",
         15426 => x"33",
         15427 => x"32",
         15428 => x"31",
         15429 => x"00",
         15430 => x"00",
         15431 => x"00",
         15432 => x"00",
         15433 => x"00",
         15434 => x"00",
         15435 => x"00",
         15436 => x"00",
         15437 => x"00",
         15438 => x"00",
         15439 => x"00",
         15440 => x"73",
         15441 => x"79",
         15442 => x"61",
         15443 => x"30",
         15444 => x"0a",
         15445 => x"6e",
         15446 => x"20",
         15447 => x"6e",
         15448 => x"65",
         15449 => x"20",
         15450 => x"74",
         15451 => x"20",
         15452 => x"65",
         15453 => x"69",
         15454 => x"6c",
         15455 => x"2e",
         15456 => x"73",
         15457 => x"79",
         15458 => x"73",
         15459 => x"00",
         15460 => x"00",
         15461 => x"73",
         15462 => x"79",
         15463 => x"66",
         15464 => x"40",
         15465 => x"6c",
         15466 => x"00",
         15467 => x"36",
         15468 => x"20",
         15469 => x"00",
         15470 => x"69",
         15471 => x"20",
         15472 => x"72",
         15473 => x"74",
         15474 => x"65",
         15475 => x"73",
         15476 => x"79",
         15477 => x"6c",
         15478 => x"6f",
         15479 => x"46",
         15480 => x"00",
         15481 => x"73",
         15482 => x"00",
         15483 => x"31",
         15484 => x"00",
         15485 => x"41",
         15486 => x"42",
         15487 => x"43",
         15488 => x"44",
         15489 => x"31",
         15490 => x"00",
         15491 => x"31",
         15492 => x"00",
         15493 => x"31",
         15494 => x"00",
         15495 => x"31",
         15496 => x"00",
         15497 => x"31",
         15498 => x"00",
         15499 => x"31",
         15500 => x"00",
         15501 => x"31",
         15502 => x"00",
         15503 => x"31",
         15504 => x"00",
         15505 => x"31",
         15506 => x"00",
         15507 => x"32",
         15508 => x"00",
         15509 => x"32",
         15510 => x"00",
         15511 => x"33",
         15512 => x"00",
         15513 => x"46",
         15514 => x"35",
         15515 => x"00",
         15516 => x"36",
         15517 => x"00",
         15518 => x"25",
         15519 => x"64",
         15520 => x"2c",
         15521 => x"25",
         15522 => x"64",
         15523 => x"32",
         15524 => x"00",
         15525 => x"25",
         15526 => x"64",
         15527 => x"3a",
         15528 => x"25",
         15529 => x"64",
         15530 => x"3a",
         15531 => x"2c",
         15532 => x"25",
         15533 => x"00",
         15534 => x"32",
         15535 => x"00",
         15536 => x"5b",
         15537 => x"25",
         15538 => x"00",
         15539 => x"70",
         15540 => x"20",
         15541 => x"73",
         15542 => x"00",
         15543 => x"3a",
         15544 => x"78",
         15545 => x"32",
         15546 => x"00",
         15547 => x"3a",
         15548 => x"78",
         15549 => x"32",
         15550 => x"00",
         15551 => x"3a",
         15552 => x"78",
         15553 => x"00",
         15554 => x"20",
         15555 => x"74",
         15556 => x"66",
         15557 => x"64",
         15558 => x"00",
         15559 => x"00",
         15560 => x"3a",
         15561 => x"7c",
         15562 => x"00",
         15563 => x"3b",
         15564 => x"00",
         15565 => x"54",
         15566 => x"54",
         15567 => x"00",
         15568 => x"90",
         15569 => x"4f",
         15570 => x"30",
         15571 => x"20",
         15572 => x"45",
         15573 => x"20",
         15574 => x"20",
         15575 => x"20",
         15576 => x"20",
         15577 => x"45",
         15578 => x"20",
         15579 => x"33",
         15580 => x"20",
         15581 => x"f3",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"05",
         15586 => x"10",
         15587 => x"18",
         15588 => x"00",
         15589 => x"45",
         15590 => x"8f",
         15591 => x"45",
         15592 => x"8e",
         15593 => x"92",
         15594 => x"55",
         15595 => x"9a",
         15596 => x"9e",
         15597 => x"4f",
         15598 => x"a6",
         15599 => x"aa",
         15600 => x"ae",
         15601 => x"b2",
         15602 => x"b6",
         15603 => x"ba",
         15604 => x"be",
         15605 => x"c2",
         15606 => x"c6",
         15607 => x"ca",
         15608 => x"ce",
         15609 => x"d2",
         15610 => x"d6",
         15611 => x"da",
         15612 => x"de",
         15613 => x"e2",
         15614 => x"e6",
         15615 => x"ea",
         15616 => x"ee",
         15617 => x"f2",
         15618 => x"f6",
         15619 => x"fa",
         15620 => x"fe",
         15621 => x"2c",
         15622 => x"5d",
         15623 => x"2a",
         15624 => x"3f",
         15625 => x"00",
         15626 => x"00",
         15627 => x"00",
         15628 => x"02",
         15629 => x"00",
         15630 => x"00",
         15631 => x"00",
         15632 => x"00",
         15633 => x"00",
         15634 => x"00",
         15635 => x"00",
         15636 => x"00",
         15637 => x"00",
         15638 => x"00",
         15639 => x"00",
         15640 => x"00",
         15641 => x"00",
         15642 => x"00",
         15643 => x"00",
         15644 => x"00",
         15645 => x"00",
         15646 => x"00",
         15647 => x"00",
         15648 => x"00",
         15649 => x"01",
         15650 => x"00",
         15651 => x"00",
         15652 => x"00",
         15653 => x"00",
         15654 => x"23",
         15655 => x"00",
         15656 => x"00",
         15657 => x"00",
         15658 => x"25",
         15659 => x"25",
         15660 => x"25",
         15661 => x"25",
         15662 => x"25",
         15663 => x"25",
         15664 => x"25",
         15665 => x"25",
         15666 => x"25",
         15667 => x"25",
         15668 => x"25",
         15669 => x"25",
         15670 => x"25",
         15671 => x"25",
         15672 => x"25",
         15673 => x"25",
         15674 => x"25",
         15675 => x"25",
         15676 => x"25",
         15677 => x"25",
         15678 => x"25",
         15679 => x"25",
         15680 => x"25",
         15681 => x"25",
         15682 => x"00",
         15683 => x"03",
         15684 => x"03",
         15685 => x"03",
         15686 => x"03",
         15687 => x"03",
         15688 => x"03",
         15689 => x"22",
         15690 => x"00",
         15691 => x"22",
         15692 => x"23",
         15693 => x"22",
         15694 => x"22",
         15695 => x"22",
         15696 => x"00",
         15697 => x"00",
         15698 => x"03",
         15699 => x"03",
         15700 => x"03",
         15701 => x"00",
         15702 => x"01",
         15703 => x"01",
         15704 => x"01",
         15705 => x"01",
         15706 => x"01",
         15707 => x"01",
         15708 => x"02",
         15709 => x"01",
         15710 => x"01",
         15711 => x"01",
         15712 => x"01",
         15713 => x"01",
         15714 => x"01",
         15715 => x"01",
         15716 => x"01",
         15717 => x"01",
         15718 => x"01",
         15719 => x"01",
         15720 => x"01",
         15721 => x"02",
         15722 => x"01",
         15723 => x"02",
         15724 => x"01",
         15725 => x"01",
         15726 => x"01",
         15727 => x"01",
         15728 => x"01",
         15729 => x"01",
         15730 => x"01",
         15731 => x"01",
         15732 => x"01",
         15733 => x"01",
         15734 => x"01",
         15735 => x"01",
         15736 => x"01",
         15737 => x"01",
         15738 => x"01",
         15739 => x"01",
         15740 => x"01",
         15741 => x"01",
         15742 => x"01",
         15743 => x"01",
         15744 => x"01",
         15745 => x"01",
         15746 => x"01",
         15747 => x"01",
         15748 => x"00",
         15749 => x"01",
         15750 => x"01",
         15751 => x"01",
         15752 => x"01",
         15753 => x"01",
         15754 => x"01",
         15755 => x"00",
         15756 => x"02",
         15757 => x"02",
         15758 => x"02",
         15759 => x"02",
         15760 => x"02",
         15761 => x"02",
         15762 => x"01",
         15763 => x"02",
         15764 => x"01",
         15765 => x"01",
         15766 => x"01",
         15767 => x"02",
         15768 => x"02",
         15769 => x"02",
         15770 => x"01",
         15771 => x"02",
         15772 => x"02",
         15773 => x"01",
         15774 => x"2c",
         15775 => x"02",
         15776 => x"01",
         15777 => x"02",
         15778 => x"02",
         15779 => x"01",
         15780 => x"02",
         15781 => x"02",
         15782 => x"02",
         15783 => x"2c",
         15784 => x"02",
         15785 => x"02",
         15786 => x"01",
         15787 => x"02",
         15788 => x"02",
         15789 => x"02",
         15790 => x"01",
         15791 => x"02",
         15792 => x"02",
         15793 => x"02",
         15794 => x"03",
         15795 => x"03",
         15796 => x"03",
         15797 => x"00",
         15798 => x"03",
         15799 => x"03",
         15800 => x"03",
         15801 => x"00",
         15802 => x"03",
         15803 => x"03",
         15804 => x"00",
         15805 => x"03",
         15806 => x"03",
         15807 => x"03",
         15808 => x"03",
         15809 => x"03",
         15810 => x"03",
         15811 => x"03",
         15812 => x"03",
         15813 => x"04",
         15814 => x"04",
         15815 => x"04",
         15816 => x"04",
         15817 => x"04",
         15818 => x"04",
         15819 => x"04",
         15820 => x"01",
         15821 => x"04",
         15822 => x"00",
         15823 => x"00",
         15824 => x"1e",
         15825 => x"1e",
         15826 => x"1f",
         15827 => x"1f",
         15828 => x"1f",
         15829 => x"1f",
         15830 => x"1f",
         15831 => x"1f",
         15832 => x"1f",
         15833 => x"1f",
         15834 => x"1f",
         15835 => x"1f",
         15836 => x"06",
         15837 => x"00",
         15838 => x"1f",
         15839 => x"1f",
         15840 => x"1f",
         15841 => x"1f",
         15842 => x"1f",
         15843 => x"1f",
         15844 => x"1f",
         15845 => x"06",
         15846 => x"06",
         15847 => x"06",
         15848 => x"00",
         15849 => x"1f",
         15850 => x"1f",
         15851 => x"00",
         15852 => x"1f",
         15853 => x"1f",
         15854 => x"1f",
         15855 => x"1f",
         15856 => x"00",
         15857 => x"21",
         15858 => x"21",
         15859 => x"02",
         15860 => x"00",
         15861 => x"24",
         15862 => x"2c",
         15863 => x"2c",
         15864 => x"2c",
         15865 => x"2c",
         15866 => x"2c",
         15867 => x"2d",
         15868 => x"ff",
         15869 => x"00",
         15870 => x"00",
         15871 => x"e6",
         15872 => x"01",
         15873 => x"00",
         15874 => x"00",
         15875 => x"e7",
         15876 => x"01",
         15877 => x"00",
         15878 => x"00",
         15879 => x"e7",
         15880 => x"03",
         15881 => x"00",
         15882 => x"00",
         15883 => x"e7",
         15884 => x"03",
         15885 => x"00",
         15886 => x"00",
         15887 => x"e7",
         15888 => x"03",
         15889 => x"00",
         15890 => x"00",
         15891 => x"e7",
         15892 => x"04",
         15893 => x"00",
         15894 => x"00",
         15895 => x"e7",
         15896 => x"04",
         15897 => x"00",
         15898 => x"00",
         15899 => x"e7",
         15900 => x"04",
         15901 => x"00",
         15902 => x"00",
         15903 => x"e7",
         15904 => x"04",
         15905 => x"00",
         15906 => x"00",
         15907 => x"e7",
         15908 => x"04",
         15909 => x"00",
         15910 => x"00",
         15911 => x"e7",
         15912 => x"04",
         15913 => x"00",
         15914 => x"00",
         15915 => x"e7",
         15916 => x"04",
         15917 => x"00",
         15918 => x"00",
         15919 => x"e7",
         15920 => x"05",
         15921 => x"00",
         15922 => x"00",
         15923 => x"e7",
         15924 => x"05",
         15925 => x"00",
         15926 => x"00",
         15927 => x"e7",
         15928 => x"05",
         15929 => x"00",
         15930 => x"00",
         15931 => x"e7",
         15932 => x"05",
         15933 => x"00",
         15934 => x"00",
         15935 => x"e7",
         15936 => x"07",
         15937 => x"00",
         15938 => x"00",
         15939 => x"e7",
         15940 => x"07",
         15941 => x"00",
         15942 => x"00",
         15943 => x"e7",
         15944 => x"08",
         15945 => x"00",
         15946 => x"00",
         15947 => x"e7",
         15948 => x"08",
         15949 => x"00",
         15950 => x"00",
         15951 => x"e7",
         15952 => x"08",
         15953 => x"00",
         15954 => x"00",
         15955 => x"e7",
         15956 => x"08",
         15957 => x"00",
         15958 => x"00",
         15959 => x"e7",
         15960 => x"08",
         15961 => x"00",
         15962 => x"00",
         15963 => x"e7",
         15964 => x"08",
         15965 => x"00",
         15966 => x"00",
         15967 => x"e7",
         15968 => x"09",
         15969 => x"00",
         15970 => x"00",
         15971 => x"e7",
         15972 => x"09",
         15973 => x"00",
         15974 => x"00",
         15975 => x"e7",
         15976 => x"09",
         15977 => x"00",
         15978 => x"00",
         15979 => x"e7",
         15980 => x"09",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"7f",
         15986 => x"00",
         15987 => x"7f",
         15988 => x"00",
         15989 => x"7f",
         15990 => x"00",
         15991 => x"00",
         15992 => x"00",
         15993 => x"ff",
         15994 => x"00",
         15995 => x"00",
         15996 => x"78",
         15997 => x"00",
         15998 => x"e1",
         15999 => x"e1",
         16000 => x"e1",
         16001 => x"00",
         16002 => x"01",
         16003 => x"01",
         16004 => x"10",
         16005 => x"00",
         16006 => x"00",
         16007 => x"00",
         16008 => x"00",
         16009 => x"00",
         16010 => x"00",
         16011 => x"00",
         16012 => x"00",
         16013 => x"00",
         16014 => x"00",
         16015 => x"00",
         16016 => x"00",
         16017 => x"00",
         16018 => x"00",
         16019 => x"00",
         16020 => x"00",
         16021 => x"00",
         16022 => x"00",
         16023 => x"00",
         16024 => x"00",
         16025 => x"00",
         16026 => x"00",
         16027 => x"00",
         16028 => x"00",
         16029 => x"00",
         16030 => x"f1",
         16031 => x"00",
         16032 => x"f1",
         16033 => x"00",
         16034 => x"f1",
         16035 => x"00",
         16036 => x"fd",
         16037 => x"5f",
         16038 => x"3a",
         16039 => x"40",
         16040 => x"f0",
         16041 => x"73",
         16042 => x"77",
         16043 => x"6b",
         16044 => x"6f",
         16045 => x"63",
         16046 => x"67",
         16047 => x"33",
         16048 => x"37",
         16049 => x"2d",
         16050 => x"2c",
         16051 => x"f3",
         16052 => x"3f",
         16053 => x"f0",
         16054 => x"f0",
         16055 => x"82",
         16056 => x"f0",
         16057 => x"58",
         16058 => x"3b",
         16059 => x"40",
         16060 => x"f0",
         16061 => x"53",
         16062 => x"57",
         16063 => x"4b",
         16064 => x"4f",
         16065 => x"43",
         16066 => x"47",
         16067 => x"33",
         16068 => x"37",
         16069 => x"2d",
         16070 => x"2c",
         16071 => x"f3",
         16072 => x"3f",
         16073 => x"f0",
         16074 => x"f0",
         16075 => x"82",
         16076 => x"f0",
         16077 => x"58",
         16078 => x"2a",
         16079 => x"60",
         16080 => x"f0",
         16081 => x"53",
         16082 => x"57",
         16083 => x"4b",
         16084 => x"4f",
         16085 => x"43",
         16086 => x"47",
         16087 => x"23",
         16088 => x"27",
         16089 => x"3d",
         16090 => x"3c",
         16091 => x"e0",
         16092 => x"3f",
         16093 => x"f0",
         16094 => x"f0",
         16095 => x"87",
         16096 => x"f0",
         16097 => x"1e",
         16098 => x"f0",
         16099 => x"00",
         16100 => x"f0",
         16101 => x"13",
         16102 => x"17",
         16103 => x"0b",
         16104 => x"0f",
         16105 => x"03",
         16106 => x"07",
         16107 => x"f0",
         16108 => x"f0",
         16109 => x"f0",
         16110 => x"f0",
         16111 => x"f0",
         16112 => x"f0",
         16113 => x"f0",
         16114 => x"f0",
         16115 => x"82",
         16116 => x"f0",
         16117 => x"cf",
         16118 => x"4d",
         16119 => x"d7",
         16120 => x"f0",
         16121 => x"41",
         16122 => x"78",
         16123 => x"6c",
         16124 => x"d5",
         16125 => x"d9",
         16126 => x"4c",
         16127 => x"7e",
         16128 => x"5f",
         16129 => x"d1",
         16130 => x"d0",
         16131 => x"c2",
         16132 => x"bb",
         16133 => x"f0",
         16134 => x"f0",
         16135 => x"82",
         16136 => x"f0",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"00",
         16165 => x"f1",
         16166 => x"00",
         16167 => x"f1",
         16168 => x"00",
         16169 => x"f1",
         16170 => x"00",
         16171 => x"f1",
         16172 => x"00",
         16173 => x"f2",
         16174 => x"00",
         16175 => x"f2",
         16176 => x"00",
         16177 => x"f2",
         16178 => x"00",
         16179 => x"f2",
         16180 => x"00",
         16181 => x"f2",
         16182 => x"00",
         16183 => x"f2",
         16184 => x"00",
         16185 => x"f2",
         16186 => x"00",
         16187 => x"f2",
         16188 => x"00",
         16189 => x"f2",
         16190 => x"00",
         16191 => x"f2",
         16192 => x"00",
         16193 => x"f2",
         16194 => x"00",
         16195 => x"f2",
         16196 => x"00",
         16197 => x"f2",
         16198 => x"00",
         16199 => x"f2",
         16200 => x"00",
         16201 => x"f2",
         16202 => x"00",
         16203 => x"f2",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"32",
         18206 => x"01",
         18207 => x"00",
         18208 => x"f2",
         18209 => x"f6",
         18210 => x"fa",
         18211 => x"fe",
         18212 => x"c2",
         18213 => x"c6",
         18214 => x"e5",
         18215 => x"ef",
         18216 => x"62",
         18217 => x"66",
         18218 => x"6b",
         18219 => x"2e",
         18220 => x"22",
         18221 => x"26",
         18222 => x"4f",
         18223 => x"57",
         18224 => x"02",
         18225 => x"06",
         18226 => x"0a",
         18227 => x"0e",
         18228 => x"12",
         18229 => x"16",
         18230 => x"1a",
         18231 => x"be",
         18232 => x"82",
         18233 => x"86",
         18234 => x"8a",
         18235 => x"8e",
         18236 => x"92",
         18237 => x"96",
         18238 => x"9a",
         18239 => x"a5",
         18240 => x"00",
         18241 => x"00",
         18242 => x"00",
         18243 => x"00",
         18244 => x"00",
         18245 => x"00",
         18246 => x"00",
         18247 => x"00",
         18248 => x"00",
         18249 => x"00",
         18250 => x"00",
         18251 => x"00",
         18252 => x"00",
         18253 => x"00",
         18254 => x"00",
         18255 => x"00",
         18256 => x"00",
         18257 => x"00",
         18258 => x"00",
         18259 => x"00",
         18260 => x"00",
         18261 => x"00",
         18262 => x"00",
         18263 => x"00",
         18264 => x"00",
         18265 => x"00",
         18266 => x"00",
         18267 => x"00",
         18268 => x"00",
         18269 => x"00",
         18270 => x"00",
         18271 => x"01",
         18272 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"b5",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"91",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"92",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"84",
           386 => x"80",
           387 => x"84",
           388 => x"80",
           389 => x"04",
           390 => x"0c",
           391 => x"84",
           392 => x"80",
           393 => x"04",
           394 => x"0c",
           395 => x"84",
           396 => x"80",
           397 => x"04",
           398 => x"0c",
           399 => x"84",
           400 => x"80",
           401 => x"04",
           402 => x"0c",
           403 => x"84",
           404 => x"80",
           405 => x"04",
           406 => x"0c",
           407 => x"84",
           408 => x"80",
           409 => x"04",
           410 => x"0c",
           411 => x"84",
           412 => x"80",
           413 => x"04",
           414 => x"0c",
           415 => x"84",
           416 => x"80",
           417 => x"04",
           418 => x"0c",
           419 => x"84",
           420 => x"80",
           421 => x"04",
           422 => x"0c",
           423 => x"84",
           424 => x"80",
           425 => x"04",
           426 => x"0c",
           427 => x"84",
           428 => x"80",
           429 => x"04",
           430 => x"0c",
           431 => x"84",
           432 => x"80",
           433 => x"04",
           434 => x"0c",
           435 => x"2d",
           436 => x"08",
           437 => x"90",
           438 => x"90",
           439 => x"e1",
           440 => x"90",
           441 => x"80",
           442 => x"bb",
           443 => x"d2",
           444 => x"bb",
           445 => x"c0",
           446 => x"84",
           447 => x"80",
           448 => x"84",
           449 => x"80",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"90",
           455 => x"90",
           456 => x"89",
           457 => x"90",
           458 => x"80",
           459 => x"bb",
           460 => x"d4",
           461 => x"bb",
           462 => x"c0",
           463 => x"84",
           464 => x"82",
           465 => x"84",
           466 => x"80",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"90",
           472 => x"90",
           473 => x"fc",
           474 => x"90",
           475 => x"80",
           476 => x"bb",
           477 => x"de",
           478 => x"bb",
           479 => x"c0",
           480 => x"84",
           481 => x"82",
           482 => x"84",
           483 => x"80",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"90",
           489 => x"90",
           490 => x"b7",
           491 => x"90",
           492 => x"80",
           493 => x"bb",
           494 => x"85",
           495 => x"bb",
           496 => x"c0",
           497 => x"84",
           498 => x"82",
           499 => x"84",
           500 => x"80",
           501 => x"04",
           502 => x"0c",
           503 => x"2d",
           504 => x"08",
           505 => x"90",
           506 => x"90",
           507 => x"94",
           508 => x"90",
           509 => x"80",
           510 => x"bb",
           511 => x"95",
           512 => x"bb",
           513 => x"c0",
           514 => x"84",
           515 => x"83",
           516 => x"84",
           517 => x"80",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"90",
           523 => x"90",
           524 => x"f0",
           525 => x"90",
           526 => x"80",
           527 => x"bb",
           528 => x"e7",
           529 => x"bb",
           530 => x"c0",
           531 => x"84",
           532 => x"82",
           533 => x"84",
           534 => x"80",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"90",
           540 => x"90",
           541 => x"86",
           542 => x"90",
           543 => x"80",
           544 => x"bb",
           545 => x"a1",
           546 => x"bb",
           547 => x"c0",
           548 => x"84",
           549 => x"82",
           550 => x"84",
           551 => x"80",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"90",
           557 => x"90",
           558 => x"a2",
           559 => x"90",
           560 => x"80",
           561 => x"bb",
           562 => x"b8",
           563 => x"bb",
           564 => x"c0",
           565 => x"84",
           566 => x"81",
           567 => x"84",
           568 => x"80",
           569 => x"04",
           570 => x"0c",
           571 => x"2d",
           572 => x"08",
           573 => x"90",
           574 => x"90",
           575 => x"a9",
           576 => x"90",
           577 => x"80",
           578 => x"bb",
           579 => x"d0",
           580 => x"bb",
           581 => x"c0",
           582 => x"84",
           583 => x"80",
           584 => x"84",
           585 => x"80",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"90",
           591 => x"90",
           592 => x"2d",
           593 => x"08",
           594 => x"90",
           595 => x"90",
           596 => x"c9",
           597 => x"90",
           598 => x"80",
           599 => x"bb",
           600 => x"de",
           601 => x"bb",
           602 => x"c0",
           603 => x"84",
           604 => x"81",
           605 => x"84",
           606 => x"80",
           607 => x"04",
           608 => x"0c",
           609 => x"2d",
           610 => x"08",
           611 => x"90",
           612 => x"10",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"51",
           621 => x"73",
           622 => x"73",
           623 => x"81",
           624 => x"10",
           625 => x"07",
           626 => x"0c",
           627 => x"72",
           628 => x"81",
           629 => x"09",
           630 => x"71",
           631 => x"0a",
           632 => x"72",
           633 => x"51",
           634 => x"84",
           635 => x"84",
           636 => x"8e",
           637 => x"70",
           638 => x"0c",
           639 => x"93",
           640 => x"81",
           641 => x"ca",
           642 => x"3d",
           643 => x"70",
           644 => x"52",
           645 => x"74",
           646 => x"e8",
           647 => x"c5",
           648 => x"0d",
           649 => x"0d",
           650 => x"85",
           651 => x"32",
           652 => x"73",
           653 => x"58",
           654 => x"52",
           655 => x"09",
           656 => x"d3",
           657 => x"77",
           658 => x"70",
           659 => x"07",
           660 => x"55",
           661 => x"80",
           662 => x"38",
           663 => x"b2",
           664 => x"8e",
           665 => x"bb",
           666 => x"84",
           667 => x"ff",
           668 => x"84",
           669 => x"75",
           670 => x"57",
           671 => x"73",
           672 => x"30",
           673 => x"9f",
           674 => x"54",
           675 => x"24",
           676 => x"75",
           677 => x"71",
           678 => x"0c",
           679 => x"04",
           680 => x"bb",
           681 => x"3d",
           682 => x"3d",
           683 => x"86",
           684 => x"99",
           685 => x"56",
           686 => x"8e",
           687 => x"53",
           688 => x"3d",
           689 => x"9d",
           690 => x"54",
           691 => x"8d",
           692 => x"fd",
           693 => x"3d",
           694 => x"76",
           695 => x"85",
           696 => x"0d",
           697 => x"0d",
           698 => x"42",
           699 => x"70",
           700 => x"85",
           701 => x"81",
           702 => x"81",
           703 => x"5b",
           704 => x"7b",
           705 => x"06",
           706 => x"7b",
           707 => x"7b",
           708 => x"38",
           709 => x"81",
           710 => x"72",
           711 => x"81",
           712 => x"5f",
           713 => x"81",
           714 => x"b0",
           715 => x"70",
           716 => x"54",
           717 => x"38",
           718 => x"a9",
           719 => x"2a",
           720 => x"81",
           721 => x"7e",
           722 => x"38",
           723 => x"07",
           724 => x"57",
           725 => x"38",
           726 => x"54",
           727 => x"84",
           728 => x"0d",
           729 => x"2a",
           730 => x"10",
           731 => x"05",
           732 => x"70",
           733 => x"70",
           734 => x"29",
           735 => x"70",
           736 => x"5a",
           737 => x"80",
           738 => x"86",
           739 => x"06",
           740 => x"bd",
           741 => x"33",
           742 => x"fe",
           743 => x"b8",
           744 => x"2e",
           745 => x"93",
           746 => x"74",
           747 => x"8a",
           748 => x"5a",
           749 => x"38",
           750 => x"7c",
           751 => x"8b",
           752 => x"33",
           753 => x"cc",
           754 => x"39",
           755 => x"70",
           756 => x"55",
           757 => x"81",
           758 => x"40",
           759 => x"38",
           760 => x"72",
           761 => x"97",
           762 => x"10",
           763 => x"05",
           764 => x"04",
           765 => x"54",
           766 => x"73",
           767 => x"7c",
           768 => x"8a",
           769 => x"7c",
           770 => x"76",
           771 => x"fe",
           772 => x"ff",
           773 => x"39",
           774 => x"60",
           775 => x"08",
           776 => x"cf",
           777 => x"41",
           778 => x"94",
           779 => x"75",
           780 => x"3f",
           781 => x"08",
           782 => x"84",
           783 => x"18",
           784 => x"53",
           785 => x"88",
           786 => x"84",
           787 => x"55",
           788 => x"81",
           789 => x"79",
           790 => x"90",
           791 => x"bb",
           792 => x"84",
           793 => x"c5",
           794 => x"bb",
           795 => x"2b",
           796 => x"40",
           797 => x"2e",
           798 => x"84",
           799 => x"fc",
           800 => x"70",
           801 => x"55",
           802 => x"70",
           803 => x"5f",
           804 => x"9e",
           805 => x"80",
           806 => x"80",
           807 => x"79",
           808 => x"38",
           809 => x"80",
           810 => x"80",
           811 => x"90",
           812 => x"83",
           813 => x"06",
           814 => x"80",
           815 => x"75",
           816 => x"81",
           817 => x"54",
           818 => x"86",
           819 => x"83",
           820 => x"70",
           821 => x"86",
           822 => x"5b",
           823 => x"54",
           824 => x"85",
           825 => x"79",
           826 => x"70",
           827 => x"83",
           828 => x"59",
           829 => x"2e",
           830 => x"7a",
           831 => x"06",
           832 => x"eb",
           833 => x"2a",
           834 => x"73",
           835 => x"7a",
           836 => x"06",
           837 => x"97",
           838 => x"06",
           839 => x"8f",
           840 => x"2a",
           841 => x"7e",
           842 => x"38",
           843 => x"80",
           844 => x"80",
           845 => x"90",
           846 => x"54",
           847 => x"9d",
           848 => x"b0",
           849 => x"3f",
           850 => x"80",
           851 => x"80",
           852 => x"90",
           853 => x"54",
           854 => x"e5",
           855 => x"06",
           856 => x"2e",
           857 => x"79",
           858 => x"29",
           859 => x"05",
           860 => x"5b",
           861 => x"75",
           862 => x"7c",
           863 => x"87",
           864 => x"79",
           865 => x"29",
           866 => x"05",
           867 => x"5b",
           868 => x"80",
           869 => x"7a",
           870 => x"81",
           871 => x"7a",
           872 => x"b9",
           873 => x"e3",
           874 => x"38",
           875 => x"2e",
           876 => x"76",
           877 => x"81",
           878 => x"84",
           879 => x"96",
           880 => x"ff",
           881 => x"52",
           882 => x"3f",
           883 => x"94",
           884 => x"06",
           885 => x"81",
           886 => x"80",
           887 => x"38",
           888 => x"80",
           889 => x"80",
           890 => x"90",
           891 => x"55",
           892 => x"fc",
           893 => x"52",
           894 => x"f4",
           895 => x"7a",
           896 => x"7a",
           897 => x"33",
           898 => x"fa",
           899 => x"c8",
           900 => x"c0",
           901 => x"f8",
           902 => x"61",
           903 => x"08",
           904 => x"cf",
           905 => x"42",
           906 => x"fd",
           907 => x"84",
           908 => x"80",
           909 => x"13",
           910 => x"2b",
           911 => x"84",
           912 => x"fc",
           913 => x"70",
           914 => x"52",
           915 => x"41",
           916 => x"2a",
           917 => x"5c",
           918 => x"c9",
           919 => x"84",
           920 => x"fc",
           921 => x"70",
           922 => x"54",
           923 => x"25",
           924 => x"7c",
           925 => x"85",
           926 => x"39",
           927 => x"83",
           928 => x"5b",
           929 => x"ff",
           930 => x"ca",
           931 => x"75",
           932 => x"57",
           933 => x"d8",
           934 => x"ff",
           935 => x"ff",
           936 => x"54",
           937 => x"ff",
           938 => x"38",
           939 => x"70",
           940 => x"33",
           941 => x"3f",
           942 => x"fc",
           943 => x"fc",
           944 => x"84",
           945 => x"fc",
           946 => x"70",
           947 => x"58",
           948 => x"7b",
           949 => x"81",
           950 => x"57",
           951 => x"38",
           952 => x"7f",
           953 => x"71",
           954 => x"40",
           955 => x"7e",
           956 => x"38",
           957 => x"bf",
           958 => x"bb",
           959 => x"ad",
           960 => x"07",
           961 => x"5b",
           962 => x"38",
           963 => x"7a",
           964 => x"80",
           965 => x"59",
           966 => x"38",
           967 => x"7f",
           968 => x"71",
           969 => x"06",
           970 => x"5f",
           971 => x"38",
           972 => x"f6",
           973 => x"84",
           974 => x"ff",
           975 => x"31",
           976 => x"5a",
           977 => x"58",
           978 => x"7a",
           979 => x"7c",
           980 => x"76",
           981 => x"f7",
           982 => x"60",
           983 => x"08",
           984 => x"5d",
           985 => x"79",
           986 => x"75",
           987 => x"3f",
           988 => x"08",
           989 => x"06",
           990 => x"90",
           991 => x"c4",
           992 => x"80",
           993 => x"58",
           994 => x"88",
           995 => x"39",
           996 => x"80",
           997 => x"80",
           998 => x"90",
           999 => x"54",
          1000 => x"fa",
          1001 => x"52",
          1002 => x"c4",
          1003 => x"7c",
          1004 => x"83",
          1005 => x"90",
          1006 => x"06",
          1007 => x"7c",
          1008 => x"83",
          1009 => x"88",
          1010 => x"5f",
          1011 => x"fb",
          1012 => x"d8",
          1013 => x"2c",
          1014 => x"90",
          1015 => x"2c",
          1016 => x"06",
          1017 => x"53",
          1018 => x"38",
          1019 => x"7c",
          1020 => x"82",
          1021 => x"81",
          1022 => x"80",
          1023 => x"38",
          1024 => x"7c",
          1025 => x"2a",
          1026 => x"3f",
          1027 => x"5b",
          1028 => x"f7",
          1029 => x"c8",
          1030 => x"31",
          1031 => x"98",
          1032 => x"f9",
          1033 => x"52",
          1034 => x"c4",
          1035 => x"7c",
          1036 => x"82",
          1037 => x"be",
          1038 => x"75",
          1039 => x"3f",
          1040 => x"08",
          1041 => x"06",
          1042 => x"90",
          1043 => x"fd",
          1044 => x"82",
          1045 => x"71",
          1046 => x"06",
          1047 => x"fd",
          1048 => x"3d",
          1049 => x"e4",
          1050 => x"52",
          1051 => x"b5",
          1052 => x"0d",
          1053 => x"0d",
          1054 => x"0b",
          1055 => x"08",
          1056 => x"70",
          1057 => x"32",
          1058 => x"51",
          1059 => x"57",
          1060 => x"77",
          1061 => x"06",
          1062 => x"74",
          1063 => x"56",
          1064 => x"77",
          1065 => x"84",
          1066 => x"52",
          1067 => x"14",
          1068 => x"2d",
          1069 => x"08",
          1070 => x"38",
          1071 => x"70",
          1072 => x"33",
          1073 => x"2e",
          1074 => x"e6",
          1075 => x"d7",
          1076 => x"e8",
          1077 => x"e6",
          1078 => x"8a",
          1079 => x"08",
          1080 => x"84",
          1081 => x"80",
          1082 => x"ff",
          1083 => x"75",
          1084 => x"0c",
          1085 => x"04",
          1086 => x"78",
          1087 => x"80",
          1088 => x"33",
          1089 => x"81",
          1090 => x"06",
          1091 => x"57",
          1092 => x"77",
          1093 => x"06",
          1094 => x"70",
          1095 => x"33",
          1096 => x"2e",
          1097 => x"98",
          1098 => x"75",
          1099 => x"0c",
          1100 => x"04",
          1101 => x"05",
          1102 => x"72",
          1103 => x"38",
          1104 => x"51",
          1105 => x"53",
          1106 => x"bb",
          1107 => x"2e",
          1108 => x"74",
          1109 => x"56",
          1110 => x"72",
          1111 => x"39",
          1112 => x"84",
          1113 => x"52",
          1114 => x"3f",
          1115 => x"04",
          1116 => x"78",
          1117 => x"33",
          1118 => x"81",
          1119 => x"56",
          1120 => x"ff",
          1121 => x"38",
          1122 => x"81",
          1123 => x"80",
          1124 => x"8c",
          1125 => x"72",
          1126 => x"25",
          1127 => x"08",
          1128 => x"34",
          1129 => x"05",
          1130 => x"15",
          1131 => x"13",
          1132 => x"76",
          1133 => x"bb",
          1134 => x"3d",
          1135 => x"52",
          1136 => x"06",
          1137 => x"08",
          1138 => x"ff",
          1139 => x"84",
          1140 => x"8c",
          1141 => x"05",
          1142 => x"76",
          1143 => x"fb",
          1144 => x"85",
          1145 => x"81",
          1146 => x"81",
          1147 => x"55",
          1148 => x"ff",
          1149 => x"38",
          1150 => x"81",
          1151 => x"b3",
          1152 => x"2a",
          1153 => x"71",
          1154 => x"c3",
          1155 => x"70",
          1156 => x"71",
          1157 => x"f0",
          1158 => x"76",
          1159 => x"08",
          1160 => x"17",
          1161 => x"ff",
          1162 => x"84",
          1163 => x"87",
          1164 => x"74",
          1165 => x"53",
          1166 => x"34",
          1167 => x"81",
          1168 => x"0c",
          1169 => x"84",
          1170 => x"87",
          1171 => x"75",
          1172 => x"08",
          1173 => x"84",
          1174 => x"52",
          1175 => x"08",
          1176 => x"b9",
          1177 => x"33",
          1178 => x"54",
          1179 => x"84",
          1180 => x"85",
          1181 => x"07",
          1182 => x"17",
          1183 => x"73",
          1184 => x"0c",
          1185 => x"04",
          1186 => x"53",
          1187 => x"34",
          1188 => x"39",
          1189 => x"75",
          1190 => x"54",
          1191 => x"81",
          1192 => x"51",
          1193 => x"ff",
          1194 => x"70",
          1195 => x"33",
          1196 => x"70",
          1197 => x"34",
          1198 => x"73",
          1199 => x"0c",
          1200 => x"04",
          1201 => x"76",
          1202 => x"55",
          1203 => x"70",
          1204 => x"38",
          1205 => x"a1",
          1206 => x"2e",
          1207 => x"70",
          1208 => x"33",
          1209 => x"05",
          1210 => x"11",
          1211 => x"38",
          1212 => x"84",
          1213 => x"0d",
          1214 => x"55",
          1215 => x"d9",
          1216 => x"75",
          1217 => x"13",
          1218 => x"53",
          1219 => x"34",
          1220 => x"70",
          1221 => x"38",
          1222 => x"13",
          1223 => x"33",
          1224 => x"11",
          1225 => x"38",
          1226 => x"3d",
          1227 => x"53",
          1228 => x"81",
          1229 => x"51",
          1230 => x"ff",
          1231 => x"31",
          1232 => x"0c",
          1233 => x"0d",
          1234 => x"0d",
          1235 => x"54",
          1236 => x"70",
          1237 => x"33",
          1238 => x"70",
          1239 => x"34",
          1240 => x"73",
          1241 => x"0c",
          1242 => x"04",
          1243 => x"75",
          1244 => x"55",
          1245 => x"70",
          1246 => x"38",
          1247 => x"05",
          1248 => x"70",
          1249 => x"34",
          1250 => x"70",
          1251 => x"84",
          1252 => x"85",
          1253 => x"fc",
          1254 => x"78",
          1255 => x"54",
          1256 => x"a1",
          1257 => x"75",
          1258 => x"57",
          1259 => x"71",
          1260 => x"81",
          1261 => x"81",
          1262 => x"80",
          1263 => x"ff",
          1264 => x"e1",
          1265 => x"70",
          1266 => x"0c",
          1267 => x"04",
          1268 => x"f1",
          1269 => x"53",
          1270 => x"80",
          1271 => x"ff",
          1272 => x"81",
          1273 => x"2e",
          1274 => x"72",
          1275 => x"84",
          1276 => x"0d",
          1277 => x"bb",
          1278 => x"3d",
          1279 => x"3d",
          1280 => x"53",
          1281 => x"80",
          1282 => x"bb",
          1283 => x"bb",
          1284 => x"05",
          1285 => x"b4",
          1286 => x"bb",
          1287 => x"84",
          1288 => x"80",
          1289 => x"84",
          1290 => x"15",
          1291 => x"34",
          1292 => x"52",
          1293 => x"08",
          1294 => x"3f",
          1295 => x"08",
          1296 => x"bb",
          1297 => x"3d",
          1298 => x"3d",
          1299 => x"71",
          1300 => x"53",
          1301 => x"2e",
          1302 => x"70",
          1303 => x"33",
          1304 => x"2e",
          1305 => x"12",
          1306 => x"2e",
          1307 => x"ea",
          1308 => x"70",
          1309 => x"52",
          1310 => x"84",
          1311 => x"0d",
          1312 => x"0d",
          1313 => x"72",
          1314 => x"54",
          1315 => x"8e",
          1316 => x"70",
          1317 => x"34",
          1318 => x"70",
          1319 => x"84",
          1320 => x"85",
          1321 => x"fa",
          1322 => x"7a",
          1323 => x"52",
          1324 => x"8b",
          1325 => x"80",
          1326 => x"bb",
          1327 => x"e0",
          1328 => x"80",
          1329 => x"73",
          1330 => x"3f",
          1331 => x"84",
          1332 => x"80",
          1333 => x"26",
          1334 => x"73",
          1335 => x"2e",
          1336 => x"81",
          1337 => x"2a",
          1338 => x"76",
          1339 => x"54",
          1340 => x"56",
          1341 => x"a8",
          1342 => x"74",
          1343 => x"74",
          1344 => x"78",
          1345 => x"11",
          1346 => x"81",
          1347 => x"06",
          1348 => x"ff",
          1349 => x"52",
          1350 => x"55",
          1351 => x"38",
          1352 => x"07",
          1353 => x"bb",
          1354 => x"3d",
          1355 => x"3d",
          1356 => x"fc",
          1357 => x"70",
          1358 => x"07",
          1359 => x"84",
          1360 => x"31",
          1361 => x"70",
          1362 => x"06",
          1363 => x"80",
          1364 => x"88",
          1365 => x"71",
          1366 => x"f0",
          1367 => x"70",
          1368 => x"2b",
          1369 => x"74",
          1370 => x"53",
          1371 => x"73",
          1372 => x"30",
          1373 => x"10",
          1374 => x"77",
          1375 => x"81",
          1376 => x"70",
          1377 => x"30",
          1378 => x"06",
          1379 => x"84",
          1380 => x"51",
          1381 => x"51",
          1382 => x"53",
          1383 => x"51",
          1384 => x"56",
          1385 => x"54",
          1386 => x"0d",
          1387 => x"0d",
          1388 => x"54",
          1389 => x"54",
          1390 => x"84",
          1391 => x"73",
          1392 => x"31",
          1393 => x"0c",
          1394 => x"0d",
          1395 => x"0d",
          1396 => x"54",
          1397 => x"80",
          1398 => x"76",
          1399 => x"3f",
          1400 => x"08",
          1401 => x"52",
          1402 => x"8d",
          1403 => x"fe",
          1404 => x"84",
          1405 => x"31",
          1406 => x"71",
          1407 => x"c5",
          1408 => x"71",
          1409 => x"38",
          1410 => x"71",
          1411 => x"31",
          1412 => x"57",
          1413 => x"80",
          1414 => x"2e",
          1415 => x"10",
          1416 => x"07",
          1417 => x"07",
          1418 => x"ff",
          1419 => x"70",
          1420 => x"72",
          1421 => x"31",
          1422 => x"56",
          1423 => x"58",
          1424 => x"da",
          1425 => x"bb",
          1426 => x"3d",
          1427 => x"3d",
          1428 => x"2c",
          1429 => x"7a",
          1430 => x"32",
          1431 => x"7d",
          1432 => x"32",
          1433 => x"57",
          1434 => x"56",
          1435 => x"55",
          1436 => x"3f",
          1437 => x"08",
          1438 => x"31",
          1439 => x"0c",
          1440 => x"04",
          1441 => x"7b",
          1442 => x"80",
          1443 => x"77",
          1444 => x"56",
          1445 => x"a0",
          1446 => x"06",
          1447 => x"15",
          1448 => x"70",
          1449 => x"73",
          1450 => x"38",
          1451 => x"80",
          1452 => x"b0",
          1453 => x"38",
          1454 => x"80",
          1455 => x"26",
          1456 => x"8a",
          1457 => x"a0",
          1458 => x"c4",
          1459 => x"74",
          1460 => x"e0",
          1461 => x"ff",
          1462 => x"d0",
          1463 => x"ff",
          1464 => x"90",
          1465 => x"38",
          1466 => x"81",
          1467 => x"54",
          1468 => x"81",
          1469 => x"78",
          1470 => x"38",
          1471 => x"13",
          1472 => x"79",
          1473 => x"56",
          1474 => x"a0",
          1475 => x"38",
          1476 => x"84",
          1477 => x"56",
          1478 => x"81",
          1479 => x"bb",
          1480 => x"3d",
          1481 => x"70",
          1482 => x"0c",
          1483 => x"56",
          1484 => x"2e",
          1485 => x"fe",
          1486 => x"15",
          1487 => x"70",
          1488 => x"73",
          1489 => x"a6",
          1490 => x"73",
          1491 => x"a0",
          1492 => x"a0",
          1493 => x"38",
          1494 => x"80",
          1495 => x"89",
          1496 => x"e1",
          1497 => x"bb",
          1498 => x"3d",
          1499 => x"58",
          1500 => x"78",
          1501 => x"55",
          1502 => x"fe",
          1503 => x"0b",
          1504 => x"0c",
          1505 => x"04",
          1506 => x"7b",
          1507 => x"80",
          1508 => x"77",
          1509 => x"56",
          1510 => x"a0",
          1511 => x"06",
          1512 => x"15",
          1513 => x"70",
          1514 => x"73",
          1515 => x"38",
          1516 => x"80",
          1517 => x"b0",
          1518 => x"38",
          1519 => x"80",
          1520 => x"26",
          1521 => x"8a",
          1522 => x"a0",
          1523 => x"c4",
          1524 => x"74",
          1525 => x"e0",
          1526 => x"ff",
          1527 => x"d0",
          1528 => x"ff",
          1529 => x"90",
          1530 => x"38",
          1531 => x"81",
          1532 => x"54",
          1533 => x"81",
          1534 => x"78",
          1535 => x"38",
          1536 => x"13",
          1537 => x"79",
          1538 => x"56",
          1539 => x"a0",
          1540 => x"38",
          1541 => x"84",
          1542 => x"56",
          1543 => x"81",
          1544 => x"bb",
          1545 => x"3d",
          1546 => x"70",
          1547 => x"0c",
          1548 => x"56",
          1549 => x"2e",
          1550 => x"fe",
          1551 => x"15",
          1552 => x"70",
          1553 => x"73",
          1554 => x"a6",
          1555 => x"73",
          1556 => x"a0",
          1557 => x"a0",
          1558 => x"38",
          1559 => x"80",
          1560 => x"89",
          1561 => x"e1",
          1562 => x"bb",
          1563 => x"3d",
          1564 => x"58",
          1565 => x"78",
          1566 => x"55",
          1567 => x"fe",
          1568 => x"0b",
          1569 => x"0c",
          1570 => x"04",
          1571 => x"3f",
          1572 => x"08",
          1573 => x"84",
          1574 => x"04",
          1575 => x"73",
          1576 => x"26",
          1577 => x"10",
          1578 => x"94",
          1579 => x"08",
          1580 => x"ac",
          1581 => x"3f",
          1582 => x"04",
          1583 => x"51",
          1584 => x"83",
          1585 => x"83",
          1586 => x"ef",
          1587 => x"3d",
          1588 => x"cf",
          1589 => x"9d",
          1590 => x"0d",
          1591 => x"84",
          1592 => x"3f",
          1593 => x"04",
          1594 => x"51",
          1595 => x"83",
          1596 => x"83",
          1597 => x"ee",
          1598 => x"3d",
          1599 => x"d0",
          1600 => x"f1",
          1601 => x"0d",
          1602 => x"ec",
          1603 => x"3f",
          1604 => x"04",
          1605 => x"51",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ee",
          1609 => x"3d",
          1610 => x"d1",
          1611 => x"c5",
          1612 => x"0d",
          1613 => x"cc",
          1614 => x"3f",
          1615 => x"04",
          1616 => x"51",
          1617 => x"83",
          1618 => x"83",
          1619 => x"ee",
          1620 => x"3d",
          1621 => x"d2",
          1622 => x"99",
          1623 => x"0d",
          1624 => x"98",
          1625 => x"3f",
          1626 => x"04",
          1627 => x"51",
          1628 => x"83",
          1629 => x"83",
          1630 => x"ed",
          1631 => x"3d",
          1632 => x"d2",
          1633 => x"ed",
          1634 => x"0d",
          1635 => x"d4",
          1636 => x"3f",
          1637 => x"04",
          1638 => x"0d",
          1639 => x"08",
          1640 => x"84",
          1641 => x"5b",
          1642 => x"81",
          1643 => x"79",
          1644 => x"07",
          1645 => x"57",
          1646 => x"57",
          1647 => x"26",
          1648 => x"57",
          1649 => x"70",
          1650 => x"51",
          1651 => x"74",
          1652 => x"81",
          1653 => x"8c",
          1654 => x"58",
          1655 => x"3f",
          1656 => x"08",
          1657 => x"84",
          1658 => x"80",
          1659 => x"51",
          1660 => x"3f",
          1661 => x"78",
          1662 => x"7b",
          1663 => x"2a",
          1664 => x"57",
          1665 => x"80",
          1666 => x"87",
          1667 => x"08",
          1668 => x"e7",
          1669 => x"38",
          1670 => x"87",
          1671 => x"f5",
          1672 => x"bb",
          1673 => x"83",
          1674 => x"78",
          1675 => x"e0",
          1676 => x"3f",
          1677 => x"84",
          1678 => x"3d",
          1679 => x"bb",
          1680 => x"c0",
          1681 => x"84",
          1682 => x"59",
          1683 => x"fb",
          1684 => x"84",
          1685 => x"52",
          1686 => x"9f",
          1687 => x"bb",
          1688 => x"84",
          1689 => x"ff",
          1690 => x"55",
          1691 => x"fe",
          1692 => x"19",
          1693 => x"59",
          1694 => x"e8",
          1695 => x"f4",
          1696 => x"bb",
          1697 => x"78",
          1698 => x"3f",
          1699 => x"08",
          1700 => x"84",
          1701 => x"83",
          1702 => x"de",
          1703 => x"94",
          1704 => x"0d",
          1705 => x"05",
          1706 => x"58",
          1707 => x"80",
          1708 => x"7a",
          1709 => x"3f",
          1710 => x"08",
          1711 => x"80",
          1712 => x"76",
          1713 => x"38",
          1714 => x"84",
          1715 => x"0d",
          1716 => x"84",
          1717 => x"61",
          1718 => x"84",
          1719 => x"7f",
          1720 => x"78",
          1721 => x"84",
          1722 => x"84",
          1723 => x"0d",
          1724 => x"0d",
          1725 => x"02",
          1726 => x"cf",
          1727 => x"73",
          1728 => x"5f",
          1729 => x"5d",
          1730 => x"2e",
          1731 => x"7a",
          1732 => x"8c",
          1733 => x"3f",
          1734 => x"51",
          1735 => x"80",
          1736 => x"27",
          1737 => x"90",
          1738 => x"38",
          1739 => x"82",
          1740 => x"18",
          1741 => x"27",
          1742 => x"72",
          1743 => x"d3",
          1744 => x"c6",
          1745 => x"84",
          1746 => x"53",
          1747 => x"ec",
          1748 => x"74",
          1749 => x"83",
          1750 => x"dd",
          1751 => x"56",
          1752 => x"80",
          1753 => x"18",
          1754 => x"53",
          1755 => x"7a",
          1756 => x"81",
          1757 => x"9f",
          1758 => x"38",
          1759 => x"73",
          1760 => x"ff",
          1761 => x"74",
          1762 => x"38",
          1763 => x"27",
          1764 => x"84",
          1765 => x"52",
          1766 => x"d4",
          1767 => x"56",
          1768 => x"c2",
          1769 => x"a4",
          1770 => x"3f",
          1771 => x"1c",
          1772 => x"51",
          1773 => x"84",
          1774 => x"98",
          1775 => x"2c",
          1776 => x"a0",
          1777 => x"38",
          1778 => x"82",
          1779 => x"1e",
          1780 => x"26",
          1781 => x"ff",
          1782 => x"84",
          1783 => x"0d",
          1784 => x"a8",
          1785 => x"3f",
          1786 => x"e6",
          1787 => x"54",
          1788 => x"fc",
          1789 => x"26",
          1790 => x"fe",
          1791 => x"d3",
          1792 => x"86",
          1793 => x"84",
          1794 => x"53",
          1795 => x"ea",
          1796 => x"79",
          1797 => x"38",
          1798 => x"72",
          1799 => x"38",
          1800 => x"83",
          1801 => x"db",
          1802 => x"14",
          1803 => x"08",
          1804 => x"51",
          1805 => x"78",
          1806 => x"38",
          1807 => x"83",
          1808 => x"db",
          1809 => x"14",
          1810 => x"08",
          1811 => x"51",
          1812 => x"73",
          1813 => x"ff",
          1814 => x"53",
          1815 => x"df",
          1816 => x"52",
          1817 => x"51",
          1818 => x"84",
          1819 => x"e8",
          1820 => x"a0",
          1821 => x"3f",
          1822 => x"dd",
          1823 => x"39",
          1824 => x"08",
          1825 => x"e9",
          1826 => x"16",
          1827 => x"39",
          1828 => x"3f",
          1829 => x"08",
          1830 => x"53",
          1831 => x"a8",
          1832 => x"38",
          1833 => x"80",
          1834 => x"81",
          1835 => x"38",
          1836 => x"db",
          1837 => x"9b",
          1838 => x"bb",
          1839 => x"2b",
          1840 => x"70",
          1841 => x"30",
          1842 => x"70",
          1843 => x"07",
          1844 => x"06",
          1845 => x"59",
          1846 => x"72",
          1847 => x"e8",
          1848 => x"9b",
          1849 => x"bb",
          1850 => x"2b",
          1851 => x"70",
          1852 => x"30",
          1853 => x"70",
          1854 => x"07",
          1855 => x"06",
          1856 => x"59",
          1857 => x"80",
          1858 => x"a9",
          1859 => x"39",
          1860 => x"bb",
          1861 => x"3d",
          1862 => x"3d",
          1863 => x"96",
          1864 => x"aa",
          1865 => x"51",
          1866 => x"83",
          1867 => x"9d",
          1868 => x"51",
          1869 => x"72",
          1870 => x"81",
          1871 => x"71",
          1872 => x"72",
          1873 => x"81",
          1874 => x"71",
          1875 => x"72",
          1876 => x"81",
          1877 => x"71",
          1878 => x"72",
          1879 => x"81",
          1880 => x"71",
          1881 => x"72",
          1882 => x"81",
          1883 => x"71",
          1884 => x"72",
          1885 => x"81",
          1886 => x"71",
          1887 => x"72",
          1888 => x"81",
          1889 => x"71",
          1890 => x"88",
          1891 => x"53",
          1892 => x"a9",
          1893 => x"3d",
          1894 => x"51",
          1895 => x"83",
          1896 => x"9c",
          1897 => x"51",
          1898 => x"a9",
          1899 => x"3d",
          1900 => x"51",
          1901 => x"83",
          1902 => x"9c",
          1903 => x"51",
          1904 => x"72",
          1905 => x"06",
          1906 => x"2e",
          1907 => x"39",
          1908 => x"e3",
          1909 => x"90",
          1910 => x"3f",
          1911 => x"d7",
          1912 => x"2a",
          1913 => x"51",
          1914 => x"2e",
          1915 => x"c2",
          1916 => x"9b",
          1917 => x"d5",
          1918 => x"d3",
          1919 => x"9b",
          1920 => x"86",
          1921 => x"06",
          1922 => x"80",
          1923 => x"38",
          1924 => x"81",
          1925 => x"3f",
          1926 => x"51",
          1927 => x"80",
          1928 => x"3f",
          1929 => x"70",
          1930 => x"52",
          1931 => x"fe",
          1932 => x"bd",
          1933 => x"9a",
          1934 => x"d5",
          1935 => x"8f",
          1936 => x"9a",
          1937 => x"84",
          1938 => x"06",
          1939 => x"80",
          1940 => x"38",
          1941 => x"81",
          1942 => x"3f",
          1943 => x"51",
          1944 => x"80",
          1945 => x"3f",
          1946 => x"70",
          1947 => x"52",
          1948 => x"fd",
          1949 => x"bd",
          1950 => x"9a",
          1951 => x"d5",
          1952 => x"cb",
          1953 => x"9a",
          1954 => x"82",
          1955 => x"06",
          1956 => x"80",
          1957 => x"38",
          1958 => x"ca",
          1959 => x"70",
          1960 => x"61",
          1961 => x"0c",
          1962 => x"60",
          1963 => x"c9",
          1964 => x"84",
          1965 => x"06",
          1966 => x"59",
          1967 => x"84",
          1968 => x"d6",
          1969 => x"ad",
          1970 => x"43",
          1971 => x"51",
          1972 => x"7e",
          1973 => x"53",
          1974 => x"51",
          1975 => x"0b",
          1976 => x"f8",
          1977 => x"ff",
          1978 => x"79",
          1979 => x"f1",
          1980 => x"2e",
          1981 => x"78",
          1982 => x"5e",
          1983 => x"83",
          1984 => x"70",
          1985 => x"80",
          1986 => x"38",
          1987 => x"7b",
          1988 => x"81",
          1989 => x"81",
          1990 => x"5d",
          1991 => x"2e",
          1992 => x"5c",
          1993 => x"be",
          1994 => x"29",
          1995 => x"05",
          1996 => x"5b",
          1997 => x"84",
          1998 => x"84",
          1999 => x"54",
          2000 => x"08",
          2001 => x"cf",
          2002 => x"84",
          2003 => x"84",
          2004 => x"7d",
          2005 => x"84",
          2006 => x"70",
          2007 => x"5d",
          2008 => x"27",
          2009 => x"3d",
          2010 => x"80",
          2011 => x"38",
          2012 => x"7e",
          2013 => x"3f",
          2014 => x"08",
          2015 => x"84",
          2016 => x"8d",
          2017 => x"bb",
          2018 => x"b8",
          2019 => x"05",
          2020 => x"3f",
          2021 => x"08",
          2022 => x"5c",
          2023 => x"2e",
          2024 => x"84",
          2025 => x"51",
          2026 => x"84",
          2027 => x"8f",
          2028 => x"38",
          2029 => x"3d",
          2030 => x"82",
          2031 => x"38",
          2032 => x"8c",
          2033 => x"81",
          2034 => x"38",
          2035 => x"53",
          2036 => x"52",
          2037 => x"d2",
          2038 => x"c0",
          2039 => x"b4",
          2040 => x"67",
          2041 => x"90",
          2042 => x"90",
          2043 => x"7c",
          2044 => x"3f",
          2045 => x"08",
          2046 => x"08",
          2047 => x"70",
          2048 => x"25",
          2049 => x"42",
          2050 => x"83",
          2051 => x"81",
          2052 => x"06",
          2053 => x"2e",
          2054 => x"1b",
          2055 => x"06",
          2056 => x"ff",
          2057 => x"81",
          2058 => x"32",
          2059 => x"81",
          2060 => x"ff",
          2061 => x"38",
          2062 => x"96",
          2063 => x"d6",
          2064 => x"c6",
          2065 => x"80",
          2066 => x"52",
          2067 => x"b1",
          2068 => x"83",
          2069 => x"70",
          2070 => x"5b",
          2071 => x"91",
          2072 => x"83",
          2073 => x"84",
          2074 => x"82",
          2075 => x"84",
          2076 => x"80",
          2077 => x"0b",
          2078 => x"ef",
          2079 => x"de",
          2080 => x"f8",
          2081 => x"82",
          2082 => x"84",
          2083 => x"80",
          2084 => x"84",
          2085 => x"51",
          2086 => x"0b",
          2087 => x"f8",
          2088 => x"ff",
          2089 => x"7d",
          2090 => x"81",
          2091 => x"38",
          2092 => x"de",
          2093 => x"a1",
          2094 => x"0b",
          2095 => x"ef",
          2096 => x"55",
          2097 => x"54",
          2098 => x"f8",
          2099 => x"a7",
          2100 => x"70",
          2101 => x"fc",
          2102 => x"39",
          2103 => x"0c",
          2104 => x"59",
          2105 => x"26",
          2106 => x"78",
          2107 => x"bf",
          2108 => x"79",
          2109 => x"53",
          2110 => x"52",
          2111 => x"ec",
          2112 => x"7e",
          2113 => x"b0",
          2114 => x"bd",
          2115 => x"84",
          2116 => x"09",
          2117 => x"aa",
          2118 => x"9a",
          2119 => x"41",
          2120 => x"83",
          2121 => x"de",
          2122 => x"51",
          2123 => x"3f",
          2124 => x"83",
          2125 => x"7b",
          2126 => x"a0",
          2127 => x"83",
          2128 => x"7c",
          2129 => x"3f",
          2130 => x"81",
          2131 => x"fa",
          2132 => x"f9",
          2133 => x"39",
          2134 => x"51",
          2135 => x"3f",
          2136 => x"81",
          2137 => x"fa",
          2138 => x"d7",
          2139 => x"85",
          2140 => x"78",
          2141 => x"c8",
          2142 => x"3f",
          2143 => x"fa",
          2144 => x"3d",
          2145 => x"53",
          2146 => x"51",
          2147 => x"84",
          2148 => x"80",
          2149 => x"38",
          2150 => x"d7",
          2151 => x"ea",
          2152 => x"79",
          2153 => x"84",
          2154 => x"fa",
          2155 => x"bb",
          2156 => x"83",
          2157 => x"d0",
          2158 => x"90",
          2159 => x"ff",
          2160 => x"ff",
          2161 => x"eb",
          2162 => x"bb",
          2163 => x"2e",
          2164 => x"68",
          2165 => x"9c",
          2166 => x"3f",
          2167 => x"04",
          2168 => x"f4",
          2169 => x"80",
          2170 => x"98",
          2171 => x"84",
          2172 => x"f9",
          2173 => x"3d",
          2174 => x"53",
          2175 => x"51",
          2176 => x"84",
          2177 => x"86",
          2178 => x"59",
          2179 => x"78",
          2180 => x"b8",
          2181 => x"3f",
          2182 => x"08",
          2183 => x"52",
          2184 => x"81",
          2185 => x"7e",
          2186 => x"ae",
          2187 => x"38",
          2188 => x"87",
          2189 => x"84",
          2190 => x"59",
          2191 => x"3d",
          2192 => x"53",
          2193 => x"51",
          2194 => x"84",
          2195 => x"80",
          2196 => x"38",
          2197 => x"f0",
          2198 => x"80",
          2199 => x"a4",
          2200 => x"84",
          2201 => x"38",
          2202 => x"22",
          2203 => x"83",
          2204 => x"cf",
          2205 => x"e6",
          2206 => x"80",
          2207 => x"51",
          2208 => x"7e",
          2209 => x"59",
          2210 => x"f8",
          2211 => x"9f",
          2212 => x"38",
          2213 => x"70",
          2214 => x"39",
          2215 => x"84",
          2216 => x"80",
          2217 => x"e0",
          2218 => x"84",
          2219 => x"f8",
          2220 => x"3d",
          2221 => x"53",
          2222 => x"51",
          2223 => x"84",
          2224 => x"80",
          2225 => x"38",
          2226 => x"f8",
          2227 => x"80",
          2228 => x"b4",
          2229 => x"84",
          2230 => x"f7",
          2231 => x"d8",
          2232 => x"a6",
          2233 => x"5d",
          2234 => x"27",
          2235 => x"65",
          2236 => x"33",
          2237 => x"7a",
          2238 => x"38",
          2239 => x"54",
          2240 => x"78",
          2241 => x"e4",
          2242 => x"3f",
          2243 => x"5c",
          2244 => x"1b",
          2245 => x"39",
          2246 => x"84",
          2247 => x"80",
          2248 => x"e4",
          2249 => x"84",
          2250 => x"f7",
          2251 => x"3d",
          2252 => x"53",
          2253 => x"51",
          2254 => x"84",
          2255 => x"80",
          2256 => x"38",
          2257 => x"f8",
          2258 => x"80",
          2259 => x"b8",
          2260 => x"84",
          2261 => x"f6",
          2262 => x"d9",
          2263 => x"aa",
          2264 => x"79",
          2265 => x"93",
          2266 => x"79",
          2267 => x"5b",
          2268 => x"65",
          2269 => x"eb",
          2270 => x"ff",
          2271 => x"ff",
          2272 => x"e8",
          2273 => x"bb",
          2274 => x"2e",
          2275 => x"b8",
          2276 => x"11",
          2277 => x"05",
          2278 => x"3f",
          2279 => x"08",
          2280 => x"70",
          2281 => x"83",
          2282 => x"cc",
          2283 => x"e6",
          2284 => x"80",
          2285 => x"51",
          2286 => x"7e",
          2287 => x"59",
          2288 => x"f6",
          2289 => x"9f",
          2290 => x"38",
          2291 => x"49",
          2292 => x"59",
          2293 => x"05",
          2294 => x"68",
          2295 => x"b8",
          2296 => x"11",
          2297 => x"05",
          2298 => x"3f",
          2299 => x"08",
          2300 => x"d8",
          2301 => x"02",
          2302 => x"33",
          2303 => x"81",
          2304 => x"3d",
          2305 => x"53",
          2306 => x"51",
          2307 => x"84",
          2308 => x"ff",
          2309 => x"b4",
          2310 => x"ff",
          2311 => x"ff",
          2312 => x"e6",
          2313 => x"bb",
          2314 => x"2e",
          2315 => x"b8",
          2316 => x"11",
          2317 => x"05",
          2318 => x"3f",
          2319 => x"08",
          2320 => x"88",
          2321 => x"fe",
          2322 => x"ff",
          2323 => x"e6",
          2324 => x"bb",
          2325 => x"38",
          2326 => x"08",
          2327 => x"98",
          2328 => x"3f",
          2329 => x"59",
          2330 => x"8f",
          2331 => x"7a",
          2332 => x"05",
          2333 => x"79",
          2334 => x"8a",
          2335 => x"3f",
          2336 => x"b8",
          2337 => x"05",
          2338 => x"3f",
          2339 => x"08",
          2340 => x"80",
          2341 => x"88",
          2342 => x"53",
          2343 => x"08",
          2344 => x"e9",
          2345 => x"bb",
          2346 => x"2e",
          2347 => x"84",
          2348 => x"51",
          2349 => x"f4",
          2350 => x"3d",
          2351 => x"53",
          2352 => x"51",
          2353 => x"84",
          2354 => x"91",
          2355 => x"88",
          2356 => x"80",
          2357 => x"38",
          2358 => x"08",
          2359 => x"fe",
          2360 => x"ff",
          2361 => x"e5",
          2362 => x"bb",
          2363 => x"38",
          2364 => x"33",
          2365 => x"2e",
          2366 => x"83",
          2367 => x"47",
          2368 => x"f8",
          2369 => x"80",
          2370 => x"fc",
          2371 => x"84",
          2372 => x"a5",
          2373 => x"5c",
          2374 => x"2e",
          2375 => x"5c",
          2376 => x"70",
          2377 => x"07",
          2378 => x"06",
          2379 => x"79",
          2380 => x"38",
          2381 => x"83",
          2382 => x"83",
          2383 => x"d6",
          2384 => x"55",
          2385 => x"53",
          2386 => x"51",
          2387 => x"83",
          2388 => x"d6",
          2389 => x"f4",
          2390 => x"71",
          2391 => x"84",
          2392 => x"3d",
          2393 => x"53",
          2394 => x"51",
          2395 => x"84",
          2396 => x"80",
          2397 => x"38",
          2398 => x"0c",
          2399 => x"05",
          2400 => x"fe",
          2401 => x"ff",
          2402 => x"e1",
          2403 => x"bb",
          2404 => x"38",
          2405 => x"64",
          2406 => x"ce",
          2407 => x"70",
          2408 => x"23",
          2409 => x"3d",
          2410 => x"53",
          2411 => x"51",
          2412 => x"84",
          2413 => x"80",
          2414 => x"38",
          2415 => x"80",
          2416 => x"7e",
          2417 => x"40",
          2418 => x"b8",
          2419 => x"11",
          2420 => x"05",
          2421 => x"3f",
          2422 => x"08",
          2423 => x"f1",
          2424 => x"3d",
          2425 => x"53",
          2426 => x"51",
          2427 => x"84",
          2428 => x"80",
          2429 => x"38",
          2430 => x"80",
          2431 => x"7c",
          2432 => x"05",
          2433 => x"39",
          2434 => x"f0",
          2435 => x"80",
          2436 => x"f0",
          2437 => x"84",
          2438 => x"81",
          2439 => x"64",
          2440 => x"64",
          2441 => x"46",
          2442 => x"39",
          2443 => x"09",
          2444 => x"98",
          2445 => x"83",
          2446 => x"80",
          2447 => x"c0",
          2448 => x"c8",
          2449 => x"91",
          2450 => x"7c",
          2451 => x"3f",
          2452 => x"83",
          2453 => x"d4",
          2454 => x"f0",
          2455 => x"fe",
          2456 => x"ff",
          2457 => x"e0",
          2458 => x"bb",
          2459 => x"2e",
          2460 => x"59",
          2461 => x"05",
          2462 => x"82",
          2463 => x"78",
          2464 => x"39",
          2465 => x"33",
          2466 => x"2e",
          2467 => x"83",
          2468 => x"47",
          2469 => x"83",
          2470 => x"5c",
          2471 => x"a1",
          2472 => x"c8",
          2473 => x"b5",
          2474 => x"f8",
          2475 => x"3f",
          2476 => x"b6",
          2477 => x"f8",
          2478 => x"3f",
          2479 => x"cc",
          2480 => x"8a",
          2481 => x"80",
          2482 => x"83",
          2483 => x"49",
          2484 => x"83",
          2485 => x"d3",
          2486 => x"c6",
          2487 => x"8a",
          2488 => x"80",
          2489 => x"83",
          2490 => x"47",
          2491 => x"83",
          2492 => x"5e",
          2493 => x"9b",
          2494 => x"d8",
          2495 => x"dd",
          2496 => x"8b",
          2497 => x"80",
          2498 => x"83",
          2499 => x"47",
          2500 => x"83",
          2501 => x"5d",
          2502 => x"9b",
          2503 => x"e0",
          2504 => x"b9",
          2505 => x"86",
          2506 => x"80",
          2507 => x"83",
          2508 => x"47",
          2509 => x"83",
          2510 => x"fc",
          2511 => x"fb",
          2512 => x"f3",
          2513 => x"05",
          2514 => x"39",
          2515 => x"80",
          2516 => x"b4",
          2517 => x"94",
          2518 => x"56",
          2519 => x"80",
          2520 => x"da",
          2521 => x"bb",
          2522 => x"2b",
          2523 => x"55",
          2524 => x"52",
          2525 => x"af",
          2526 => x"bb",
          2527 => x"77",
          2528 => x"94",
          2529 => x"56",
          2530 => x"80",
          2531 => x"da",
          2532 => x"bb",
          2533 => x"2b",
          2534 => x"55",
          2535 => x"52",
          2536 => x"83",
          2537 => x"bb",
          2538 => x"77",
          2539 => x"83",
          2540 => x"94",
          2541 => x"80",
          2542 => x"c0",
          2543 => x"81",
          2544 => x"81",
          2545 => x"83",
          2546 => x"a1",
          2547 => x"5e",
          2548 => x"0b",
          2549 => x"88",
          2550 => x"72",
          2551 => x"e8",
          2552 => x"bd",
          2553 => x"3f",
          2554 => x"ba",
          2555 => x"8d",
          2556 => x"c0",
          2557 => x"c4",
          2558 => x"3f",
          2559 => x"70",
          2560 => x"94",
          2561 => x"d3",
          2562 => x"d3",
          2563 => x"15",
          2564 => x"d3",
          2565 => x"f2",
          2566 => x"3f",
          2567 => x"51",
          2568 => x"80",
          2569 => x"80",
          2570 => x"3f",
          2571 => x"52",
          2572 => x"51",
          2573 => x"ec",
          2574 => x"04",
          2575 => x"77",
          2576 => x"56",
          2577 => x"53",
          2578 => x"81",
          2579 => x"33",
          2580 => x"06",
          2581 => x"a0",
          2582 => x"06",
          2583 => x"15",
          2584 => x"81",
          2585 => x"53",
          2586 => x"2e",
          2587 => x"81",
          2588 => x"73",
          2589 => x"82",
          2590 => x"72",
          2591 => x"e7",
          2592 => x"33",
          2593 => x"06",
          2594 => x"70",
          2595 => x"38",
          2596 => x"80",
          2597 => x"73",
          2598 => x"38",
          2599 => x"e1",
          2600 => x"81",
          2601 => x"54",
          2602 => x"09",
          2603 => x"38",
          2604 => x"a2",
          2605 => x"70",
          2606 => x"07",
          2607 => x"72",
          2608 => x"38",
          2609 => x"81",
          2610 => x"71",
          2611 => x"51",
          2612 => x"84",
          2613 => x"0d",
          2614 => x"2e",
          2615 => x"80",
          2616 => x"38",
          2617 => x"80",
          2618 => x"81",
          2619 => x"54",
          2620 => x"2e",
          2621 => x"54",
          2622 => x"15",
          2623 => x"53",
          2624 => x"2e",
          2625 => x"fe",
          2626 => x"39",
          2627 => x"76",
          2628 => x"8b",
          2629 => x"84",
          2630 => x"86",
          2631 => x"86",
          2632 => x"52",
          2633 => x"dc",
          2634 => x"84",
          2635 => x"e5",
          2636 => x"bb",
          2637 => x"3d",
          2638 => x"3d",
          2639 => x"11",
          2640 => x"52",
          2641 => x"70",
          2642 => x"98",
          2643 => x"33",
          2644 => x"82",
          2645 => x"26",
          2646 => x"84",
          2647 => x"83",
          2648 => x"26",
          2649 => x"85",
          2650 => x"84",
          2651 => x"26",
          2652 => x"86",
          2653 => x"85",
          2654 => x"26",
          2655 => x"88",
          2656 => x"86",
          2657 => x"e7",
          2658 => x"38",
          2659 => x"54",
          2660 => x"87",
          2661 => x"cc",
          2662 => x"87",
          2663 => x"0c",
          2664 => x"c0",
          2665 => x"82",
          2666 => x"c0",
          2667 => x"83",
          2668 => x"c0",
          2669 => x"84",
          2670 => x"c0",
          2671 => x"85",
          2672 => x"c0",
          2673 => x"86",
          2674 => x"c0",
          2675 => x"74",
          2676 => x"a4",
          2677 => x"c0",
          2678 => x"80",
          2679 => x"98",
          2680 => x"52",
          2681 => x"84",
          2682 => x"0d",
          2683 => x"0d",
          2684 => x"c0",
          2685 => x"81",
          2686 => x"c0",
          2687 => x"5e",
          2688 => x"87",
          2689 => x"08",
          2690 => x"1c",
          2691 => x"98",
          2692 => x"79",
          2693 => x"87",
          2694 => x"08",
          2695 => x"1c",
          2696 => x"98",
          2697 => x"79",
          2698 => x"87",
          2699 => x"08",
          2700 => x"1c",
          2701 => x"98",
          2702 => x"7b",
          2703 => x"87",
          2704 => x"08",
          2705 => x"1c",
          2706 => x"0c",
          2707 => x"ff",
          2708 => x"83",
          2709 => x"58",
          2710 => x"57",
          2711 => x"56",
          2712 => x"55",
          2713 => x"54",
          2714 => x"53",
          2715 => x"ff",
          2716 => x"d9",
          2717 => x"bf",
          2718 => x"3d",
          2719 => x"3d",
          2720 => x"05",
          2721 => x"81",
          2722 => x"72",
          2723 => x"de",
          2724 => x"84",
          2725 => x"70",
          2726 => x"52",
          2727 => x"09",
          2728 => x"38",
          2729 => x"e3",
          2730 => x"bb",
          2731 => x"3d",
          2732 => x"51",
          2733 => x"3f",
          2734 => x"08",
          2735 => x"98",
          2736 => x"71",
          2737 => x"81",
          2738 => x"72",
          2739 => x"9e",
          2740 => x"84",
          2741 => x"70",
          2742 => x"52",
          2743 => x"d2",
          2744 => x"fd",
          2745 => x"70",
          2746 => x"88",
          2747 => x"51",
          2748 => x"3f",
          2749 => x"08",
          2750 => x"98",
          2751 => x"71",
          2752 => x"38",
          2753 => x"81",
          2754 => x"83",
          2755 => x"38",
          2756 => x"84",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"33",
          2760 => x"33",
          2761 => x"06",
          2762 => x"70",
          2763 => x"f4",
          2764 => x"94",
          2765 => x"96",
          2766 => x"06",
          2767 => x"70",
          2768 => x"38",
          2769 => x"70",
          2770 => x"51",
          2771 => x"72",
          2772 => x"06",
          2773 => x"2e",
          2774 => x"93",
          2775 => x"52",
          2776 => x"73",
          2777 => x"51",
          2778 => x"80",
          2779 => x"2e",
          2780 => x"c0",
          2781 => x"74",
          2782 => x"84",
          2783 => x"86",
          2784 => x"71",
          2785 => x"81",
          2786 => x"70",
          2787 => x"81",
          2788 => x"53",
          2789 => x"cb",
          2790 => x"2a",
          2791 => x"71",
          2792 => x"38",
          2793 => x"84",
          2794 => x"2a",
          2795 => x"53",
          2796 => x"cf",
          2797 => x"ff",
          2798 => x"8f",
          2799 => x"30",
          2800 => x"51",
          2801 => x"83",
          2802 => x"83",
          2803 => x"fa",
          2804 => x"55",
          2805 => x"70",
          2806 => x"70",
          2807 => x"e7",
          2808 => x"83",
          2809 => x"70",
          2810 => x"54",
          2811 => x"80",
          2812 => x"38",
          2813 => x"94",
          2814 => x"2a",
          2815 => x"53",
          2816 => x"80",
          2817 => x"71",
          2818 => x"81",
          2819 => x"70",
          2820 => x"81",
          2821 => x"53",
          2822 => x"8a",
          2823 => x"2a",
          2824 => x"71",
          2825 => x"81",
          2826 => x"87",
          2827 => x"52",
          2828 => x"86",
          2829 => x"94",
          2830 => x"72",
          2831 => x"75",
          2832 => x"73",
          2833 => x"76",
          2834 => x"0c",
          2835 => x"04",
          2836 => x"70",
          2837 => x"51",
          2838 => x"72",
          2839 => x"06",
          2840 => x"2e",
          2841 => x"93",
          2842 => x"52",
          2843 => x"ff",
          2844 => x"c0",
          2845 => x"70",
          2846 => x"81",
          2847 => x"52",
          2848 => x"d7",
          2849 => x"0d",
          2850 => x"80",
          2851 => x"2a",
          2852 => x"52",
          2853 => x"84",
          2854 => x"c0",
          2855 => x"83",
          2856 => x"87",
          2857 => x"08",
          2858 => x"0c",
          2859 => x"94",
          2860 => x"c8",
          2861 => x"9e",
          2862 => x"f3",
          2863 => x"c0",
          2864 => x"83",
          2865 => x"87",
          2866 => x"08",
          2867 => x"0c",
          2868 => x"ac",
          2869 => x"d8",
          2870 => x"9e",
          2871 => x"f3",
          2872 => x"c0",
          2873 => x"83",
          2874 => x"87",
          2875 => x"08",
          2876 => x"0c",
          2877 => x"bc",
          2878 => x"e8",
          2879 => x"9e",
          2880 => x"f3",
          2881 => x"c0",
          2882 => x"83",
          2883 => x"87",
          2884 => x"08",
          2885 => x"f3",
          2886 => x"c0",
          2887 => x"83",
          2888 => x"87",
          2889 => x"08",
          2890 => x"0c",
          2891 => x"8c",
          2892 => x"80",
          2893 => x"83",
          2894 => x"80",
          2895 => x"9e",
          2896 => x"84",
          2897 => x"51",
          2898 => x"82",
          2899 => x"83",
          2900 => x"80",
          2901 => x"9e",
          2902 => x"88",
          2903 => x"51",
          2904 => x"80",
          2905 => x"81",
          2906 => x"f4",
          2907 => x"0b",
          2908 => x"90",
          2909 => x"80",
          2910 => x"52",
          2911 => x"2e",
          2912 => x"52",
          2913 => x"87",
          2914 => x"87",
          2915 => x"08",
          2916 => x"80",
          2917 => x"52",
          2918 => x"83",
          2919 => x"71",
          2920 => x"34",
          2921 => x"c0",
          2922 => x"70",
          2923 => x"06",
          2924 => x"70",
          2925 => x"38",
          2926 => x"83",
          2927 => x"80",
          2928 => x"9e",
          2929 => x"90",
          2930 => x"51",
          2931 => x"80",
          2932 => x"81",
          2933 => x"f4",
          2934 => x"0b",
          2935 => x"90",
          2936 => x"80",
          2937 => x"52",
          2938 => x"2e",
          2939 => x"52",
          2940 => x"8b",
          2941 => x"87",
          2942 => x"08",
          2943 => x"80",
          2944 => x"52",
          2945 => x"83",
          2946 => x"71",
          2947 => x"34",
          2948 => x"c0",
          2949 => x"70",
          2950 => x"06",
          2951 => x"70",
          2952 => x"38",
          2953 => x"83",
          2954 => x"80",
          2955 => x"9e",
          2956 => x"80",
          2957 => x"51",
          2958 => x"80",
          2959 => x"81",
          2960 => x"f4",
          2961 => x"0b",
          2962 => x"90",
          2963 => x"80",
          2964 => x"52",
          2965 => x"83",
          2966 => x"71",
          2967 => x"34",
          2968 => x"90",
          2969 => x"06",
          2970 => x"53",
          2971 => x"f4",
          2972 => x"0b",
          2973 => x"90",
          2974 => x"80",
          2975 => x"52",
          2976 => x"83",
          2977 => x"71",
          2978 => x"34",
          2979 => x"90",
          2980 => x"06",
          2981 => x"53",
          2982 => x"f4",
          2983 => x"0b",
          2984 => x"90",
          2985 => x"06",
          2986 => x"70",
          2987 => x"38",
          2988 => x"83",
          2989 => x"87",
          2990 => x"08",
          2991 => x"70",
          2992 => x"34",
          2993 => x"04",
          2994 => x"82",
          2995 => x"0d",
          2996 => x"51",
          2997 => x"3f",
          2998 => x"33",
          2999 => x"a0",
          3000 => x"a8",
          3001 => x"3f",
          3002 => x"33",
          3003 => x"f0",
          3004 => x"8b",
          3005 => x"85",
          3006 => x"f4",
          3007 => x"75",
          3008 => x"83",
          3009 => x"55",
          3010 => x"38",
          3011 => x"33",
          3012 => x"cc",
          3013 => x"8f",
          3014 => x"84",
          3015 => x"f4",
          3016 => x"73",
          3017 => x"83",
          3018 => x"55",
          3019 => x"38",
          3020 => x"33",
          3021 => x"c5",
          3022 => x"87",
          3023 => x"83",
          3024 => x"f4",
          3025 => x"74",
          3026 => x"83",
          3027 => x"56",
          3028 => x"38",
          3029 => x"33",
          3030 => x"e1",
          3031 => x"c0",
          3032 => x"3f",
          3033 => x"08",
          3034 => x"cc",
          3035 => x"9a",
          3036 => x"ec",
          3037 => x"da",
          3038 => x"b5",
          3039 => x"f3",
          3040 => x"83",
          3041 => x"ff",
          3042 => x"83",
          3043 => x"c1",
          3044 => x"f3",
          3045 => x"83",
          3046 => x"ff",
          3047 => x"83",
          3048 => x"56",
          3049 => x"52",
          3050 => x"fb",
          3051 => x"84",
          3052 => x"c0",
          3053 => x"31",
          3054 => x"bb",
          3055 => x"83",
          3056 => x"ff",
          3057 => x"83",
          3058 => x"55",
          3059 => x"83",
          3060 => x"55",
          3061 => x"87",
          3062 => x"83",
          3063 => x"56",
          3064 => x"52",
          3065 => x"bf",
          3066 => x"84",
          3067 => x"c0",
          3068 => x"31",
          3069 => x"bb",
          3070 => x"83",
          3071 => x"ff",
          3072 => x"87",
          3073 => x"83",
          3074 => x"56",
          3075 => x"52",
          3076 => x"93",
          3077 => x"84",
          3078 => x"c0",
          3079 => x"31",
          3080 => x"bb",
          3081 => x"83",
          3082 => x"ff",
          3083 => x"83",
          3084 => x"55",
          3085 => x"ff",
          3086 => x"9f",
          3087 => x"f8",
          3088 => x"3f",
          3089 => x"51",
          3090 => x"83",
          3091 => x"52",
          3092 => x"51",
          3093 => x"3f",
          3094 => x"08",
          3095 => x"f4",
          3096 => x"a6",
          3097 => x"f0",
          3098 => x"db",
          3099 => x"b3",
          3100 => x"db",
          3101 => x"bf",
          3102 => x"f3",
          3103 => x"83",
          3104 => x"ff",
          3105 => x"83",
          3106 => x"56",
          3107 => x"52",
          3108 => x"93",
          3109 => x"84",
          3110 => x"c0",
          3111 => x"31",
          3112 => x"bb",
          3113 => x"83",
          3114 => x"ff",
          3115 => x"83",
          3116 => x"55",
          3117 => x"fe",
          3118 => x"cb",
          3119 => x"80",
          3120 => x"b1",
          3121 => x"8e",
          3122 => x"80",
          3123 => x"38",
          3124 => x"83",
          3125 => x"ff",
          3126 => x"83",
          3127 => x"56",
          3128 => x"fc",
          3129 => x"39",
          3130 => x"51",
          3131 => x"3f",
          3132 => x"33",
          3133 => x"2e",
          3134 => x"d7",
          3135 => x"a0",
          3136 => x"f1",
          3137 => x"87",
          3138 => x"80",
          3139 => x"38",
          3140 => x"f4",
          3141 => x"83",
          3142 => x"ff",
          3143 => x"83",
          3144 => x"56",
          3145 => x"fc",
          3146 => x"39",
          3147 => x"33",
          3148 => x"d4",
          3149 => x"d2",
          3150 => x"91",
          3151 => x"80",
          3152 => x"38",
          3153 => x"f4",
          3154 => x"83",
          3155 => x"ff",
          3156 => x"83",
          3157 => x"54",
          3158 => x"fb",
          3159 => x"39",
          3160 => x"08",
          3161 => x"08",
          3162 => x"83",
          3163 => x"ff",
          3164 => x"83",
          3165 => x"56",
          3166 => x"fb",
          3167 => x"39",
          3168 => x"08",
          3169 => x"08",
          3170 => x"83",
          3171 => x"ff",
          3172 => x"83",
          3173 => x"54",
          3174 => x"fa",
          3175 => x"39",
          3176 => x"08",
          3177 => x"08",
          3178 => x"83",
          3179 => x"ff",
          3180 => x"83",
          3181 => x"55",
          3182 => x"fa",
          3183 => x"39",
          3184 => x"08",
          3185 => x"08",
          3186 => x"83",
          3187 => x"ff",
          3188 => x"83",
          3189 => x"56",
          3190 => x"fa",
          3191 => x"39",
          3192 => x"08",
          3193 => x"08",
          3194 => x"83",
          3195 => x"ff",
          3196 => x"83",
          3197 => x"54",
          3198 => x"f9",
          3199 => x"39",
          3200 => x"51",
          3201 => x"3f",
          3202 => x"51",
          3203 => x"3f",
          3204 => x"33",
          3205 => x"2e",
          3206 => x"c4",
          3207 => x"0d",
          3208 => x"33",
          3209 => x"26",
          3210 => x"10",
          3211 => x"8c",
          3212 => x"08",
          3213 => x"b4",
          3214 => x"ce",
          3215 => x"0d",
          3216 => x"bc",
          3217 => x"c2",
          3218 => x"0d",
          3219 => x"c4",
          3220 => x"b6",
          3221 => x"0d",
          3222 => x"cc",
          3223 => x"aa",
          3224 => x"0d",
          3225 => x"d4",
          3226 => x"9e",
          3227 => x"0d",
          3228 => x"dc",
          3229 => x"92",
          3230 => x"0d",
          3231 => x"80",
          3232 => x"0b",
          3233 => x"84",
          3234 => x"f4",
          3235 => x"c0",
          3236 => x"04",
          3237 => x"aa",
          3238 => x"3d",
          3239 => x"81",
          3240 => x"80",
          3241 => x"ec",
          3242 => x"87",
          3243 => x"bb",
          3244 => x"ed",
          3245 => x"57",
          3246 => x"f4",
          3247 => x"55",
          3248 => x"76",
          3249 => x"8e",
          3250 => x"84",
          3251 => x"a4",
          3252 => x"c0",
          3253 => x"bb",
          3254 => x"17",
          3255 => x"0b",
          3256 => x"08",
          3257 => x"84",
          3258 => x"ff",
          3259 => x"55",
          3260 => x"34",
          3261 => x"30",
          3262 => x"9f",
          3263 => x"55",
          3264 => x"85",
          3265 => x"b0",
          3266 => x"ec",
          3267 => x"08",
          3268 => x"87",
          3269 => x"bb",
          3270 => x"38",
          3271 => x"9a",
          3272 => x"bb",
          3273 => x"3d",
          3274 => x"e3",
          3275 => x"ad",
          3276 => x"76",
          3277 => x"06",
          3278 => x"52",
          3279 => x"89",
          3280 => x"ff",
          3281 => x"ab",
          3282 => x"84",
          3283 => x"76",
          3284 => x"83",
          3285 => x"ff",
          3286 => x"80",
          3287 => x"84",
          3288 => x"0d",
          3289 => x"0d",
          3290 => x"ad",
          3291 => x"72",
          3292 => x"57",
          3293 => x"73",
          3294 => x"92",
          3295 => x"8d",
          3296 => x"75",
          3297 => x"83",
          3298 => x"70",
          3299 => x"ff",
          3300 => x"84",
          3301 => x"53",
          3302 => x"08",
          3303 => x"f7",
          3304 => x"84",
          3305 => x"84",
          3306 => x"73",
          3307 => x"88",
          3308 => x"2e",
          3309 => x"16",
          3310 => x"06",
          3311 => x"76",
          3312 => x"80",
          3313 => x"bb",
          3314 => x"3d",
          3315 => x"1a",
          3316 => x"ff",
          3317 => x"ff",
          3318 => x"c7",
          3319 => x"bb",
          3320 => x"2e",
          3321 => x"1b",
          3322 => x"76",
          3323 => x"3f",
          3324 => x"08",
          3325 => x"54",
          3326 => x"c9",
          3327 => x"70",
          3328 => x"57",
          3329 => x"27",
          3330 => x"ff",
          3331 => x"33",
          3332 => x"76",
          3333 => x"e5",
          3334 => x"70",
          3335 => x"55",
          3336 => x"2e",
          3337 => x"fe",
          3338 => x"75",
          3339 => x"80",
          3340 => x"59",
          3341 => x"39",
          3342 => x"84",
          3343 => x"f4",
          3344 => x"56",
          3345 => x"3f",
          3346 => x"08",
          3347 => x"83",
          3348 => x"53",
          3349 => x"77",
          3350 => x"fa",
          3351 => x"84",
          3352 => x"ba",
          3353 => x"ff",
          3354 => x"84",
          3355 => x"55",
          3356 => x"bb",
          3357 => x"9d",
          3358 => x"84",
          3359 => x"70",
          3360 => x"80",
          3361 => x"53",
          3362 => x"16",
          3363 => x"52",
          3364 => x"f6",
          3365 => x"2e",
          3366 => x"ff",
          3367 => x"0b",
          3368 => x"0c",
          3369 => x"04",
          3370 => x"b6",
          3371 => x"3d",
          3372 => x"08",
          3373 => x"be",
          3374 => x"5b",
          3375 => x"80",
          3376 => x"34",
          3377 => x"33",
          3378 => x"f4",
          3379 => x"f4",
          3380 => x"74",
          3381 => x"76",
          3382 => x"56",
          3383 => x"2e",
          3384 => x"77",
          3385 => x"88",
          3386 => x"78",
          3387 => x"78",
          3388 => x"77",
          3389 => x"f8",
          3390 => x"b5",
          3391 => x"80",
          3392 => x"3f",
          3393 => x"08",
          3394 => x"98",
          3395 => x"79",
          3396 => x"d7",
          3397 => x"ff",
          3398 => x"c0",
          3399 => x"2b",
          3400 => x"84",
          3401 => x"70",
          3402 => x"97",
          3403 => x"2c",
          3404 => x"10",
          3405 => x"05",
          3406 => x"70",
          3407 => x"49",
          3408 => x"5b",
          3409 => x"81",
          3410 => x"2e",
          3411 => x"78",
          3412 => x"a8",
          3413 => x"80",
          3414 => x"ff",
          3415 => x"98",
          3416 => x"80",
          3417 => x"ec",
          3418 => x"16",
          3419 => x"56",
          3420 => x"83",
          3421 => x"33",
          3422 => x"62",
          3423 => x"83",
          3424 => x"08",
          3425 => x"56",
          3426 => x"2e",
          3427 => x"76",
          3428 => x"38",
          3429 => x"bc",
          3430 => x"76",
          3431 => x"ba",
          3432 => x"70",
          3433 => x"98",
          3434 => x"bc",
          3435 => x"2b",
          3436 => x"71",
          3437 => x"70",
          3438 => x"df",
          3439 => x"5f",
          3440 => x"58",
          3441 => x"7a",
          3442 => x"b1",
          3443 => x"e2",
          3444 => x"51",
          3445 => x"84",
          3446 => x"98",
          3447 => x"2c",
          3448 => x"ff",
          3449 => x"06",
          3450 => x"7d",
          3451 => x"8f",
          3452 => x"fe",
          3453 => x"57",
          3454 => x"38",
          3455 => x"0a",
          3456 => x"0a",
          3457 => x"2c",
          3458 => x"06",
          3459 => x"76",
          3460 => x"c0",
          3461 => x"16",
          3462 => x"51",
          3463 => x"83",
          3464 => x"33",
          3465 => x"62",
          3466 => x"83",
          3467 => x"08",
          3468 => x"43",
          3469 => x"2e",
          3470 => x"76",
          3471 => x"bc",
          3472 => x"39",
          3473 => x"80",
          3474 => x"38",
          3475 => x"81",
          3476 => x"39",
          3477 => x"fe",
          3478 => x"84",
          3479 => x"76",
          3480 => x"34",
          3481 => x"76",
          3482 => x"55",
          3483 => x"fd",
          3484 => x"10",
          3485 => x"a4",
          3486 => x"08",
          3487 => x"e8",
          3488 => x"0c",
          3489 => x"e2",
          3490 => x"0b",
          3491 => x"34",
          3492 => x"e2",
          3493 => x"75",
          3494 => x"e3",
          3495 => x"e8",
          3496 => x"51",
          3497 => x"3f",
          3498 => x"33",
          3499 => x"7a",
          3500 => x"34",
          3501 => x"84",
          3502 => x"70",
          3503 => x"84",
          3504 => x"5a",
          3505 => x"78",
          3506 => x"38",
          3507 => x"08",
          3508 => x"42",
          3509 => x"c8",
          3510 => x"70",
          3511 => x"ff",
          3512 => x"fc",
          3513 => x"93",
          3514 => x"38",
          3515 => x"90",
          3516 => x"10",
          3517 => x"05",
          3518 => x"58",
          3519 => x"38",
          3520 => x"e2",
          3521 => x"7c",
          3522 => x"c4",
          3523 => x"c8",
          3524 => x"74",
          3525 => x"38",
          3526 => x"08",
          3527 => x"ff",
          3528 => x"84",
          3529 => x"52",
          3530 => x"b4",
          3531 => x"e6",
          3532 => x"88",
          3533 => x"b8",
          3534 => x"c8",
          3535 => x"59",
          3536 => x"c8",
          3537 => x"ff",
          3538 => x"cc",
          3539 => x"ff",
          3540 => x"75",
          3541 => x"34",
          3542 => x"7c",
          3543 => x"f4",
          3544 => x"75",
          3545 => x"ff",
          3546 => x"ff",
          3547 => x"76",
          3548 => x"38",
          3549 => x"83",
          3550 => x"70",
          3551 => x"75",
          3552 => x"7c",
          3553 => x"f7",
          3554 => x"10",
          3555 => x"05",
          3556 => x"59",
          3557 => x"fa",
          3558 => x"51",
          3559 => x"3f",
          3560 => x"08",
          3561 => x"34",
          3562 => x"08",
          3563 => x"81",
          3564 => x"52",
          3565 => x"b7",
          3566 => x"e2",
          3567 => x"e2",
          3568 => x"56",
          3569 => x"ff",
          3570 => x"e6",
          3571 => x"88",
          3572 => x"9c",
          3573 => x"e8",
          3574 => x"51",
          3575 => x"3f",
          3576 => x"08",
          3577 => x"ff",
          3578 => x"84",
          3579 => x"ff",
          3580 => x"84",
          3581 => x"74",
          3582 => x"55",
          3583 => x"e2",
          3584 => x"81",
          3585 => x"e2",
          3586 => x"57",
          3587 => x"27",
          3588 => x"84",
          3589 => x"52",
          3590 => x"76",
          3591 => x"34",
          3592 => x"33",
          3593 => x"b2",
          3594 => x"e2",
          3595 => x"81",
          3596 => x"e2",
          3597 => x"57",
          3598 => x"27",
          3599 => x"84",
          3600 => x"52",
          3601 => x"76",
          3602 => x"34",
          3603 => x"33",
          3604 => x"b2",
          3605 => x"e2",
          3606 => x"81",
          3607 => x"e2",
          3608 => x"57",
          3609 => x"26",
          3610 => x"f9",
          3611 => x"e2",
          3612 => x"e2",
          3613 => x"56",
          3614 => x"f9",
          3615 => x"15",
          3616 => x"e2",
          3617 => x"98",
          3618 => x"2c",
          3619 => x"06",
          3620 => x"61",
          3621 => x"ef",
          3622 => x"e8",
          3623 => x"51",
          3624 => x"3f",
          3625 => x"33",
          3626 => x"70",
          3627 => x"e2",
          3628 => x"57",
          3629 => x"77",
          3630 => x"38",
          3631 => x"08",
          3632 => x"ff",
          3633 => x"74",
          3634 => x"29",
          3635 => x"05",
          3636 => x"84",
          3637 => x"5d",
          3638 => x"7b",
          3639 => x"38",
          3640 => x"08",
          3641 => x"ff",
          3642 => x"74",
          3643 => x"29",
          3644 => x"05",
          3645 => x"84",
          3646 => x"5d",
          3647 => x"75",
          3648 => x"38",
          3649 => x"7b",
          3650 => x"18",
          3651 => x"84",
          3652 => x"52",
          3653 => x"ff",
          3654 => x"75",
          3655 => x"29",
          3656 => x"05",
          3657 => x"84",
          3658 => x"5c",
          3659 => x"7a",
          3660 => x"38",
          3661 => x"81",
          3662 => x"34",
          3663 => x"08",
          3664 => x"51",
          3665 => x"3f",
          3666 => x"0a",
          3667 => x"0a",
          3668 => x"2c",
          3669 => x"33",
          3670 => x"79",
          3671 => x"a7",
          3672 => x"39",
          3673 => x"33",
          3674 => x"2e",
          3675 => x"84",
          3676 => x"52",
          3677 => x"af",
          3678 => x"e2",
          3679 => x"05",
          3680 => x"e2",
          3681 => x"81",
          3682 => x"dd",
          3683 => x"c4",
          3684 => x"41",
          3685 => x"84",
          3686 => x"52",
          3687 => x"af",
          3688 => x"e2",
          3689 => x"51",
          3690 => x"84",
          3691 => x"81",
          3692 => x"77",
          3693 => x"84",
          3694 => x"57",
          3695 => x"80",
          3696 => x"f4",
          3697 => x"10",
          3698 => x"9c",
          3699 => x"57",
          3700 => x"8b",
          3701 => x"82",
          3702 => x"06",
          3703 => x"05",
          3704 => x"53",
          3705 => x"e8",
          3706 => x"bb",
          3707 => x"0c",
          3708 => x"33",
          3709 => x"83",
          3710 => x"70",
          3711 => x"83",
          3712 => x"5b",
          3713 => x"3f",
          3714 => x"33",
          3715 => x"83",
          3716 => x"70",
          3717 => x"5e",
          3718 => x"38",
          3719 => x"08",
          3720 => x"2e",
          3721 => x"f4",
          3722 => x"77",
          3723 => x"de",
          3724 => x"84",
          3725 => x"80",
          3726 => x"c4",
          3727 => x"bb",
          3728 => x"3d",
          3729 => x"e2",
          3730 => x"74",
          3731 => x"38",
          3732 => x"08",
          3733 => x"ff",
          3734 => x"84",
          3735 => x"52",
          3736 => x"ae",
          3737 => x"e6",
          3738 => x"88",
          3739 => x"80",
          3740 => x"c8",
          3741 => x"42",
          3742 => x"c8",
          3743 => x"ff",
          3744 => x"cc",
          3745 => x"80",
          3746 => x"fe",
          3747 => x"84",
          3748 => x"80",
          3749 => x"c4",
          3750 => x"39",
          3751 => x"33",
          3752 => x"06",
          3753 => x"80",
          3754 => x"38",
          3755 => x"33",
          3756 => x"79",
          3757 => x"34",
          3758 => x"77",
          3759 => x"34",
          3760 => x"08",
          3761 => x"ff",
          3762 => x"84",
          3763 => x"70",
          3764 => x"98",
          3765 => x"c4",
          3766 => x"5a",
          3767 => x"24",
          3768 => x"84",
          3769 => x"52",
          3770 => x"ad",
          3771 => x"e2",
          3772 => x"98",
          3773 => x"2c",
          3774 => x"33",
          3775 => x"56",
          3776 => x"f3",
          3777 => x"e6",
          3778 => x"88",
          3779 => x"e0",
          3780 => x"80",
          3781 => x"80",
          3782 => x"98",
          3783 => x"c4",
          3784 => x"55",
          3785 => x"f3",
          3786 => x"e6",
          3787 => x"88",
          3788 => x"bc",
          3789 => x"80",
          3790 => x"80",
          3791 => x"98",
          3792 => x"c4",
          3793 => x"55",
          3794 => x"ff",
          3795 => x"af",
          3796 => x"57",
          3797 => x"77",
          3798 => x"e8",
          3799 => x"33",
          3800 => x"8c",
          3801 => x"80",
          3802 => x"80",
          3803 => x"98",
          3804 => x"c4",
          3805 => x"5b",
          3806 => x"fe",
          3807 => x"16",
          3808 => x"33",
          3809 => x"e6",
          3810 => x"76",
          3811 => x"ab",
          3812 => x"81",
          3813 => x"81",
          3814 => x"70",
          3815 => x"e2",
          3816 => x"57",
          3817 => x"24",
          3818 => x"fe",
          3819 => x"7c",
          3820 => x"81",
          3821 => x"e2",
          3822 => x"74",
          3823 => x"38",
          3824 => x"08",
          3825 => x"ff",
          3826 => x"84",
          3827 => x"52",
          3828 => x"ab",
          3829 => x"e6",
          3830 => x"88",
          3831 => x"90",
          3832 => x"c8",
          3833 => x"5d",
          3834 => x"c8",
          3835 => x"ff",
          3836 => x"cc",
          3837 => x"80",
          3838 => x"8e",
          3839 => x"84",
          3840 => x"80",
          3841 => x"c4",
          3842 => x"bb",
          3843 => x"3d",
          3844 => x"e2",
          3845 => x"81",
          3846 => x"58",
          3847 => x"f1",
          3848 => x"e2",
          3849 => x"76",
          3850 => x"38",
          3851 => x"70",
          3852 => x"42",
          3853 => x"a1",
          3854 => x"5b",
          3855 => x"1c",
          3856 => x"80",
          3857 => x"ff",
          3858 => x"98",
          3859 => x"c8",
          3860 => x"58",
          3861 => x"e1",
          3862 => x"55",
          3863 => x"c8",
          3864 => x"ff",
          3865 => x"59",
          3866 => x"79",
          3867 => x"c4",
          3868 => x"61",
          3869 => x"81",
          3870 => x"84",
          3871 => x"75",
          3872 => x"c8",
          3873 => x"80",
          3874 => x"ff",
          3875 => x"98",
          3876 => x"ff",
          3877 => x"5c",
          3878 => x"24",
          3879 => x"77",
          3880 => x"98",
          3881 => x"ff",
          3882 => x"5a",
          3883 => x"f0",
          3884 => x"e6",
          3885 => x"88",
          3886 => x"b4",
          3887 => x"80",
          3888 => x"80",
          3889 => x"98",
          3890 => x"c4",
          3891 => x"42",
          3892 => x"f0",
          3893 => x"e6",
          3894 => x"88",
          3895 => x"90",
          3896 => x"80",
          3897 => x"80",
          3898 => x"98",
          3899 => x"c4",
          3900 => x"42",
          3901 => x"ff",
          3902 => x"83",
          3903 => x"51",
          3904 => x"3f",
          3905 => x"08",
          3906 => x"0c",
          3907 => x"08",
          3908 => x"c0",
          3909 => x"f2",
          3910 => x"ec",
          3911 => x"86",
          3912 => x"83",
          3913 => x"77",
          3914 => x"80",
          3915 => x"e6",
          3916 => x"7b",
          3917 => x"52",
          3918 => x"b4",
          3919 => x"80",
          3920 => x"80",
          3921 => x"98",
          3922 => x"c4",
          3923 => x"57",
          3924 => x"da",
          3925 => x"c8",
          3926 => x"2b",
          3927 => x"79",
          3928 => x"5c",
          3929 => x"75",
          3930 => x"93",
          3931 => x"39",
          3932 => x"08",
          3933 => x"81",
          3934 => x"9c",
          3935 => x"76",
          3936 => x"bb",
          3937 => x"84",
          3938 => x"75",
          3939 => x"38",
          3940 => x"f4",
          3941 => x"f4",
          3942 => x"74",
          3943 => x"d9",
          3944 => x"81",
          3945 => x"83",
          3946 => x"51",
          3947 => x"3f",
          3948 => x"f4",
          3949 => x"3d",
          3950 => x"40",
          3951 => x"74",
          3952 => x"97",
          3953 => x"0c",
          3954 => x"18",
          3955 => x"80",
          3956 => x"38",
          3957 => x"75",
          3958 => x"ce",
          3959 => x"84",
          3960 => x"c4",
          3961 => x"84",
          3962 => x"06",
          3963 => x"75",
          3964 => x"ff",
          3965 => x"93",
          3966 => x"c4",
          3967 => x"c8",
          3968 => x"5d",
          3969 => x"f2",
          3970 => x"e6",
          3971 => x"88",
          3972 => x"dc",
          3973 => x"e8",
          3974 => x"51",
          3975 => x"3f",
          3976 => x"08",
          3977 => x"ff",
          3978 => x"84",
          3979 => x"ff",
          3980 => x"84",
          3981 => x"78",
          3982 => x"55",
          3983 => x"51",
          3984 => x"3f",
          3985 => x"08",
          3986 => x"34",
          3987 => x"08",
          3988 => x"81",
          3989 => x"52",
          3990 => x"aa",
          3991 => x"84",
          3992 => x"84",
          3993 => x"57",
          3994 => x"80",
          3995 => x"38",
          3996 => x"08",
          3997 => x"ff",
          3998 => x"84",
          3999 => x"52",
          4000 => x"a5",
          4001 => x"e6",
          4002 => x"88",
          4003 => x"e0",
          4004 => x"c8",
          4005 => x"57",
          4006 => x"c8",
          4007 => x"ff",
          4008 => x"39",
          4009 => x"a9",
          4010 => x"bb",
          4011 => x"e2",
          4012 => x"bb",
          4013 => x"ff",
          4014 => x"53",
          4015 => x"51",
          4016 => x"3f",
          4017 => x"81",
          4018 => x"e2",
          4019 => x"e2",
          4020 => x"52",
          4021 => x"80",
          4022 => x"38",
          4023 => x"08",
          4024 => x"ff",
          4025 => x"84",
          4026 => x"52",
          4027 => x"a4",
          4028 => x"e6",
          4029 => x"88",
          4030 => x"f4",
          4031 => x"c8",
          4032 => x"5b",
          4033 => x"c8",
          4034 => x"ff",
          4035 => x"39",
          4036 => x"80",
          4037 => x"c8",
          4038 => x"84",
          4039 => x"7b",
          4040 => x"0c",
          4041 => x"04",
          4042 => x"08",
          4043 => x"2e",
          4044 => x"75",
          4045 => x"f2",
          4046 => x"84",
          4047 => x"c4",
          4048 => x"84",
          4049 => x"06",
          4050 => x"75",
          4051 => x"ff",
          4052 => x"84",
          4053 => x"84",
          4054 => x"56",
          4055 => x"2e",
          4056 => x"84",
          4057 => x"52",
          4058 => x"a4",
          4059 => x"e6",
          4060 => x"a0",
          4061 => x"f8",
          4062 => x"e8",
          4063 => x"51",
          4064 => x"3f",
          4065 => x"33",
          4066 => x"78",
          4067 => x"34",
          4068 => x"06",
          4069 => x"74",
          4070 => x"bf",
          4071 => x"f4",
          4072 => x"2b",
          4073 => x"83",
          4074 => x"81",
          4075 => x"52",
          4076 => x"dd",
          4077 => x"bb",
          4078 => x"0c",
          4079 => x"33",
          4080 => x"83",
          4081 => x"70",
          4082 => x"83",
          4083 => x"5b",
          4084 => x"3f",
          4085 => x"33",
          4086 => x"83",
          4087 => x"70",
          4088 => x"5e",
          4089 => x"f4",
          4090 => x"53",
          4091 => x"51",
          4092 => x"3f",
          4093 => x"33",
          4094 => x"81",
          4095 => x"56",
          4096 => x"83",
          4097 => x"83",
          4098 => x"f4",
          4099 => x"3d",
          4100 => x"54",
          4101 => x"52",
          4102 => x"d9",
          4103 => x"f4",
          4104 => x"8a",
          4105 => x"fc",
          4106 => x"ec",
          4107 => x"de",
          4108 => x"0b",
          4109 => x"34",
          4110 => x"e2",
          4111 => x"84",
          4112 => x"b5",
          4113 => x"93",
          4114 => x"74",
          4115 => x"a8",
          4116 => x"84",
          4117 => x"38",
          4118 => x"08",
          4119 => x"5d",
          4120 => x"08",
          4121 => x"52",
          4122 => x"b7",
          4123 => x"bb",
          4124 => x"84",
          4125 => x"7b",
          4126 => x"06",
          4127 => x"84",
          4128 => x"51",
          4129 => x"3f",
          4130 => x"08",
          4131 => x"84",
          4132 => x"25",
          4133 => x"84",
          4134 => x"ff",
          4135 => x"57",
          4136 => x"34",
          4137 => x"06",
          4138 => x"33",
          4139 => x"83",
          4140 => x"70",
          4141 => x"57",
          4142 => x"8a",
          4143 => x"2b",
          4144 => x"83",
          4145 => x"81",
          4146 => x"57",
          4147 => x"fb",
          4148 => x"84",
          4149 => x"83",
          4150 => x"70",
          4151 => x"f4",
          4152 => x"08",
          4153 => x"e3",
          4154 => x"ff",
          4155 => x"83",
          4156 => x"70",
          4157 => x"f4",
          4158 => x"08",
          4159 => x"74",
          4160 => x"1d",
          4161 => x"06",
          4162 => x"7d",
          4163 => x"80",
          4164 => x"2e",
          4165 => x"fe",
          4166 => x"e7",
          4167 => x"d0",
          4168 => x"79",
          4169 => x"ff",
          4170 => x"83",
          4171 => x"81",
          4172 => x"ff",
          4173 => x"93",
          4174 => x"e0",
          4175 => x"83",
          4176 => x"ff",
          4177 => x"51",
          4178 => x"3f",
          4179 => x"33",
          4180 => x"87",
          4181 => x"f4",
          4182 => x"1b",
          4183 => x"40",
          4184 => x"e7",
          4185 => x"84",
          4186 => x"83",
          4187 => x"70",
          4188 => x"f4",
          4189 => x"08",
          4190 => x"e3",
          4191 => x"ff",
          4192 => x"83",
          4193 => x"70",
          4194 => x"f4",
          4195 => x"08",
          4196 => x"74",
          4197 => x"ea",
          4198 => x"39",
          4199 => x"f4",
          4200 => x"39",
          4201 => x"f4",
          4202 => x"39",
          4203 => x"51",
          4204 => x"3f",
          4205 => x"38",
          4206 => x"f2",
          4207 => x"80",
          4208 => x"02",
          4209 => x"c7",
          4210 => x"53",
          4211 => x"81",
          4212 => x"81",
          4213 => x"38",
          4214 => x"83",
          4215 => x"82",
          4216 => x"38",
          4217 => x"80",
          4218 => x"b0",
          4219 => x"57",
          4220 => x"a0",
          4221 => x"2e",
          4222 => x"83",
          4223 => x"75",
          4224 => x"34",
          4225 => x"b2",
          4226 => x"b0",
          4227 => x"2b",
          4228 => x"07",
          4229 => x"07",
          4230 => x"7f",
          4231 => x"5b",
          4232 => x"94",
          4233 => x"70",
          4234 => x"0c",
          4235 => x"84",
          4236 => x"76",
          4237 => x"38",
          4238 => x"a2",
          4239 => x"b0",
          4240 => x"d6",
          4241 => x"31",
          4242 => x"a0",
          4243 => x"15",
          4244 => x"70",
          4245 => x"34",
          4246 => x"72",
          4247 => x"3d",
          4248 => x"c7",
          4249 => x"83",
          4250 => x"70",
          4251 => x"83",
          4252 => x"71",
          4253 => x"74",
          4254 => x"58",
          4255 => x"c7",
          4256 => x"84",
          4257 => x"70",
          4258 => x"84",
          4259 => x"70",
          4260 => x"83",
          4261 => x"70",
          4262 => x"06",
          4263 => x"5d",
          4264 => x"5e",
          4265 => x"73",
          4266 => x"38",
          4267 => x"75",
          4268 => x"81",
          4269 => x"81",
          4270 => x"81",
          4271 => x"83",
          4272 => x"62",
          4273 => x"70",
          4274 => x"5d",
          4275 => x"5b",
          4276 => x"26",
          4277 => x"fa",
          4278 => x"76",
          4279 => x"7d",
          4280 => x"5f",
          4281 => x"5c",
          4282 => x"fe",
          4283 => x"7d",
          4284 => x"77",
          4285 => x"38",
          4286 => x"81",
          4287 => x"83",
          4288 => x"74",
          4289 => x"56",
          4290 => x"86",
          4291 => x"59",
          4292 => x"80",
          4293 => x"f8",
          4294 => x"ff",
          4295 => x"f7",
          4296 => x"ff",
          4297 => x"b2",
          4298 => x"29",
          4299 => x"57",
          4300 => x"57",
          4301 => x"81",
          4302 => x"81",
          4303 => x"81",
          4304 => x"71",
          4305 => x"54",
          4306 => x"2e",
          4307 => x"80",
          4308 => x"b4",
          4309 => x"83",
          4310 => x"83",
          4311 => x"70",
          4312 => x"90",
          4313 => x"88",
          4314 => x"07",
          4315 => x"56",
          4316 => x"79",
          4317 => x"38",
          4318 => x"72",
          4319 => x"83",
          4320 => x"70",
          4321 => x"70",
          4322 => x"83",
          4323 => x"71",
          4324 => x"86",
          4325 => x"11",
          4326 => x"56",
          4327 => x"c7",
          4328 => x"14",
          4329 => x"33",
          4330 => x"06",
          4331 => x"33",
          4332 => x"06",
          4333 => x"22",
          4334 => x"ff",
          4335 => x"29",
          4336 => x"5a",
          4337 => x"5f",
          4338 => x"79",
          4339 => x"38",
          4340 => x"15",
          4341 => x"19",
          4342 => x"81",
          4343 => x"81",
          4344 => x"71",
          4345 => x"ff",
          4346 => x"81",
          4347 => x"75",
          4348 => x"5b",
          4349 => x"7b",
          4350 => x"38",
          4351 => x"53",
          4352 => x"16",
          4353 => x"5b",
          4354 => x"e2",
          4355 => x"06",
          4356 => x"da",
          4357 => x"39",
          4358 => x"7b",
          4359 => x"9a",
          4360 => x"0d",
          4361 => x"8c",
          4362 => x"73",
          4363 => x"34",
          4364 => x"81",
          4365 => x"8e",
          4366 => x"80",
          4367 => x"ff",
          4368 => x"87",
          4369 => x"56",
          4370 => x"80",
          4371 => x"8e",
          4372 => x"8a",
          4373 => x"74",
          4374 => x"75",
          4375 => x"83",
          4376 => x"3f",
          4377 => x"e0",
          4378 => x"54",
          4379 => x"86",
          4380 => x"73",
          4381 => x"07",
          4382 => x"75",
          4383 => x"70",
          4384 => x"80",
          4385 => x"53",
          4386 => x"86",
          4387 => x"08",
          4388 => x"81",
          4389 => x"72",
          4390 => x"f3",
          4391 => x"81",
          4392 => x"07",
          4393 => x"34",
          4394 => x"84",
          4395 => x"80",
          4396 => x"84",
          4397 => x"0d",
          4398 => x"f8",
          4399 => x"84",
          4400 => x"3d",
          4401 => x"05",
          4402 => x"05",
          4403 => x"84",
          4404 => x"5b",
          4405 => x"53",
          4406 => x"82",
          4407 => x"b8",
          4408 => x"fa",
          4409 => x"fa",
          4410 => x"71",
          4411 => x"c7",
          4412 => x"83",
          4413 => x"5f",
          4414 => x"71",
          4415 => x"70",
          4416 => x"06",
          4417 => x"33",
          4418 => x"53",
          4419 => x"83",
          4420 => x"fa",
          4421 => x"05",
          4422 => x"fa",
          4423 => x"fa",
          4424 => x"05",
          4425 => x"06",
          4426 => x"06",
          4427 => x"72",
          4428 => x"8c",
          4429 => x"53",
          4430 => x"b4",
          4431 => x"b2",
          4432 => x"ff",
          4433 => x"b8",
          4434 => x"55",
          4435 => x"26",
          4436 => x"84",
          4437 => x"76",
          4438 => x"58",
          4439 => x"9f",
          4440 => x"38",
          4441 => x"70",
          4442 => x"e0",
          4443 => x"e0",
          4444 => x"72",
          4445 => x"54",
          4446 => x"81",
          4447 => x"81",
          4448 => x"b8",
          4449 => x"e3",
          4450 => x"9f",
          4451 => x"83",
          4452 => x"84",
          4453 => x"54",
          4454 => x"e0",
          4455 => x"74",
          4456 => x"05",
          4457 => x"14",
          4458 => x"74",
          4459 => x"84",
          4460 => x"ff",
          4461 => x"83",
          4462 => x"75",
          4463 => x"ff",
          4464 => x"ff",
          4465 => x"54",
          4466 => x"81",
          4467 => x"74",
          4468 => x"84",
          4469 => x"71",
          4470 => x"55",
          4471 => x"86",
          4472 => x"58",
          4473 => x"80",
          4474 => x"06",
          4475 => x"06",
          4476 => x"19",
          4477 => x"57",
          4478 => x"b9",
          4479 => x"d6",
          4480 => x"e0",
          4481 => x"84",
          4482 => x"33",
          4483 => x"05",
          4484 => x"70",
          4485 => x"33",
          4486 => x"05",
          4487 => x"15",
          4488 => x"33",
          4489 => x"33",
          4490 => x"19",
          4491 => x"55",
          4492 => x"ce",
          4493 => x"72",
          4494 => x"0c",
          4495 => x"04",
          4496 => x"b4",
          4497 => x"b2",
          4498 => x"ff",
          4499 => x"b8",
          4500 => x"55",
          4501 => x"27",
          4502 => x"77",
          4503 => x"dd",
          4504 => x"ff",
          4505 => x"83",
          4506 => x"56",
          4507 => x"2e",
          4508 => x"fe",
          4509 => x"76",
          4510 => x"84",
          4511 => x"71",
          4512 => x"72",
          4513 => x"52",
          4514 => x"73",
          4515 => x"38",
          4516 => x"33",
          4517 => x"15",
          4518 => x"55",
          4519 => x"0b",
          4520 => x"34",
          4521 => x"81",
          4522 => x"ff",
          4523 => x"80",
          4524 => x"38",
          4525 => x"e0",
          4526 => x"75",
          4527 => x"57",
          4528 => x"53",
          4529 => x"fd",
          4530 => x"0b",
          4531 => x"33",
          4532 => x"89",
          4533 => x"b6",
          4534 => x"84",
          4535 => x"33",
          4536 => x"b8",
          4537 => x"fc",
          4538 => x"3d",
          4539 => x"84",
          4540 => x"33",
          4541 => x"86",
          4542 => x"70",
          4543 => x"c4",
          4544 => x"70",
          4545 => x"b8",
          4546 => x"71",
          4547 => x"38",
          4548 => x"b5",
          4549 => x"84",
          4550 => x"86",
          4551 => x"80",
          4552 => x"b5",
          4553 => x"b4",
          4554 => x"ff",
          4555 => x"72",
          4556 => x"38",
          4557 => x"70",
          4558 => x"34",
          4559 => x"bb",
          4560 => x"3d",
          4561 => x"fa",
          4562 => x"73",
          4563 => x"70",
          4564 => x"06",
          4565 => x"54",
          4566 => x"b4",
          4567 => x"83",
          4568 => x"72",
          4569 => x"f7",
          4570 => x"55",
          4571 => x"75",
          4572 => x"70",
          4573 => x"fa",
          4574 => x"0b",
          4575 => x"0c",
          4576 => x"04",
          4577 => x"33",
          4578 => x"70",
          4579 => x"2c",
          4580 => x"56",
          4581 => x"83",
          4582 => x"80",
          4583 => x"84",
          4584 => x"0d",
          4585 => x"b5",
          4586 => x"84",
          4587 => x"ff",
          4588 => x"51",
          4589 => x"83",
          4590 => x"72",
          4591 => x"34",
          4592 => x"bb",
          4593 => x"3d",
          4594 => x"0b",
          4595 => x"34",
          4596 => x"33",
          4597 => x"33",
          4598 => x"52",
          4599 => x"fe",
          4600 => x"12",
          4601 => x"fa",
          4602 => x"d0",
          4603 => x"0d",
          4604 => x"33",
          4605 => x"26",
          4606 => x"10",
          4607 => x"98",
          4608 => x"08",
          4609 => x"b0",
          4610 => x"f0",
          4611 => x"2b",
          4612 => x"70",
          4613 => x"07",
          4614 => x"51",
          4615 => x"2e",
          4616 => x"9c",
          4617 => x"0b",
          4618 => x"34",
          4619 => x"bb",
          4620 => x"3d",
          4621 => x"fa",
          4622 => x"9f",
          4623 => x"51",
          4624 => x"b0",
          4625 => x"84",
          4626 => x"83",
          4627 => x"83",
          4628 => x"80",
          4629 => x"70",
          4630 => x"34",
          4631 => x"fa",
          4632 => x"fe",
          4633 => x"51",
          4634 => x"b0",
          4635 => x"80",
          4636 => x"fa",
          4637 => x"0b",
          4638 => x"0c",
          4639 => x"04",
          4640 => x"33",
          4641 => x"84",
          4642 => x"83",
          4643 => x"ff",
          4644 => x"fa",
          4645 => x"07",
          4646 => x"fa",
          4647 => x"a5",
          4648 => x"b0",
          4649 => x"06",
          4650 => x"70",
          4651 => x"34",
          4652 => x"83",
          4653 => x"81",
          4654 => x"07",
          4655 => x"fa",
          4656 => x"81",
          4657 => x"b0",
          4658 => x"06",
          4659 => x"70",
          4660 => x"34",
          4661 => x"83",
          4662 => x"81",
          4663 => x"70",
          4664 => x"34",
          4665 => x"83",
          4666 => x"81",
          4667 => x"d0",
          4668 => x"83",
          4669 => x"fe",
          4670 => x"fa",
          4671 => x"bf",
          4672 => x"51",
          4673 => x"b0",
          4674 => x"39",
          4675 => x"33",
          4676 => x"80",
          4677 => x"70",
          4678 => x"34",
          4679 => x"83",
          4680 => x"81",
          4681 => x"c0",
          4682 => x"83",
          4683 => x"fe",
          4684 => x"fa",
          4685 => x"af",
          4686 => x"51",
          4687 => x"b0",
          4688 => x"39",
          4689 => x"33",
          4690 => x"51",
          4691 => x"b0",
          4692 => x"39",
          4693 => x"33",
          4694 => x"82",
          4695 => x"83",
          4696 => x"fd",
          4697 => x"3d",
          4698 => x"05",
          4699 => x"05",
          4700 => x"33",
          4701 => x"33",
          4702 => x"33",
          4703 => x"33",
          4704 => x"33",
          4705 => x"5d",
          4706 => x"82",
          4707 => x"38",
          4708 => x"a5",
          4709 => x"2e",
          4710 => x"7d",
          4711 => x"34",
          4712 => x"b8",
          4713 => x"83",
          4714 => x"7b",
          4715 => x"23",
          4716 => x"b5",
          4717 => x"0d",
          4718 => x"2e",
          4719 => x"db",
          4720 => x"84",
          4721 => x"81",
          4722 => x"fc",
          4723 => x"83",
          4724 => x"a8",
          4725 => x"b5",
          4726 => x"83",
          4727 => x"79",
          4728 => x"f8",
          4729 => x"b8",
          4730 => x"84",
          4731 => x"55",
          4732 => x"53",
          4733 => x"e4",
          4734 => x"80",
          4735 => x"84",
          4736 => x"80",
          4737 => x"fc",
          4738 => x"fa",
          4739 => x"83",
          4740 => x"7c",
          4741 => x"34",
          4742 => x"04",
          4743 => x"b8",
          4744 => x"0b",
          4745 => x"34",
          4746 => x"fa",
          4747 => x"0b",
          4748 => x"34",
          4749 => x"fa",
          4750 => x"ba",
          4751 => x"84",
          4752 => x"57",
          4753 => x"33",
          4754 => x"7b",
          4755 => x"7a",
          4756 => x"94",
          4757 => x"b2",
          4758 => x"84",
          4759 => x"5a",
          4760 => x"27",
          4761 => x"10",
          4762 => x"05",
          4763 => x"59",
          4764 => x"51",
          4765 => x"3f",
          4766 => x"81",
          4767 => x"ba",
          4768 => x"5b",
          4769 => x"26",
          4770 => x"d3",
          4771 => x"fe",
          4772 => x"84",
          4773 => x"80",
          4774 => x"fc",
          4775 => x"fa",
          4776 => x"83",
          4777 => x"7c",
          4778 => x"34",
          4779 => x"04",
          4780 => x"b8",
          4781 => x"0b",
          4782 => x"34",
          4783 => x"fa",
          4784 => x"0b",
          4785 => x"34",
          4786 => x"fa",
          4787 => x"f8",
          4788 => x"90",
          4789 => x"bb",
          4790 => x"83",
          4791 => x"fe",
          4792 => x"80",
          4793 => x"e8",
          4794 => x"be",
          4795 => x"bb",
          4796 => x"fd",
          4797 => x"f8",
          4798 => x"52",
          4799 => x"51",
          4800 => x"3f",
          4801 => x"81",
          4802 => x"5a",
          4803 => x"3d",
          4804 => x"84",
          4805 => x"33",
          4806 => x"33",
          4807 => x"33",
          4808 => x"33",
          4809 => x"12",
          4810 => x"80",
          4811 => x"b2",
          4812 => x"59",
          4813 => x"29",
          4814 => x"ff",
          4815 => x"f9",
          4816 => x"59",
          4817 => x"57",
          4818 => x"81",
          4819 => x"89",
          4820 => x"38",
          4821 => x"81",
          4822 => x"81",
          4823 => x"38",
          4824 => x"82",
          4825 => x"b8",
          4826 => x"fa",
          4827 => x"fa",
          4828 => x"72",
          4829 => x"56",
          4830 => x"80",
          4831 => x"c7",
          4832 => x"34",
          4833 => x"33",
          4834 => x"33",
          4835 => x"22",
          4836 => x"12",
          4837 => x"53",
          4838 => x"b6",
          4839 => x"fa",
          4840 => x"71",
          4841 => x"54",
          4842 => x"33",
          4843 => x"80",
          4844 => x"b8",
          4845 => x"81",
          4846 => x"fa",
          4847 => x"fa",
          4848 => x"72",
          4849 => x"5b",
          4850 => x"83",
          4851 => x"84",
          4852 => x"34",
          4853 => x"81",
          4854 => x"55",
          4855 => x"81",
          4856 => x"b8",
          4857 => x"77",
          4858 => x"ff",
          4859 => x"83",
          4860 => x"84",
          4861 => x"53",
          4862 => x"8c",
          4863 => x"fc",
          4864 => x"80",
          4865 => x"38",
          4866 => x"bb",
          4867 => x"3d",
          4868 => x"8d",
          4869 => x"75",
          4870 => x"f7",
          4871 => x"2e",
          4872 => x"fe",
          4873 => x"52",
          4874 => x"96",
          4875 => x"83",
          4876 => x"ff",
          4877 => x"fa",
          4878 => x"53",
          4879 => x"13",
          4880 => x"75",
          4881 => x"81",
          4882 => x"38",
          4883 => x"52",
          4884 => x"ba",
          4885 => x"70",
          4886 => x"54",
          4887 => x"26",
          4888 => x"76",
          4889 => x"fd",
          4890 => x"13",
          4891 => x"06",
          4892 => x"73",
          4893 => x"fe",
          4894 => x"83",
          4895 => x"fe",
          4896 => x"52",
          4897 => x"de",
          4898 => x"84",
          4899 => x"89",
          4900 => x"75",
          4901 => x"09",
          4902 => x"ca",
          4903 => x"b5",
          4904 => x"ff",
          4905 => x"05",
          4906 => x"38",
          4907 => x"83",
          4908 => x"76",
          4909 => x"fc",
          4910 => x"fa",
          4911 => x"81",
          4912 => x"ff",
          4913 => x"fe",
          4914 => x"53",
          4915 => x"b5",
          4916 => x"39",
          4917 => x"fa",
          4918 => x"52",
          4919 => x"e2",
          4920 => x"39",
          4921 => x"51",
          4922 => x"fe",
          4923 => x"3d",
          4924 => x"f3",
          4925 => x"ba",
          4926 => x"59",
          4927 => x"81",
          4928 => x"82",
          4929 => x"38",
          4930 => x"84",
          4931 => x"8a",
          4932 => x"38",
          4933 => x"84",
          4934 => x"89",
          4935 => x"38",
          4936 => x"33",
          4937 => x"33",
          4938 => x"33",
          4939 => x"05",
          4940 => x"84",
          4941 => x"33",
          4942 => x"80",
          4943 => x"b8",
          4944 => x"fa",
          4945 => x"fa",
          4946 => x"71",
          4947 => x"5a",
          4948 => x"83",
          4949 => x"34",
          4950 => x"33",
          4951 => x"62",
          4952 => x"83",
          4953 => x"7f",
          4954 => x"80",
          4955 => x"b8",
          4956 => x"81",
          4957 => x"fa",
          4958 => x"fa",
          4959 => x"72",
          4960 => x"40",
          4961 => x"83",
          4962 => x"84",
          4963 => x"34",
          4964 => x"81",
          4965 => x"58",
          4966 => x"81",
          4967 => x"b8",
          4968 => x"79",
          4969 => x"ff",
          4970 => x"83",
          4971 => x"80",
          4972 => x"84",
          4973 => x"0d",
          4974 => x"2e",
          4975 => x"b7",
          4976 => x"fd",
          4977 => x"2e",
          4978 => x"78",
          4979 => x"89",
          4980 => x"0b",
          4981 => x"0c",
          4982 => x"33",
          4983 => x"33",
          4984 => x"33",
          4985 => x"05",
          4986 => x"84",
          4987 => x"33",
          4988 => x"80",
          4989 => x"b8",
          4990 => x"fa",
          4991 => x"fa",
          4992 => x"71",
          4993 => x"5f",
          4994 => x"83",
          4995 => x"34",
          4996 => x"33",
          4997 => x"19",
          4998 => x"fa",
          4999 => x"c7",
          5000 => x"34",
          5001 => x"33",
          5002 => x"06",
          5003 => x"22",
          5004 => x"33",
          5005 => x"11",
          5006 => x"58",
          5007 => x"b0",
          5008 => x"99",
          5009 => x"81",
          5010 => x"81",
          5011 => x"60",
          5012 => x"ca",
          5013 => x"fa",
          5014 => x"0b",
          5015 => x"0c",
          5016 => x"04",
          5017 => x"82",
          5018 => x"9b",
          5019 => x"38",
          5020 => x"09",
          5021 => x"a8",
          5022 => x"83",
          5023 => x"80",
          5024 => x"84",
          5025 => x"0d",
          5026 => x"2e",
          5027 => x"d0",
          5028 => x"89",
          5029 => x"38",
          5030 => x"33",
          5031 => x"57",
          5032 => x"84",
          5033 => x"ba",
          5034 => x"77",
          5035 => x"59",
          5036 => x"ba",
          5037 => x"80",
          5038 => x"84",
          5039 => x"0d",
          5040 => x"2e",
          5041 => x"80",
          5042 => x"80",
          5043 => x"f8",
          5044 => x"b4",
          5045 => x"b5",
          5046 => x"29",
          5047 => x"40",
          5048 => x"19",
          5049 => x"a0",
          5050 => x"84",
          5051 => x"83",
          5052 => x"83",
          5053 => x"72",
          5054 => x"41",
          5055 => x"78",
          5056 => x"1f",
          5057 => x"b4",
          5058 => x"29",
          5059 => x"83",
          5060 => x"86",
          5061 => x"1b",
          5062 => x"f8",
          5063 => x"ff",
          5064 => x"b2",
          5065 => x"b5",
          5066 => x"29",
          5067 => x"43",
          5068 => x"fa",
          5069 => x"84",
          5070 => x"34",
          5071 => x"fe",
          5072 => x"52",
          5073 => x"fa",
          5074 => x"83",
          5075 => x"fe",
          5076 => x"b8",
          5077 => x"fa",
          5078 => x"81",
          5079 => x"fa",
          5080 => x"71",
          5081 => x"c7",
          5082 => x"83",
          5083 => x"40",
          5084 => x"7e",
          5085 => x"83",
          5086 => x"83",
          5087 => x"5a",
          5088 => x"5c",
          5089 => x"86",
          5090 => x"81",
          5091 => x"1a",
          5092 => x"fc",
          5093 => x"56",
          5094 => x"b5",
          5095 => x"39",
          5096 => x"ba",
          5097 => x"0b",
          5098 => x"34",
          5099 => x"ba",
          5100 => x"0b",
          5101 => x"34",
          5102 => x"ba",
          5103 => x"0b",
          5104 => x"0c",
          5105 => x"04",
          5106 => x"33",
          5107 => x"34",
          5108 => x"33",
          5109 => x"34",
          5110 => x"33",
          5111 => x"34",
          5112 => x"ba",
          5113 => x"0b",
          5114 => x"0c",
          5115 => x"04",
          5116 => x"2e",
          5117 => x"fa",
          5118 => x"fa",
          5119 => x"b8",
          5120 => x"81",
          5121 => x"fa",
          5122 => x"81",
          5123 => x"75",
          5124 => x"c7",
          5125 => x"83",
          5126 => x"5c",
          5127 => x"29",
          5128 => x"ff",
          5129 => x"f9",
          5130 => x"5c",
          5131 => x"5b",
          5132 => x"2e",
          5133 => x"78",
          5134 => x"ff",
          5135 => x"75",
          5136 => x"57",
          5137 => x"b5",
          5138 => x"ff",
          5139 => x"ff",
          5140 => x"ff",
          5141 => x"29",
          5142 => x"5b",
          5143 => x"33",
          5144 => x"80",
          5145 => x"b8",
          5146 => x"fa",
          5147 => x"fa",
          5148 => x"71",
          5149 => x"5e",
          5150 => x"0b",
          5151 => x"18",
          5152 => x"b4",
          5153 => x"29",
          5154 => x"56",
          5155 => x"33",
          5156 => x"80",
          5157 => x"b8",
          5158 => x"81",
          5159 => x"fa",
          5160 => x"fa",
          5161 => x"72",
          5162 => x"5d",
          5163 => x"83",
          5164 => x"7f",
          5165 => x"05",
          5166 => x"70",
          5167 => x"5c",
          5168 => x"26",
          5169 => x"84",
          5170 => x"5a",
          5171 => x"38",
          5172 => x"77",
          5173 => x"34",
          5174 => x"33",
          5175 => x"06",
          5176 => x"56",
          5177 => x"78",
          5178 => x"d8",
          5179 => x"2e",
          5180 => x"78",
          5181 => x"a8",
          5182 => x"84",
          5183 => x"83",
          5184 => x"bf",
          5185 => x"b4",
          5186 => x"38",
          5187 => x"83",
          5188 => x"58",
          5189 => x"80",
          5190 => x"b5",
          5191 => x"81",
          5192 => x"3f",
          5193 => x"bb",
          5194 => x"3d",
          5195 => x"fa",
          5196 => x"b8",
          5197 => x"81",
          5198 => x"fa",
          5199 => x"81",
          5200 => x"75",
          5201 => x"c7",
          5202 => x"83",
          5203 => x"5c",
          5204 => x"29",
          5205 => x"ff",
          5206 => x"f9",
          5207 => x"53",
          5208 => x"5b",
          5209 => x"2e",
          5210 => x"80",
          5211 => x"ff",
          5212 => x"ff",
          5213 => x"ff",
          5214 => x"29",
          5215 => x"40",
          5216 => x"33",
          5217 => x"80",
          5218 => x"b8",
          5219 => x"fa",
          5220 => x"fa",
          5221 => x"71",
          5222 => x"41",
          5223 => x"0b",
          5224 => x"1c",
          5225 => x"b4",
          5226 => x"29",
          5227 => x"83",
          5228 => x"86",
          5229 => x"1a",
          5230 => x"f8",
          5231 => x"ff",
          5232 => x"b2",
          5233 => x"b5",
          5234 => x"29",
          5235 => x"5a",
          5236 => x"fa",
          5237 => x"99",
          5238 => x"60",
          5239 => x"81",
          5240 => x"58",
          5241 => x"81",
          5242 => x"b8",
          5243 => x"77",
          5244 => x"ff",
          5245 => x"83",
          5246 => x"81",
          5247 => x"ff",
          5248 => x"7b",
          5249 => x"a7",
          5250 => x"b4",
          5251 => x"f8",
          5252 => x"b5",
          5253 => x"ff",
          5254 => x"ff",
          5255 => x"ff",
          5256 => x"29",
          5257 => x"43",
          5258 => x"84",
          5259 => x"86",
          5260 => x"1b",
          5261 => x"f8",
          5262 => x"b5",
          5263 => x"b2",
          5264 => x"29",
          5265 => x"5e",
          5266 => x"83",
          5267 => x"34",
          5268 => x"33",
          5269 => x"1e",
          5270 => x"fa",
          5271 => x"c7",
          5272 => x"34",
          5273 => x"33",
          5274 => x"06",
          5275 => x"22",
          5276 => x"33",
          5277 => x"11",
          5278 => x"40",
          5279 => x"b0",
          5280 => x"d6",
          5281 => x"81",
          5282 => x"ff",
          5283 => x"79",
          5284 => x"d6",
          5285 => x"fa",
          5286 => x"df",
          5287 => x"84",
          5288 => x"80",
          5289 => x"84",
          5290 => x"0d",
          5291 => x"b6",
          5292 => x"84",
          5293 => x"33",
          5294 => x"fa",
          5295 => x"81",
          5296 => x"ff",
          5297 => x"ca",
          5298 => x"84",
          5299 => x"80",
          5300 => x"84",
          5301 => x"0d",
          5302 => x"b6",
          5303 => x"84",
          5304 => x"33",
          5305 => x"fa",
          5306 => x"b8",
          5307 => x"fa",
          5308 => x"5b",
          5309 => x"fc",
          5310 => x"ba",
          5311 => x"3d",
          5312 => x"d8",
          5313 => x"88",
          5314 => x"bb",
          5315 => x"2e",
          5316 => x"84",
          5317 => x"81",
          5318 => x"75",
          5319 => x"34",
          5320 => x"fe",
          5321 => x"80",
          5322 => x"61",
          5323 => x"05",
          5324 => x"39",
          5325 => x"17",
          5326 => x"b9",
          5327 => x"7b",
          5328 => x"b4",
          5329 => x"f8",
          5330 => x"b5",
          5331 => x"5c",
          5332 => x"84",
          5333 => x"83",
          5334 => x"83",
          5335 => x"72",
          5336 => x"41",
          5337 => x"b9",
          5338 => x"7f",
          5339 => x"80",
          5340 => x"b8",
          5341 => x"fa",
          5342 => x"fa",
          5343 => x"71",
          5344 => x"43",
          5345 => x"83",
          5346 => x"34",
          5347 => x"33",
          5348 => x"1b",
          5349 => x"fa",
          5350 => x"86",
          5351 => x"05",
          5352 => x"f8",
          5353 => x"ff",
          5354 => x"b2",
          5355 => x"b5",
          5356 => x"29",
          5357 => x"5a",
          5358 => x"fa",
          5359 => x"99",
          5360 => x"81",
          5361 => x"ff",
          5362 => x"60",
          5363 => x"a2",
          5364 => x"f9",
          5365 => x"90",
          5366 => x"1a",
          5367 => x"fa",
          5368 => x"0b",
          5369 => x"0c",
          5370 => x"33",
          5371 => x"2e",
          5372 => x"84",
          5373 => x"56",
          5374 => x"38",
          5375 => x"51",
          5376 => x"80",
          5377 => x"84",
          5378 => x"0d",
          5379 => x"ec",
          5380 => x"b4",
          5381 => x"ed",
          5382 => x"b5",
          5383 => x"ee",
          5384 => x"83",
          5385 => x"ff",
          5386 => x"fa",
          5387 => x"ba",
          5388 => x"fa",
          5389 => x"ba",
          5390 => x"fa",
          5391 => x"ba",
          5392 => x"9e",
          5393 => x"85",
          5394 => x"80",
          5395 => x"38",
          5396 => x"22",
          5397 => x"2e",
          5398 => x"ff",
          5399 => x"fa",
          5400 => x"05",
          5401 => x"b4",
          5402 => x"54",
          5403 => x"e5",
          5404 => x"3d",
          5405 => x"fe",
          5406 => x"76",
          5407 => x"aa",
          5408 => x"84",
          5409 => x"06",
          5410 => x"33",
          5411 => x"41",
          5412 => x"fe",
          5413 => x"52",
          5414 => x"51",
          5415 => x"3f",
          5416 => x"80",
          5417 => x"85",
          5418 => x"79",
          5419 => x"5b",
          5420 => x"fe",
          5421 => x"10",
          5422 => x"05",
          5423 => x"57",
          5424 => x"26",
          5425 => x"75",
          5426 => x"c8",
          5427 => x"7e",
          5428 => x"ba",
          5429 => x"7d",
          5430 => x"a4",
          5431 => x"b4",
          5432 => x"d9",
          5433 => x"31",
          5434 => x"9f",
          5435 => x"5a",
          5436 => x"5c",
          5437 => x"b4",
          5438 => x"39",
          5439 => x"33",
          5440 => x"2e",
          5441 => x"84",
          5442 => x"ff",
          5443 => x"ff",
          5444 => x"f8",
          5445 => x"5f",
          5446 => x"fd",
          5447 => x"83",
          5448 => x"fd",
          5449 => x"0b",
          5450 => x"34",
          5451 => x"33",
          5452 => x"06",
          5453 => x"80",
          5454 => x"38",
          5455 => x"75",
          5456 => x"34",
          5457 => x"80",
          5458 => x"b5",
          5459 => x"b4",
          5460 => x"f7",
          5461 => x"57",
          5462 => x"25",
          5463 => x"81",
          5464 => x"83",
          5465 => x"fc",
          5466 => x"ba",
          5467 => x"7f",
          5468 => x"e0",
          5469 => x"b5",
          5470 => x"d9",
          5471 => x"31",
          5472 => x"9f",
          5473 => x"5a",
          5474 => x"5a",
          5475 => x"b5",
          5476 => x"39",
          5477 => x"33",
          5478 => x"2e",
          5479 => x"84",
          5480 => x"41",
          5481 => x"09",
          5482 => x"b6",
          5483 => x"f8",
          5484 => x"b5",
          5485 => x"b4",
          5486 => x"29",
          5487 => x"a0",
          5488 => x"fa",
          5489 => x"51",
          5490 => x"60",
          5491 => x"83",
          5492 => x"83",
          5493 => x"87",
          5494 => x"06",
          5495 => x"5d",
          5496 => x"80",
          5497 => x"38",
          5498 => x"f9",
          5499 => x"f2",
          5500 => x"85",
          5501 => x"80",
          5502 => x"38",
          5503 => x"22",
          5504 => x"2e",
          5505 => x"fb",
          5506 => x"0b",
          5507 => x"34",
          5508 => x"84",
          5509 => x"56",
          5510 => x"90",
          5511 => x"ba",
          5512 => x"fa",
          5513 => x"7c",
          5514 => x"f8",
          5515 => x"59",
          5516 => x"7d",
          5517 => x"75",
          5518 => x"fa",
          5519 => x"a2",
          5520 => x"85",
          5521 => x"80",
          5522 => x"38",
          5523 => x"33",
          5524 => x"33",
          5525 => x"84",
          5526 => x"ff",
          5527 => x"56",
          5528 => x"83",
          5529 => x"76",
          5530 => x"34",
          5531 => x"83",
          5532 => x"fe",
          5533 => x"80",
          5534 => x"85",
          5535 => x"76",
          5536 => x"c7",
          5537 => x"84",
          5538 => x"70",
          5539 => x"83",
          5540 => x"fe",
          5541 => x"81",
          5542 => x"ff",
          5543 => x"85",
          5544 => x"58",
          5545 => x"0b",
          5546 => x"33",
          5547 => x"80",
          5548 => x"84",
          5549 => x"56",
          5550 => x"83",
          5551 => x"81",
          5552 => x"ff",
          5553 => x"f3",
          5554 => x"39",
          5555 => x"33",
          5556 => x"27",
          5557 => x"84",
          5558 => x"ff",
          5559 => x"ff",
          5560 => x"d9",
          5561 => x"70",
          5562 => x"84",
          5563 => x"70",
          5564 => x"ff",
          5565 => x"52",
          5566 => x"5c",
          5567 => x"83",
          5568 => x"79",
          5569 => x"23",
          5570 => x"06",
          5571 => x"5f",
          5572 => x"83",
          5573 => x"76",
          5574 => x"34",
          5575 => x"33",
          5576 => x"40",
          5577 => x"f9",
          5578 => x"56",
          5579 => x"b5",
          5580 => x"39",
          5581 => x"33",
          5582 => x"2e",
          5583 => x"84",
          5584 => x"84",
          5585 => x"40",
          5586 => x"26",
          5587 => x"83",
          5588 => x"84",
          5589 => x"70",
          5590 => x"83",
          5591 => x"71",
          5592 => x"86",
          5593 => x"05",
          5594 => x"22",
          5595 => x"7e",
          5596 => x"83",
          5597 => x"83",
          5598 => x"46",
          5599 => x"5f",
          5600 => x"2e",
          5601 => x"79",
          5602 => x"06",
          5603 => x"5d",
          5604 => x"24",
          5605 => x"84",
          5606 => x"56",
          5607 => x"8e",
          5608 => x"16",
          5609 => x"fa",
          5610 => x"81",
          5611 => x"7c",
          5612 => x"80",
          5613 => x"e5",
          5614 => x"f7",
          5615 => x"76",
          5616 => x"38",
          5617 => x"75",
          5618 => x"34",
          5619 => x"06",
          5620 => x"22",
          5621 => x"5a",
          5622 => x"90",
          5623 => x"31",
          5624 => x"81",
          5625 => x"71",
          5626 => x"5b",
          5627 => x"c7",
          5628 => x"86",
          5629 => x"7f",
          5630 => x"7f",
          5631 => x"71",
          5632 => x"42",
          5633 => x"79",
          5634 => x"d6",
          5635 => x"d6",
          5636 => x"e0",
          5637 => x"84",
          5638 => x"33",
          5639 => x"05",
          5640 => x"70",
          5641 => x"33",
          5642 => x"05",
          5643 => x"18",
          5644 => x"33",
          5645 => x"33",
          5646 => x"1d",
          5647 => x"58",
          5648 => x"f7",
          5649 => x"e0",
          5650 => x"84",
          5651 => x"33",
          5652 => x"05",
          5653 => x"70",
          5654 => x"33",
          5655 => x"05",
          5656 => x"18",
          5657 => x"33",
          5658 => x"33",
          5659 => x"1d",
          5660 => x"58",
          5661 => x"ff",
          5662 => x"e6",
          5663 => x"85",
          5664 => x"80",
          5665 => x"38",
          5666 => x"ba",
          5667 => x"d8",
          5668 => x"ce",
          5669 => x"84",
          5670 => x"ff",
          5671 => x"85",
          5672 => x"40",
          5673 => x"2e",
          5674 => x"ba",
          5675 => x"75",
          5676 => x"81",
          5677 => x"38",
          5678 => x"33",
          5679 => x"ff",
          5680 => x"b4",
          5681 => x"5c",
          5682 => x"2e",
          5683 => x"84",
          5684 => x"40",
          5685 => x"f6",
          5686 => x"81",
          5687 => x"60",
          5688 => x"fe",
          5689 => x"26",
          5690 => x"07",
          5691 => x"f2",
          5692 => x"10",
          5693 => x"29",
          5694 => x"c7",
          5695 => x"70",
          5696 => x"86",
          5697 => x"05",
          5698 => x"58",
          5699 => x"8b",
          5700 => x"83",
          5701 => x"8b",
          5702 => x"fa",
          5703 => x"98",
          5704 => x"2b",
          5705 => x"2b",
          5706 => x"79",
          5707 => x"5f",
          5708 => x"27",
          5709 => x"77",
          5710 => x"59",
          5711 => x"70",
          5712 => x"0c",
          5713 => x"ee",
          5714 => x"f8",
          5715 => x"f7",
          5716 => x"7e",
          5717 => x"60",
          5718 => x"83",
          5719 => x"7d",
          5720 => x"05",
          5721 => x"5a",
          5722 => x"8c",
          5723 => x"31",
          5724 => x"29",
          5725 => x"40",
          5726 => x"57",
          5727 => x"26",
          5728 => x"83",
          5729 => x"84",
          5730 => x"59",
          5731 => x"e0",
          5732 => x"79",
          5733 => x"05",
          5734 => x"17",
          5735 => x"26",
          5736 => x"a0",
          5737 => x"19",
          5738 => x"70",
          5739 => x"34",
          5740 => x"75",
          5741 => x"38",
          5742 => x"ff",
          5743 => x"ff",
          5744 => x"fe",
          5745 => x"fa",
          5746 => x"80",
          5747 => x"84",
          5748 => x"06",
          5749 => x"07",
          5750 => x"7b",
          5751 => x"09",
          5752 => x"38",
          5753 => x"83",
          5754 => x"81",
          5755 => x"ff",
          5756 => x"f5",
          5757 => x"fa",
          5758 => x"5e",
          5759 => x"1e",
          5760 => x"83",
          5761 => x"84",
          5762 => x"83",
          5763 => x"84",
          5764 => x"42",
          5765 => x"fa",
          5766 => x"fa",
          5767 => x"07",
          5768 => x"fa",
          5769 => x"18",
          5770 => x"06",
          5771 => x"fb",
          5772 => x"b0",
          5773 => x"06",
          5774 => x"75",
          5775 => x"34",
          5776 => x"fa",
          5777 => x"fb",
          5778 => x"56",
          5779 => x"b0",
          5780 => x"83",
          5781 => x"81",
          5782 => x"07",
          5783 => x"fa",
          5784 => x"39",
          5785 => x"33",
          5786 => x"90",
          5787 => x"83",
          5788 => x"ff",
          5789 => x"f1",
          5790 => x"b0",
          5791 => x"70",
          5792 => x"59",
          5793 => x"39",
          5794 => x"33",
          5795 => x"56",
          5796 => x"b0",
          5797 => x"39",
          5798 => x"33",
          5799 => x"90",
          5800 => x"83",
          5801 => x"fe",
          5802 => x"fa",
          5803 => x"ef",
          5804 => x"07",
          5805 => x"fa",
          5806 => x"ea",
          5807 => x"b0",
          5808 => x"06",
          5809 => x"56",
          5810 => x"b0",
          5811 => x"39",
          5812 => x"33",
          5813 => x"a0",
          5814 => x"83",
          5815 => x"fe",
          5816 => x"fa",
          5817 => x"fe",
          5818 => x"56",
          5819 => x"b0",
          5820 => x"39",
          5821 => x"33",
          5822 => x"84",
          5823 => x"83",
          5824 => x"fe",
          5825 => x"fa",
          5826 => x"fa",
          5827 => x"56",
          5828 => x"b0",
          5829 => x"39",
          5830 => x"33",
          5831 => x"56",
          5832 => x"b0",
          5833 => x"39",
          5834 => x"33",
          5835 => x"56",
          5836 => x"b0",
          5837 => x"39",
          5838 => x"33",
          5839 => x"56",
          5840 => x"b0",
          5841 => x"39",
          5842 => x"33",
          5843 => x"80",
          5844 => x"75",
          5845 => x"34",
          5846 => x"83",
          5847 => x"81",
          5848 => x"07",
          5849 => x"fa",
          5850 => x"ba",
          5851 => x"83",
          5852 => x"80",
          5853 => x"d2",
          5854 => x"ff",
          5855 => x"ec",
          5856 => x"b4",
          5857 => x"ed",
          5858 => x"b5",
          5859 => x"ee",
          5860 => x"83",
          5861 => x"80",
          5862 => x"80",
          5863 => x"39",
          5864 => x"ba",
          5865 => x"0b",
          5866 => x"0c",
          5867 => x"04",
          5868 => x"b5",
          5869 => x"b5",
          5870 => x"ff",
          5871 => x"05",
          5872 => x"39",
          5873 => x"42",
          5874 => x"11",
          5875 => x"51",
          5876 => x"3f",
          5877 => x"08",
          5878 => x"bb",
          5879 => x"ba",
          5880 => x"0b",
          5881 => x"34",
          5882 => x"bb",
          5883 => x"3d",
          5884 => x"83",
          5885 => x"ef",
          5886 => x"ba",
          5887 => x"11",
          5888 => x"84",
          5889 => x"7b",
          5890 => x"06",
          5891 => x"ca",
          5892 => x"ba",
          5893 => x"80",
          5894 => x"84",
          5895 => x"80",
          5896 => x"b5",
          5897 => x"81",
          5898 => x"3f",
          5899 => x"33",
          5900 => x"06",
          5901 => x"56",
          5902 => x"80",
          5903 => x"b5",
          5904 => x"81",
          5905 => x"3f",
          5906 => x"8a",
          5907 => x"90",
          5908 => x"39",
          5909 => x"33",
          5910 => x"09",
          5911 => x"72",
          5912 => x"57",
          5913 => x"75",
          5914 => x"d9",
          5915 => x"f8",
          5916 => x"60",
          5917 => x"38",
          5918 => x"b5",
          5919 => x"39",
          5920 => x"33",
          5921 => x"09",
          5922 => x"72",
          5923 => x"57",
          5924 => x"83",
          5925 => x"81",
          5926 => x"f7",
          5927 => x"59",
          5928 => x"78",
          5929 => x"38",
          5930 => x"bb",
          5931 => x"f7",
          5932 => x"ff",
          5933 => x"81",
          5934 => x"a6",
          5935 => x"b4",
          5936 => x"f8",
          5937 => x"ff",
          5938 => x"b5",
          5939 => x"29",
          5940 => x"a0",
          5941 => x"fa",
          5942 => x"5f",
          5943 => x"05",
          5944 => x"ff",
          5945 => x"8a",
          5946 => x"44",
          5947 => x"77",
          5948 => x"f5",
          5949 => x"ff",
          5950 => x"11",
          5951 => x"7b",
          5952 => x"38",
          5953 => x"33",
          5954 => x"27",
          5955 => x"ff",
          5956 => x"83",
          5957 => x"7c",
          5958 => x"ff",
          5959 => x"80",
          5960 => x"df",
          5961 => x"f7",
          5962 => x"76",
          5963 => x"38",
          5964 => x"75",
          5965 => x"34",
          5966 => x"06",
          5967 => x"22",
          5968 => x"5a",
          5969 => x"90",
          5970 => x"31",
          5971 => x"81",
          5972 => x"71",
          5973 => x"5f",
          5974 => x"c7",
          5975 => x"86",
          5976 => x"7c",
          5977 => x"7f",
          5978 => x"71",
          5979 => x"41",
          5980 => x"79",
          5981 => x"ea",
          5982 => x"d6",
          5983 => x"e0",
          5984 => x"84",
          5985 => x"33",
          5986 => x"05",
          5987 => x"70",
          5988 => x"33",
          5989 => x"05",
          5990 => x"18",
          5991 => x"33",
          5992 => x"33",
          5993 => x"1d",
          5994 => x"58",
          5995 => x"ec",
          5996 => x"e0",
          5997 => x"84",
          5998 => x"33",
          5999 => x"05",
          6000 => x"70",
          6001 => x"33",
          6002 => x"05",
          6003 => x"18",
          6004 => x"33",
          6005 => x"33",
          6006 => x"1d",
          6007 => x"58",
          6008 => x"ff",
          6009 => x"fa",
          6010 => x"b6",
          6011 => x"84",
          6012 => x"33",
          6013 => x"fa",
          6014 => x"b8",
          6015 => x"fa",
          6016 => x"b8",
          6017 => x"5c",
          6018 => x"e9",
          6019 => x"d2",
          6020 => x"f7",
          6021 => x"ff",
          6022 => x"5c",
          6023 => x"61",
          6024 => x"76",
          6025 => x"fa",
          6026 => x"81",
          6027 => x"19",
          6028 => x"7a",
          6029 => x"80",
          6030 => x"fa",
          6031 => x"b8",
          6032 => x"81",
          6033 => x"12",
          6034 => x"80",
          6035 => x"8d",
          6036 => x"75",
          6037 => x"34",
          6038 => x"83",
          6039 => x"81",
          6040 => x"f8",
          6041 => x"59",
          6042 => x"7f",
          6043 => x"38",
          6044 => x"c5",
          6045 => x"2e",
          6046 => x"f4",
          6047 => x"fa",
          6048 => x"81",
          6049 => x"fa",
          6050 => x"44",
          6051 => x"76",
          6052 => x"81",
          6053 => x"38",
          6054 => x"ff",
          6055 => x"83",
          6056 => x"fd",
          6057 => x"1a",
          6058 => x"fa",
          6059 => x"e7",
          6060 => x"31",
          6061 => x"fa",
          6062 => x"90",
          6063 => x"58",
          6064 => x"26",
          6065 => x"80",
          6066 => x"05",
          6067 => x"fa",
          6068 => x"70",
          6069 => x"34",
          6070 => x"f4",
          6071 => x"76",
          6072 => x"58",
          6073 => x"b0",
          6074 => x"81",
          6075 => x"79",
          6076 => x"38",
          6077 => x"79",
          6078 => x"75",
          6079 => x"23",
          6080 => x"80",
          6081 => x"b4",
          6082 => x"39",
          6083 => x"b2",
          6084 => x"39",
          6085 => x"fa",
          6086 => x"8e",
          6087 => x"83",
          6088 => x"f1",
          6089 => x"fa",
          6090 => x"5a",
          6091 => x"1a",
          6092 => x"80",
          6093 => x"89",
          6094 => x"39",
          6095 => x"02",
          6096 => x"84",
          6097 => x"54",
          6098 => x"2e",
          6099 => x"51",
          6100 => x"80",
          6101 => x"84",
          6102 => x"0d",
          6103 => x"73",
          6104 => x"3f",
          6105 => x"bb",
          6106 => x"3d",
          6107 => x"3d",
          6108 => x"05",
          6109 => x"0b",
          6110 => x"33",
          6111 => x"06",
          6112 => x"11",
          6113 => x"55",
          6114 => x"2e",
          6115 => x"81",
          6116 => x"83",
          6117 => x"74",
          6118 => x"bb",
          6119 => x"3d",
          6120 => x"f8",
          6121 => x"82",
          6122 => x"2e",
          6123 => x"73",
          6124 => x"71",
          6125 => x"70",
          6126 => x"5d",
          6127 => x"83",
          6128 => x"ff",
          6129 => x"7b",
          6130 => x"81",
          6131 => x"7b",
          6132 => x"32",
          6133 => x"80",
          6134 => x"5c",
          6135 => x"80",
          6136 => x"38",
          6137 => x"33",
          6138 => x"33",
          6139 => x"33",
          6140 => x"12",
          6141 => x"80",
          6142 => x"b2",
          6143 => x"5d",
          6144 => x"05",
          6145 => x"ff",
          6146 => x"89",
          6147 => x"55",
          6148 => x"2e",
          6149 => x"81",
          6150 => x"87",
          6151 => x"34",
          6152 => x"c0",
          6153 => x"87",
          6154 => x"08",
          6155 => x"2e",
          6156 => x"8e",
          6157 => x"57",
          6158 => x"b4",
          6159 => x"14",
          6160 => x"06",
          6161 => x"f9",
          6162 => x"38",
          6163 => x"f8",
          6164 => x"70",
          6165 => x"83",
          6166 => x"33",
          6167 => x"72",
          6168 => x"c1",
          6169 => x"ff",
          6170 => x"38",
          6171 => x"b8",
          6172 => x"81",
          6173 => x"79",
          6174 => x"85",
          6175 => x"83",
          6176 => x"34",
          6177 => x"14",
          6178 => x"ae",
          6179 => x"14",
          6180 => x"06",
          6181 => x"74",
          6182 => x"38",
          6183 => x"33",
          6184 => x"70",
          6185 => x"56",
          6186 => x"f8",
          6187 => x"81",
          6188 => x"86",
          6189 => x"70",
          6190 => x"54",
          6191 => x"2e",
          6192 => x"81",
          6193 => x"dd",
          6194 => x"81",
          6195 => x"80",
          6196 => x"38",
          6197 => x"f8",
          6198 => x"0b",
          6199 => x"33",
          6200 => x"08",
          6201 => x"33",
          6202 => x"e0",
          6203 => x"df",
          6204 => x"42",
          6205 => x"56",
          6206 => x"16",
          6207 => x"81",
          6208 => x"38",
          6209 => x"16",
          6210 => x"80",
          6211 => x"38",
          6212 => x"16",
          6213 => x"81",
          6214 => x"38",
          6215 => x"16",
          6216 => x"81",
          6217 => x"81",
          6218 => x"73",
          6219 => x"8d",
          6220 => x"cc",
          6221 => x"72",
          6222 => x"da",
          6223 => x"ff",
          6224 => x"81",
          6225 => x"8c",
          6226 => x"cc",
          6227 => x"81",
          6228 => x"80",
          6229 => x"d8",
          6230 => x"05",
          6231 => x"9c",
          6232 => x"73",
          6233 => x"ec",
          6234 => x"87",
          6235 => x"08",
          6236 => x"0c",
          6237 => x"70",
          6238 => x"57",
          6239 => x"27",
          6240 => x"76",
          6241 => x"34",
          6242 => x"e0",
          6243 => x"19",
          6244 => x"26",
          6245 => x"72",
          6246 => x"c9",
          6247 => x"79",
          6248 => x"f9",
          6249 => x"73",
          6250 => x"38",
          6251 => x"87",
          6252 => x"08",
          6253 => x"7d",
          6254 => x"38",
          6255 => x"f9",
          6256 => x"54",
          6257 => x"83",
          6258 => x"73",
          6259 => x"34",
          6260 => x"9c",
          6261 => x"8c",
          6262 => x"ff",
          6263 => x"81",
          6264 => x"83",
          6265 => x"33",
          6266 => x"80",
          6267 => x"34",
          6268 => x"fc",
          6269 => x"f8",
          6270 => x"72",
          6271 => x"9c",
          6272 => x"2e",
          6273 => x"80",
          6274 => x"81",
          6275 => x"8a",
          6276 => x"fe",
          6277 => x"74",
          6278 => x"59",
          6279 => x"9b",
          6280 => x"2e",
          6281 => x"83",
          6282 => x"81",
          6283 => x"38",
          6284 => x"80",
          6285 => x"81",
          6286 => x"87",
          6287 => x"98",
          6288 => x"72",
          6289 => x"38",
          6290 => x"9c",
          6291 => x"70",
          6292 => x"76",
          6293 => x"06",
          6294 => x"71",
          6295 => x"53",
          6296 => x"80",
          6297 => x"38",
          6298 => x"10",
          6299 => x"76",
          6300 => x"78",
          6301 => x"94",
          6302 => x"5b",
          6303 => x"87",
          6304 => x"08",
          6305 => x"0c",
          6306 => x"39",
          6307 => x"81",
          6308 => x"38",
          6309 => x"06",
          6310 => x"39",
          6311 => x"9b",
          6312 => x"2e",
          6313 => x"80",
          6314 => x"fa",
          6315 => x"72",
          6316 => x"e8",
          6317 => x"32",
          6318 => x"80",
          6319 => x"40",
          6320 => x"8a",
          6321 => x"2e",
          6322 => x"f9",
          6323 => x"ff",
          6324 => x"38",
          6325 => x"10",
          6326 => x"f9",
          6327 => x"33",
          6328 => x"7c",
          6329 => x"38",
          6330 => x"81",
          6331 => x"57",
          6332 => x"e2",
          6333 => x"fb",
          6334 => x"80",
          6335 => x"38",
          6336 => x"33",
          6337 => x"91",
          6338 => x"ff",
          6339 => x"51",
          6340 => x"78",
          6341 => x"0c",
          6342 => x"04",
          6343 => x"81",
          6344 => x"f6",
          6345 => x"ff",
          6346 => x"83",
          6347 => x"33",
          6348 => x"7a",
          6349 => x"15",
          6350 => x"39",
          6351 => x"f8",
          6352 => x"ff",
          6353 => x"b8",
          6354 => x"0b",
          6355 => x"15",
          6356 => x"39",
          6357 => x"06",
          6358 => x"ff",
          6359 => x"38",
          6360 => x"16",
          6361 => x"75",
          6362 => x"38",
          6363 => x"06",
          6364 => x"2e",
          6365 => x"fb",
          6366 => x"f8",
          6367 => x"fa",
          6368 => x"98",
          6369 => x"55",
          6370 => x"fb",
          6371 => x"c0",
          6372 => x"83",
          6373 => x"76",
          6374 => x"59",
          6375 => x"ff",
          6376 => x"b8",
          6377 => x"ca",
          6378 => x"f8",
          6379 => x"09",
          6380 => x"72",
          6381 => x"72",
          6382 => x"34",
          6383 => x"f8",
          6384 => x"f8",
          6385 => x"f8",
          6386 => x"83",
          6387 => x"83",
          6388 => x"5d",
          6389 => x"5c",
          6390 => x"9c",
          6391 => x"2e",
          6392 => x"fc",
          6393 => x"59",
          6394 => x"fc",
          6395 => x"81",
          6396 => x"06",
          6397 => x"fd",
          6398 => x"76",
          6399 => x"54",
          6400 => x"80",
          6401 => x"fb",
          6402 => x"75",
          6403 => x"54",
          6404 => x"fb",
          6405 => x"f7",
          6406 => x"0b",
          6407 => x"33",
          6408 => x"83",
          6409 => x"73",
          6410 => x"34",
          6411 => x"95",
          6412 => x"83",
          6413 => x"84",
          6414 => x"38",
          6415 => x"f8",
          6416 => x"ff",
          6417 => x"f7",
          6418 => x"ff",
          6419 => x"57",
          6420 => x"79",
          6421 => x"80",
          6422 => x"fa",
          6423 => x"81",
          6424 => x"15",
          6425 => x"73",
          6426 => x"80",
          6427 => x"fa",
          6428 => x"b8",
          6429 => x"81",
          6430 => x"ff",
          6431 => x"75",
          6432 => x"80",
          6433 => x"fa",
          6434 => x"59",
          6435 => x"81",
          6436 => x"ff",
          6437 => x"ff",
          6438 => x"39",
          6439 => x"95",
          6440 => x"08",
          6441 => x"e8",
          6442 => x"9d",
          6443 => x"83",
          6444 => x"83",
          6445 => x"59",
          6446 => x"80",
          6447 => x"51",
          6448 => x"82",
          6449 => x"fa",
          6450 => x"0b",
          6451 => x"08",
          6452 => x"a3",
          6453 => x"13",
          6454 => x"90",
          6455 => x"e0",
          6456 => x"0b",
          6457 => x"08",
          6458 => x"0b",
          6459 => x"80",
          6460 => x"80",
          6461 => x"c0",
          6462 => x"83",
          6463 => x"55",
          6464 => x"05",
          6465 => x"98",
          6466 => x"87",
          6467 => x"08",
          6468 => x"2e",
          6469 => x"14",
          6470 => x"98",
          6471 => x"52",
          6472 => x"87",
          6473 => x"fe",
          6474 => x"87",
          6475 => x"08",
          6476 => x"70",
          6477 => x"c8",
          6478 => x"71",
          6479 => x"c0",
          6480 => x"98",
          6481 => x"ce",
          6482 => x"87",
          6483 => x"08",
          6484 => x"98",
          6485 => x"74",
          6486 => x"38",
          6487 => x"87",
          6488 => x"08",
          6489 => x"73",
          6490 => x"71",
          6491 => x"db",
          6492 => x"98",
          6493 => x"72",
          6494 => x"38",
          6495 => x"55",
          6496 => x"81",
          6497 => x"53",
          6498 => x"98",
          6499 => x"ff",
          6500 => x"fe",
          6501 => x"ff",
          6502 => x"76",
          6503 => x"0c",
          6504 => x"04",
          6505 => x"bb",
          6506 => x"3d",
          6507 => x"3d",
          6508 => x"84",
          6509 => x"33",
          6510 => x"0b",
          6511 => x"08",
          6512 => x"87",
          6513 => x"06",
          6514 => x"2a",
          6515 => x"55",
          6516 => x"15",
          6517 => x"2a",
          6518 => x"15",
          6519 => x"2a",
          6520 => x"15",
          6521 => x"15",
          6522 => x"90",
          6523 => x"82",
          6524 => x"f5",
          6525 => x"80",
          6526 => x"85",
          6527 => x"90",
          6528 => x"fe",
          6529 => x"34",
          6530 => x"90",
          6531 => x"87",
          6532 => x"08",
          6533 => x"08",
          6534 => x"90",
          6535 => x"c0",
          6536 => x"52",
          6537 => x"9c",
          6538 => x"72",
          6539 => x"81",
          6540 => x"c0",
          6541 => x"56",
          6542 => x"27",
          6543 => x"81",
          6544 => x"38",
          6545 => x"a4",
          6546 => x"55",
          6547 => x"80",
          6548 => x"55",
          6549 => x"80",
          6550 => x"c0",
          6551 => x"80",
          6552 => x"53",
          6553 => x"9c",
          6554 => x"c0",
          6555 => x"55",
          6556 => x"f6",
          6557 => x"33",
          6558 => x"9c",
          6559 => x"70",
          6560 => x"38",
          6561 => x"2e",
          6562 => x"c0",
          6563 => x"55",
          6564 => x"83",
          6565 => x"71",
          6566 => x"70",
          6567 => x"57",
          6568 => x"2e",
          6569 => x"74",
          6570 => x"52",
          6571 => x"38",
          6572 => x"81",
          6573 => x"75",
          6574 => x"c6",
          6575 => x"80",
          6576 => x"52",
          6577 => x"92",
          6578 => x"81",
          6579 => x"71",
          6580 => x"53",
          6581 => x"26",
          6582 => x"84",
          6583 => x"88",
          6584 => x"81",
          6585 => x"84",
          6586 => x"0d",
          6587 => x"c2",
          6588 => x"0d",
          6589 => x"05",
          6590 => x"56",
          6591 => x"83",
          6592 => x"77",
          6593 => x"fc",
          6594 => x"70",
          6595 => x"07",
          6596 => x"57",
          6597 => x"34",
          6598 => x"51",
          6599 => x"34",
          6600 => x"52",
          6601 => x"34",
          6602 => x"34",
          6603 => x"90",
          6604 => x"11",
          6605 => x"56",
          6606 => x"70",
          6607 => x"38",
          6608 => x"05",
          6609 => x"70",
          6610 => x"34",
          6611 => x"f0",
          6612 => x"90",
          6613 => x"82",
          6614 => x"f5",
          6615 => x"80",
          6616 => x"85",
          6617 => x"90",
          6618 => x"fe",
          6619 => x"34",
          6620 => x"90",
          6621 => x"87",
          6622 => x"08",
          6623 => x"08",
          6624 => x"90",
          6625 => x"c0",
          6626 => x"52",
          6627 => x"9c",
          6628 => x"72",
          6629 => x"81",
          6630 => x"c0",
          6631 => x"56",
          6632 => x"27",
          6633 => x"81",
          6634 => x"38",
          6635 => x"a4",
          6636 => x"55",
          6637 => x"80",
          6638 => x"55",
          6639 => x"80",
          6640 => x"c0",
          6641 => x"80",
          6642 => x"53",
          6643 => x"9c",
          6644 => x"c0",
          6645 => x"55",
          6646 => x"f6",
          6647 => x"33",
          6648 => x"9c",
          6649 => x"70",
          6650 => x"38",
          6651 => x"2e",
          6652 => x"c0",
          6653 => x"55",
          6654 => x"83",
          6655 => x"71",
          6656 => x"70",
          6657 => x"57",
          6658 => x"2e",
          6659 => x"81",
          6660 => x"71",
          6661 => x"74",
          6662 => x"ff",
          6663 => x"80",
          6664 => x"81",
          6665 => x"bb",
          6666 => x"3d",
          6667 => x"51",
          6668 => x"3d",
          6669 => x"90",
          6670 => x"d0",
          6671 => x"0b",
          6672 => x"08",
          6673 => x"0b",
          6674 => x"80",
          6675 => x"80",
          6676 => x"c0",
          6677 => x"83",
          6678 => x"56",
          6679 => x"05",
          6680 => x"98",
          6681 => x"87",
          6682 => x"08",
          6683 => x"2e",
          6684 => x"15",
          6685 => x"98",
          6686 => x"52",
          6687 => x"87",
          6688 => x"fe",
          6689 => x"87",
          6690 => x"08",
          6691 => x"70",
          6692 => x"c8",
          6693 => x"71",
          6694 => x"c0",
          6695 => x"98",
          6696 => x"ce",
          6697 => x"87",
          6698 => x"08",
          6699 => x"98",
          6700 => x"70",
          6701 => x"38",
          6702 => x"87",
          6703 => x"08",
          6704 => x"73",
          6705 => x"71",
          6706 => x"db",
          6707 => x"98",
          6708 => x"72",
          6709 => x"38",
          6710 => x"53",
          6711 => x"81",
          6712 => x"52",
          6713 => x"8a",
          6714 => x"ff",
          6715 => x"fe",
          6716 => x"39",
          6717 => x"83",
          6718 => x"fe",
          6719 => x"82",
          6720 => x"f9",
          6721 => x"ba",
          6722 => x"71",
          6723 => x"70",
          6724 => x"06",
          6725 => x"73",
          6726 => x"81",
          6727 => x"8b",
          6728 => x"2b",
          6729 => x"70",
          6730 => x"33",
          6731 => x"71",
          6732 => x"5c",
          6733 => x"53",
          6734 => x"52",
          6735 => x"80",
          6736 => x"af",
          6737 => x"82",
          6738 => x"12",
          6739 => x"2b",
          6740 => x"07",
          6741 => x"33",
          6742 => x"71",
          6743 => x"90",
          6744 => x"53",
          6745 => x"56",
          6746 => x"24",
          6747 => x"84",
          6748 => x"14",
          6749 => x"2b",
          6750 => x"07",
          6751 => x"88",
          6752 => x"56",
          6753 => x"13",
          6754 => x"ff",
          6755 => x"87",
          6756 => x"ba",
          6757 => x"17",
          6758 => x"85",
          6759 => x"88",
          6760 => x"88",
          6761 => x"59",
          6762 => x"84",
          6763 => x"85",
          6764 => x"ba",
          6765 => x"52",
          6766 => x"13",
          6767 => x"87",
          6768 => x"ba",
          6769 => x"74",
          6770 => x"73",
          6771 => x"84",
          6772 => x"16",
          6773 => x"12",
          6774 => x"2b",
          6775 => x"80",
          6776 => x"2a",
          6777 => x"52",
          6778 => x"75",
          6779 => x"89",
          6780 => x"86",
          6781 => x"13",
          6782 => x"2b",
          6783 => x"07",
          6784 => x"16",
          6785 => x"33",
          6786 => x"07",
          6787 => x"58",
          6788 => x"53",
          6789 => x"84",
          6790 => x"85",
          6791 => x"ba",
          6792 => x"16",
          6793 => x"85",
          6794 => x"8b",
          6795 => x"2b",
          6796 => x"5a",
          6797 => x"86",
          6798 => x"13",
          6799 => x"2b",
          6800 => x"2a",
          6801 => x"52",
          6802 => x"34",
          6803 => x"34",
          6804 => x"08",
          6805 => x"81",
          6806 => x"88",
          6807 => x"ff",
          6808 => x"88",
          6809 => x"54",
          6810 => x"34",
          6811 => x"34",
          6812 => x"08",
          6813 => x"33",
          6814 => x"71",
          6815 => x"83",
          6816 => x"05",
          6817 => x"12",
          6818 => x"2b",
          6819 => x"2b",
          6820 => x"06",
          6821 => x"88",
          6822 => x"53",
          6823 => x"57",
          6824 => x"82",
          6825 => x"83",
          6826 => x"ba",
          6827 => x"17",
          6828 => x"12",
          6829 => x"2b",
          6830 => x"07",
          6831 => x"33",
          6832 => x"71",
          6833 => x"81",
          6834 => x"70",
          6835 => x"52",
          6836 => x"57",
          6837 => x"73",
          6838 => x"14",
          6839 => x"f4",
          6840 => x"82",
          6841 => x"12",
          6842 => x"2b",
          6843 => x"07",
          6844 => x"33",
          6845 => x"71",
          6846 => x"90",
          6847 => x"53",
          6848 => x"57",
          6849 => x"80",
          6850 => x"38",
          6851 => x"13",
          6852 => x"2b",
          6853 => x"80",
          6854 => x"2a",
          6855 => x"76",
          6856 => x"81",
          6857 => x"ba",
          6858 => x"17",
          6859 => x"12",
          6860 => x"2b",
          6861 => x"07",
          6862 => x"14",
          6863 => x"33",
          6864 => x"07",
          6865 => x"57",
          6866 => x"58",
          6867 => x"72",
          6868 => x"75",
          6869 => x"89",
          6870 => x"f9",
          6871 => x"84",
          6872 => x"58",
          6873 => x"2e",
          6874 => x"80",
          6875 => x"77",
          6876 => x"3f",
          6877 => x"04",
          6878 => x"0b",
          6879 => x"0c",
          6880 => x"84",
          6881 => x"82",
          6882 => x"76",
          6883 => x"f4",
          6884 => x"ed",
          6885 => x"f4",
          6886 => x"75",
          6887 => x"81",
          6888 => x"ba",
          6889 => x"76",
          6890 => x"81",
          6891 => x"34",
          6892 => x"08",
          6893 => x"17",
          6894 => x"87",
          6895 => x"ba",
          6896 => x"ba",
          6897 => x"05",
          6898 => x"07",
          6899 => x"ff",
          6900 => x"2a",
          6901 => x"56",
          6902 => x"34",
          6903 => x"34",
          6904 => x"22",
          6905 => x"10",
          6906 => x"08",
          6907 => x"55",
          6908 => x"15",
          6909 => x"83",
          6910 => x"ee",
          6911 => x"0d",
          6912 => x"53",
          6913 => x"72",
          6914 => x"fb",
          6915 => x"82",
          6916 => x"ff",
          6917 => x"51",
          6918 => x"ff",
          6919 => x"f4",
          6920 => x"33",
          6921 => x"71",
          6922 => x"70",
          6923 => x"58",
          6924 => x"ff",
          6925 => x"2e",
          6926 => x"75",
          6927 => x"17",
          6928 => x"12",
          6929 => x"2b",
          6930 => x"ff",
          6931 => x"31",
          6932 => x"ff",
          6933 => x"27",
          6934 => x"5c",
          6935 => x"74",
          6936 => x"70",
          6937 => x"38",
          6938 => x"58",
          6939 => x"85",
          6940 => x"88",
          6941 => x"5a",
          6942 => x"73",
          6943 => x"2e",
          6944 => x"74",
          6945 => x"76",
          6946 => x"11",
          6947 => x"12",
          6948 => x"2b",
          6949 => x"ff",
          6950 => x"56",
          6951 => x"59",
          6952 => x"83",
          6953 => x"80",
          6954 => x"26",
          6955 => x"78",
          6956 => x"2e",
          6957 => x"72",
          6958 => x"88",
          6959 => x"70",
          6960 => x"11",
          6961 => x"80",
          6962 => x"2a",
          6963 => x"56",
          6964 => x"34",
          6965 => x"34",
          6966 => x"08",
          6967 => x"2a",
          6968 => x"82",
          6969 => x"83",
          6970 => x"ba",
          6971 => x"19",
          6972 => x"12",
          6973 => x"2b",
          6974 => x"2b",
          6975 => x"06",
          6976 => x"83",
          6977 => x"70",
          6978 => x"58",
          6979 => x"52",
          6980 => x"12",
          6981 => x"ff",
          6982 => x"83",
          6983 => x"ba",
          6984 => x"54",
          6985 => x"72",
          6986 => x"84",
          6987 => x"70",
          6988 => x"33",
          6989 => x"71",
          6990 => x"83",
          6991 => x"05",
          6992 => x"53",
          6993 => x"15",
          6994 => x"15",
          6995 => x"f4",
          6996 => x"55",
          6997 => x"11",
          6998 => x"33",
          6999 => x"07",
          7000 => x"54",
          7001 => x"70",
          7002 => x"71",
          7003 => x"84",
          7004 => x"70",
          7005 => x"33",
          7006 => x"71",
          7007 => x"83",
          7008 => x"05",
          7009 => x"5a",
          7010 => x"15",
          7011 => x"15",
          7012 => x"f4",
          7013 => x"55",
          7014 => x"11",
          7015 => x"33",
          7016 => x"07",
          7017 => x"54",
          7018 => x"70",
          7019 => x"79",
          7020 => x"84",
          7021 => x"18",
          7022 => x"70",
          7023 => x"0c",
          7024 => x"04",
          7025 => x"87",
          7026 => x"8b",
          7027 => x"2b",
          7028 => x"84",
          7029 => x"18",
          7030 => x"2b",
          7031 => x"2a",
          7032 => x"53",
          7033 => x"84",
          7034 => x"85",
          7035 => x"ba",
          7036 => x"19",
          7037 => x"85",
          7038 => x"8b",
          7039 => x"2b",
          7040 => x"86",
          7041 => x"15",
          7042 => x"2b",
          7043 => x"2a",
          7044 => x"52",
          7045 => x"52",
          7046 => x"34",
          7047 => x"34",
          7048 => x"08",
          7049 => x"81",
          7050 => x"88",
          7051 => x"ff",
          7052 => x"88",
          7053 => x"54",
          7054 => x"34",
          7055 => x"34",
          7056 => x"08",
          7057 => x"51",
          7058 => x"f9",
          7059 => x"84",
          7060 => x"58",
          7061 => x"2e",
          7062 => x"54",
          7063 => x"73",
          7064 => x"0c",
          7065 => x"04",
          7066 => x"91",
          7067 => x"84",
          7068 => x"84",
          7069 => x"0d",
          7070 => x"f4",
          7071 => x"f4",
          7072 => x"0b",
          7073 => x"23",
          7074 => x"53",
          7075 => x"ff",
          7076 => x"cb",
          7077 => x"ba",
          7078 => x"76",
          7079 => x"0b",
          7080 => x"84",
          7081 => x"54",
          7082 => x"34",
          7083 => x"15",
          7084 => x"f4",
          7085 => x"86",
          7086 => x"0b",
          7087 => x"84",
          7088 => x"84",
          7089 => x"ff",
          7090 => x"80",
          7091 => x"ff",
          7092 => x"88",
          7093 => x"55",
          7094 => x"17",
          7095 => x"17",
          7096 => x"f0",
          7097 => x"10",
          7098 => x"f4",
          7099 => x"05",
          7100 => x"82",
          7101 => x"0b",
          7102 => x"77",
          7103 => x"2e",
          7104 => x"fe",
          7105 => x"3d",
          7106 => x"41",
          7107 => x"84",
          7108 => x"59",
          7109 => x"61",
          7110 => x"38",
          7111 => x"85",
          7112 => x"80",
          7113 => x"38",
          7114 => x"60",
          7115 => x"7f",
          7116 => x"2a",
          7117 => x"83",
          7118 => x"55",
          7119 => x"ff",
          7120 => x"78",
          7121 => x"70",
          7122 => x"06",
          7123 => x"7a",
          7124 => x"81",
          7125 => x"88",
          7126 => x"75",
          7127 => x"ff",
          7128 => x"10",
          7129 => x"05",
          7130 => x"61",
          7131 => x"81",
          7132 => x"88",
          7133 => x"90",
          7134 => x"2c",
          7135 => x"46",
          7136 => x"43",
          7137 => x"59",
          7138 => x"42",
          7139 => x"85",
          7140 => x"15",
          7141 => x"33",
          7142 => x"07",
          7143 => x"10",
          7144 => x"81",
          7145 => x"98",
          7146 => x"2b",
          7147 => x"53",
          7148 => x"80",
          7149 => x"c9",
          7150 => x"27",
          7151 => x"63",
          7152 => x"62",
          7153 => x"38",
          7154 => x"85",
          7155 => x"1b",
          7156 => x"25",
          7157 => x"63",
          7158 => x"79",
          7159 => x"38",
          7160 => x"33",
          7161 => x"71",
          7162 => x"83",
          7163 => x"11",
          7164 => x"12",
          7165 => x"2b",
          7166 => x"07",
          7167 => x"52",
          7168 => x"58",
          7169 => x"8c",
          7170 => x"1e",
          7171 => x"83",
          7172 => x"8b",
          7173 => x"2b",
          7174 => x"86",
          7175 => x"12",
          7176 => x"2b",
          7177 => x"07",
          7178 => x"14",
          7179 => x"33",
          7180 => x"07",
          7181 => x"59",
          7182 => x"5b",
          7183 => x"5c",
          7184 => x"84",
          7185 => x"85",
          7186 => x"ba",
          7187 => x"17",
          7188 => x"85",
          7189 => x"8b",
          7190 => x"2b",
          7191 => x"86",
          7192 => x"15",
          7193 => x"2b",
          7194 => x"2a",
          7195 => x"52",
          7196 => x"57",
          7197 => x"34",
          7198 => x"34",
          7199 => x"08",
          7200 => x"81",
          7201 => x"88",
          7202 => x"ff",
          7203 => x"88",
          7204 => x"5e",
          7205 => x"34",
          7206 => x"34",
          7207 => x"08",
          7208 => x"11",
          7209 => x"33",
          7210 => x"71",
          7211 => x"74",
          7212 => x"81",
          7213 => x"88",
          7214 => x"88",
          7215 => x"45",
          7216 => x"55",
          7217 => x"34",
          7218 => x"34",
          7219 => x"08",
          7220 => x"33",
          7221 => x"71",
          7222 => x"83",
          7223 => x"05",
          7224 => x"83",
          7225 => x"88",
          7226 => x"88",
          7227 => x"45",
          7228 => x"55",
          7229 => x"1a",
          7230 => x"1a",
          7231 => x"f4",
          7232 => x"82",
          7233 => x"12",
          7234 => x"2b",
          7235 => x"62",
          7236 => x"2b",
          7237 => x"5d",
          7238 => x"05",
          7239 => x"a4",
          7240 => x"f4",
          7241 => x"05",
          7242 => x"1c",
          7243 => x"ff",
          7244 => x"5f",
          7245 => x"81",
          7246 => x"54",
          7247 => x"84",
          7248 => x"0d",
          7249 => x"f4",
          7250 => x"f4",
          7251 => x"0b",
          7252 => x"23",
          7253 => x"53",
          7254 => x"ff",
          7255 => x"c6",
          7256 => x"ba",
          7257 => x"60",
          7258 => x"0b",
          7259 => x"84",
          7260 => x"5d",
          7261 => x"34",
          7262 => x"1e",
          7263 => x"f4",
          7264 => x"86",
          7265 => x"0b",
          7266 => x"84",
          7267 => x"84",
          7268 => x"ff",
          7269 => x"80",
          7270 => x"ff",
          7271 => x"88",
          7272 => x"5b",
          7273 => x"18",
          7274 => x"18",
          7275 => x"f0",
          7276 => x"10",
          7277 => x"f4",
          7278 => x"05",
          7279 => x"82",
          7280 => x"0b",
          7281 => x"84",
          7282 => x"57",
          7283 => x"38",
          7284 => x"82",
          7285 => x"54",
          7286 => x"fe",
          7287 => x"51",
          7288 => x"84",
          7289 => x"84",
          7290 => x"95",
          7291 => x"61",
          7292 => x"f4",
          7293 => x"2b",
          7294 => x"44",
          7295 => x"33",
          7296 => x"71",
          7297 => x"81",
          7298 => x"70",
          7299 => x"44",
          7300 => x"63",
          7301 => x"81",
          7302 => x"84",
          7303 => x"05",
          7304 => x"57",
          7305 => x"19",
          7306 => x"19",
          7307 => x"f4",
          7308 => x"70",
          7309 => x"33",
          7310 => x"07",
          7311 => x"8f",
          7312 => x"74",
          7313 => x"ff",
          7314 => x"88",
          7315 => x"47",
          7316 => x"5d",
          7317 => x"05",
          7318 => x"ff",
          7319 => x"63",
          7320 => x"84",
          7321 => x"1e",
          7322 => x"34",
          7323 => x"34",
          7324 => x"f4",
          7325 => x"05",
          7326 => x"3f",
          7327 => x"bc",
          7328 => x"31",
          7329 => x"ff",
          7330 => x"fa",
          7331 => x"81",
          7332 => x"76",
          7333 => x"ff",
          7334 => x"17",
          7335 => x"33",
          7336 => x"07",
          7337 => x"10",
          7338 => x"81",
          7339 => x"98",
          7340 => x"2b",
          7341 => x"53",
          7342 => x"45",
          7343 => x"25",
          7344 => x"ff",
          7345 => x"78",
          7346 => x"38",
          7347 => x"8b",
          7348 => x"83",
          7349 => x"5b",
          7350 => x"fc",
          7351 => x"8f",
          7352 => x"f4",
          7353 => x"f4",
          7354 => x"0b",
          7355 => x"23",
          7356 => x"53",
          7357 => x"ff",
          7358 => x"c3",
          7359 => x"ba",
          7360 => x"7e",
          7361 => x"0b",
          7362 => x"84",
          7363 => x"59",
          7364 => x"34",
          7365 => x"1a",
          7366 => x"f4",
          7367 => x"86",
          7368 => x"0b",
          7369 => x"84",
          7370 => x"84",
          7371 => x"ff",
          7372 => x"80",
          7373 => x"ff",
          7374 => x"88",
          7375 => x"57",
          7376 => x"88",
          7377 => x"64",
          7378 => x"84",
          7379 => x"70",
          7380 => x"84",
          7381 => x"05",
          7382 => x"43",
          7383 => x"05",
          7384 => x"83",
          7385 => x"ee",
          7386 => x"24",
          7387 => x"61",
          7388 => x"06",
          7389 => x"27",
          7390 => x"fc",
          7391 => x"80",
          7392 => x"38",
          7393 => x"fb",
          7394 => x"73",
          7395 => x"0c",
          7396 => x"04",
          7397 => x"11",
          7398 => x"33",
          7399 => x"71",
          7400 => x"7a",
          7401 => x"33",
          7402 => x"71",
          7403 => x"83",
          7404 => x"05",
          7405 => x"85",
          7406 => x"88",
          7407 => x"88",
          7408 => x"45",
          7409 => x"58",
          7410 => x"56",
          7411 => x"05",
          7412 => x"85",
          7413 => x"ba",
          7414 => x"17",
          7415 => x"85",
          7416 => x"8b",
          7417 => x"2b",
          7418 => x"86",
          7419 => x"15",
          7420 => x"2b",
          7421 => x"2a",
          7422 => x"48",
          7423 => x"41",
          7424 => x"05",
          7425 => x"87",
          7426 => x"ba",
          7427 => x"70",
          7428 => x"33",
          7429 => x"07",
          7430 => x"06",
          7431 => x"5f",
          7432 => x"7b",
          7433 => x"81",
          7434 => x"ba",
          7435 => x"1f",
          7436 => x"83",
          7437 => x"8b",
          7438 => x"2b",
          7439 => x"73",
          7440 => x"33",
          7441 => x"07",
          7442 => x"5e",
          7443 => x"43",
          7444 => x"76",
          7445 => x"81",
          7446 => x"ba",
          7447 => x"1f",
          7448 => x"12",
          7449 => x"2b",
          7450 => x"07",
          7451 => x"14",
          7452 => x"33",
          7453 => x"07",
          7454 => x"40",
          7455 => x"40",
          7456 => x"78",
          7457 => x"60",
          7458 => x"84",
          7459 => x"70",
          7460 => x"33",
          7461 => x"71",
          7462 => x"66",
          7463 => x"70",
          7464 => x"52",
          7465 => x"05",
          7466 => x"fe",
          7467 => x"84",
          7468 => x"1e",
          7469 => x"83",
          7470 => x"5c",
          7471 => x"39",
          7472 => x"0b",
          7473 => x"0c",
          7474 => x"84",
          7475 => x"82",
          7476 => x"7f",
          7477 => x"f4",
          7478 => x"a5",
          7479 => x"f4",
          7480 => x"76",
          7481 => x"81",
          7482 => x"ba",
          7483 => x"7f",
          7484 => x"81",
          7485 => x"34",
          7486 => x"08",
          7487 => x"15",
          7488 => x"87",
          7489 => x"ba",
          7490 => x"ba",
          7491 => x"05",
          7492 => x"07",
          7493 => x"ff",
          7494 => x"2a",
          7495 => x"5e",
          7496 => x"34",
          7497 => x"34",
          7498 => x"22",
          7499 => x"10",
          7500 => x"08",
          7501 => x"5c",
          7502 => x"1c",
          7503 => x"83",
          7504 => x"51",
          7505 => x"7f",
          7506 => x"39",
          7507 => x"87",
          7508 => x"8b",
          7509 => x"2b",
          7510 => x"84",
          7511 => x"1d",
          7512 => x"2b",
          7513 => x"2a",
          7514 => x"43",
          7515 => x"61",
          7516 => x"63",
          7517 => x"34",
          7518 => x"08",
          7519 => x"11",
          7520 => x"33",
          7521 => x"71",
          7522 => x"74",
          7523 => x"33",
          7524 => x"71",
          7525 => x"70",
          7526 => x"5f",
          7527 => x"56",
          7528 => x"64",
          7529 => x"78",
          7530 => x"34",
          7531 => x"08",
          7532 => x"81",
          7533 => x"88",
          7534 => x"ff",
          7535 => x"88",
          7536 => x"58",
          7537 => x"34",
          7538 => x"34",
          7539 => x"08",
          7540 => x"33",
          7541 => x"71",
          7542 => x"83",
          7543 => x"05",
          7544 => x"12",
          7545 => x"2b",
          7546 => x"2b",
          7547 => x"06",
          7548 => x"88",
          7549 => x"5d",
          7550 => x"5d",
          7551 => x"82",
          7552 => x"83",
          7553 => x"ba",
          7554 => x"1f",
          7555 => x"12",
          7556 => x"2b",
          7557 => x"07",
          7558 => x"33",
          7559 => x"71",
          7560 => x"81",
          7561 => x"70",
          7562 => x"5d",
          7563 => x"5a",
          7564 => x"60",
          7565 => x"81",
          7566 => x"83",
          7567 => x"5b",
          7568 => x"86",
          7569 => x"16",
          7570 => x"2b",
          7571 => x"07",
          7572 => x"18",
          7573 => x"33",
          7574 => x"07",
          7575 => x"5e",
          7576 => x"41",
          7577 => x"1e",
          7578 => x"1e",
          7579 => x"f4",
          7580 => x"84",
          7581 => x"12",
          7582 => x"2b",
          7583 => x"07",
          7584 => x"14",
          7585 => x"33",
          7586 => x"07",
          7587 => x"44",
          7588 => x"5a",
          7589 => x"7c",
          7590 => x"34",
          7591 => x"05",
          7592 => x"f4",
          7593 => x"33",
          7594 => x"71",
          7595 => x"81",
          7596 => x"70",
          7597 => x"5b",
          7598 => x"75",
          7599 => x"16",
          7600 => x"f4",
          7601 => x"70",
          7602 => x"33",
          7603 => x"71",
          7604 => x"74",
          7605 => x"81",
          7606 => x"88",
          7607 => x"83",
          7608 => x"f8",
          7609 => x"63",
          7610 => x"54",
          7611 => x"59",
          7612 => x"7f",
          7613 => x"7b",
          7614 => x"84",
          7615 => x"70",
          7616 => x"81",
          7617 => x"8b",
          7618 => x"2b",
          7619 => x"70",
          7620 => x"33",
          7621 => x"07",
          7622 => x"06",
          7623 => x"5d",
          7624 => x"5b",
          7625 => x"75",
          7626 => x"81",
          7627 => x"ba",
          7628 => x"1f",
          7629 => x"83",
          7630 => x"8b",
          7631 => x"2b",
          7632 => x"86",
          7633 => x"12",
          7634 => x"2b",
          7635 => x"07",
          7636 => x"14",
          7637 => x"33",
          7638 => x"07",
          7639 => x"59",
          7640 => x"5c",
          7641 => x"5d",
          7642 => x"77",
          7643 => x"79",
          7644 => x"84",
          7645 => x"70",
          7646 => x"33",
          7647 => x"71",
          7648 => x"83",
          7649 => x"05",
          7650 => x"87",
          7651 => x"88",
          7652 => x"88",
          7653 => x"5e",
          7654 => x"41",
          7655 => x"16",
          7656 => x"16",
          7657 => x"f4",
          7658 => x"33",
          7659 => x"71",
          7660 => x"81",
          7661 => x"70",
          7662 => x"5c",
          7663 => x"79",
          7664 => x"1a",
          7665 => x"f4",
          7666 => x"82",
          7667 => x"12",
          7668 => x"2b",
          7669 => x"07",
          7670 => x"33",
          7671 => x"71",
          7672 => x"70",
          7673 => x"5c",
          7674 => x"5a",
          7675 => x"79",
          7676 => x"1a",
          7677 => x"f4",
          7678 => x"70",
          7679 => x"33",
          7680 => x"71",
          7681 => x"74",
          7682 => x"33",
          7683 => x"71",
          7684 => x"70",
          7685 => x"5c",
          7686 => x"5a",
          7687 => x"82",
          7688 => x"83",
          7689 => x"ba",
          7690 => x"1f",
          7691 => x"83",
          7692 => x"88",
          7693 => x"57",
          7694 => x"83",
          7695 => x"5a",
          7696 => x"84",
          7697 => x"b4",
          7698 => x"ba",
          7699 => x"84",
          7700 => x"05",
          7701 => x"ff",
          7702 => x"44",
          7703 => x"39",
          7704 => x"87",
          7705 => x"8b",
          7706 => x"2b",
          7707 => x"84",
          7708 => x"1d",
          7709 => x"2b",
          7710 => x"2a",
          7711 => x"43",
          7712 => x"61",
          7713 => x"63",
          7714 => x"34",
          7715 => x"08",
          7716 => x"11",
          7717 => x"33",
          7718 => x"71",
          7719 => x"74",
          7720 => x"33",
          7721 => x"71",
          7722 => x"70",
          7723 => x"41",
          7724 => x"59",
          7725 => x"64",
          7726 => x"7a",
          7727 => x"34",
          7728 => x"08",
          7729 => x"81",
          7730 => x"88",
          7731 => x"ff",
          7732 => x"88",
          7733 => x"42",
          7734 => x"34",
          7735 => x"34",
          7736 => x"08",
          7737 => x"33",
          7738 => x"71",
          7739 => x"83",
          7740 => x"05",
          7741 => x"12",
          7742 => x"2b",
          7743 => x"2b",
          7744 => x"06",
          7745 => x"88",
          7746 => x"5c",
          7747 => x"45",
          7748 => x"82",
          7749 => x"83",
          7750 => x"ba",
          7751 => x"1f",
          7752 => x"12",
          7753 => x"2b",
          7754 => x"07",
          7755 => x"33",
          7756 => x"71",
          7757 => x"81",
          7758 => x"70",
          7759 => x"5f",
          7760 => x"59",
          7761 => x"7d",
          7762 => x"1e",
          7763 => x"ff",
          7764 => x"f3",
          7765 => x"60",
          7766 => x"a1",
          7767 => x"84",
          7768 => x"bb",
          7769 => x"2e",
          7770 => x"53",
          7771 => x"bb",
          7772 => x"fe",
          7773 => x"73",
          7774 => x"3f",
          7775 => x"7b",
          7776 => x"38",
          7777 => x"f9",
          7778 => x"7a",
          7779 => x"f4",
          7780 => x"76",
          7781 => x"38",
          7782 => x"8a",
          7783 => x"bb",
          7784 => x"3d",
          7785 => x"51",
          7786 => x"84",
          7787 => x"54",
          7788 => x"08",
          7789 => x"38",
          7790 => x"52",
          7791 => x"08",
          7792 => x"bd",
          7793 => x"bb",
          7794 => x"3d",
          7795 => x"ff",
          7796 => x"ba",
          7797 => x"80",
          7798 => x"f0",
          7799 => x"80",
          7800 => x"84",
          7801 => x"fe",
          7802 => x"84",
          7803 => x"55",
          7804 => x"81",
          7805 => x"34",
          7806 => x"08",
          7807 => x"15",
          7808 => x"85",
          7809 => x"ba",
          7810 => x"76",
          7811 => x"81",
          7812 => x"34",
          7813 => x"08",
          7814 => x"22",
          7815 => x"80",
          7816 => x"83",
          7817 => x"70",
          7818 => x"51",
          7819 => x"88",
          7820 => x"89",
          7821 => x"ba",
          7822 => x"10",
          7823 => x"ba",
          7824 => x"f8",
          7825 => x"76",
          7826 => x"81",
          7827 => x"34",
          7828 => x"80",
          7829 => x"38",
          7830 => x"ff",
          7831 => x"8f",
          7832 => x"81",
          7833 => x"26",
          7834 => x"bb",
          7835 => x"52",
          7836 => x"84",
          7837 => x"0d",
          7838 => x"0d",
          7839 => x"33",
          7840 => x"71",
          7841 => x"38",
          7842 => x"bb",
          7843 => x"84",
          7844 => x"06",
          7845 => x"38",
          7846 => x"80",
          7847 => x"bb",
          7848 => x"53",
          7849 => x"84",
          7850 => x"0d",
          7851 => x"0d",
          7852 => x"02",
          7853 => x"05",
          7854 => x"57",
          7855 => x"76",
          7856 => x"38",
          7857 => x"17",
          7858 => x"81",
          7859 => x"55",
          7860 => x"73",
          7861 => x"87",
          7862 => x"0c",
          7863 => x"52",
          7864 => x"ca",
          7865 => x"84",
          7866 => x"06",
          7867 => x"2e",
          7868 => x"c0",
          7869 => x"54",
          7870 => x"79",
          7871 => x"38",
          7872 => x"80",
          7873 => x"80",
          7874 => x"81",
          7875 => x"74",
          7876 => x"0c",
          7877 => x"04",
          7878 => x"81",
          7879 => x"ff",
          7880 => x"56",
          7881 => x"ff",
          7882 => x"39",
          7883 => x"7c",
          7884 => x"8c",
          7885 => x"33",
          7886 => x"59",
          7887 => x"74",
          7888 => x"84",
          7889 => x"33",
          7890 => x"06",
          7891 => x"73",
          7892 => x"58",
          7893 => x"c0",
          7894 => x"78",
          7895 => x"76",
          7896 => x"3f",
          7897 => x"08",
          7898 => x"55",
          7899 => x"a7",
          7900 => x"98",
          7901 => x"73",
          7902 => x"78",
          7903 => x"74",
          7904 => x"06",
          7905 => x"2e",
          7906 => x"54",
          7907 => x"84",
          7908 => x"8b",
          7909 => x"84",
          7910 => x"19",
          7911 => x"06",
          7912 => x"79",
          7913 => x"ac",
          7914 => x"fc",
          7915 => x"02",
          7916 => x"05",
          7917 => x"05",
          7918 => x"53",
          7919 => x"53",
          7920 => x"87",
          7921 => x"80",
          7922 => x"72",
          7923 => x"83",
          7924 => x"38",
          7925 => x"c0",
          7926 => x"81",
          7927 => x"2e",
          7928 => x"71",
          7929 => x"70",
          7930 => x"38",
          7931 => x"84",
          7932 => x"86",
          7933 => x"88",
          7934 => x"0c",
          7935 => x"84",
          7936 => x"0d",
          7937 => x"75",
          7938 => x"84",
          7939 => x"86",
          7940 => x"71",
          7941 => x"c0",
          7942 => x"53",
          7943 => x"38",
          7944 => x"81",
          7945 => x"51",
          7946 => x"2e",
          7947 => x"c0",
          7948 => x"55",
          7949 => x"87",
          7950 => x"08",
          7951 => x"38",
          7952 => x"87",
          7953 => x"14",
          7954 => x"82",
          7955 => x"80",
          7956 => x"38",
          7957 => x"06",
          7958 => x"38",
          7959 => x"f6",
          7960 => x"58",
          7961 => x"19",
          7962 => x"56",
          7963 => x"2e",
          7964 => x"a8",
          7965 => x"56",
          7966 => x"81",
          7967 => x"53",
          7968 => x"18",
          7969 => x"a3",
          7970 => x"84",
          7971 => x"83",
          7972 => x"78",
          7973 => x"0c",
          7974 => x"04",
          7975 => x"18",
          7976 => x"18",
          7977 => x"19",
          7978 => x"fc",
          7979 => x"59",
          7980 => x"08",
          7981 => x"81",
          7982 => x"84",
          7983 => x"83",
          7984 => x"18",
          7985 => x"1a",
          7986 => x"1a",
          7987 => x"84",
          7988 => x"56",
          7989 => x"27",
          7990 => x"82",
          7991 => x"74",
          7992 => x"81",
          7993 => x"38",
          7994 => x"1b",
          7995 => x"81",
          7996 => x"fc",
          7997 => x"78",
          7998 => x"75",
          7999 => x"81",
          8000 => x"38",
          8001 => x"57",
          8002 => x"09",
          8003 => x"ee",
          8004 => x"5a",
          8005 => x"56",
          8006 => x"70",
          8007 => x"34",
          8008 => x"76",
          8009 => x"d5",
          8010 => x"19",
          8011 => x"0b",
          8012 => x"34",
          8013 => x"34",
          8014 => x"b9",
          8015 => x"e1",
          8016 => x"34",
          8017 => x"bb",
          8018 => x"f2",
          8019 => x"19",
          8020 => x"0b",
          8021 => x"34",
          8022 => x"84",
          8023 => x"80",
          8024 => x"9f",
          8025 => x"18",
          8026 => x"84",
          8027 => x"74",
          8028 => x"7a",
          8029 => x"34",
          8030 => x"56",
          8031 => x"19",
          8032 => x"2a",
          8033 => x"a3",
          8034 => x"18",
          8035 => x"84",
          8036 => x"7a",
          8037 => x"74",
          8038 => x"34",
          8039 => x"56",
          8040 => x"19",
          8041 => x"2a",
          8042 => x"a7",
          8043 => x"18",
          8044 => x"70",
          8045 => x"5b",
          8046 => x"53",
          8047 => x"18",
          8048 => x"e8",
          8049 => x"19",
          8050 => x"80",
          8051 => x"33",
          8052 => x"3f",
          8053 => x"08",
          8054 => x"b7",
          8055 => x"39",
          8056 => x"60",
          8057 => x"59",
          8058 => x"76",
          8059 => x"9c",
          8060 => x"26",
          8061 => x"58",
          8062 => x"84",
          8063 => x"0d",
          8064 => x"33",
          8065 => x"82",
          8066 => x"38",
          8067 => x"82",
          8068 => x"81",
          8069 => x"06",
          8070 => x"81",
          8071 => x"89",
          8072 => x"08",
          8073 => x"80",
          8074 => x"08",
          8075 => x"38",
          8076 => x"5c",
          8077 => x"09",
          8078 => x"de",
          8079 => x"78",
          8080 => x"52",
          8081 => x"51",
          8082 => x"84",
          8083 => x"80",
          8084 => x"ff",
          8085 => x"78",
          8086 => x"7a",
          8087 => x"79",
          8088 => x"17",
          8089 => x"81",
          8090 => x"2a",
          8091 => x"05",
          8092 => x"59",
          8093 => x"79",
          8094 => x"80",
          8095 => x"33",
          8096 => x"5d",
          8097 => x"09",
          8098 => x"b5",
          8099 => x"78",
          8100 => x"52",
          8101 => x"51",
          8102 => x"84",
          8103 => x"80",
          8104 => x"ff",
          8105 => x"78",
          8106 => x"79",
          8107 => x"7a",
          8108 => x"17",
          8109 => x"70",
          8110 => x"07",
          8111 => x"71",
          8112 => x"5d",
          8113 => x"79",
          8114 => x"76",
          8115 => x"84",
          8116 => x"8f",
          8117 => x"75",
          8118 => x"18",
          8119 => x"b4",
          8120 => x"2e",
          8121 => x"0b",
          8122 => x"71",
          8123 => x"7b",
          8124 => x"81",
          8125 => x"38",
          8126 => x"53",
          8127 => x"81",
          8128 => x"f7",
          8129 => x"bb",
          8130 => x"2e",
          8131 => x"59",
          8132 => x"b4",
          8133 => x"fd",
          8134 => x"10",
          8135 => x"77",
          8136 => x"81",
          8137 => x"33",
          8138 => x"07",
          8139 => x"0c",
          8140 => x"3d",
          8141 => x"83",
          8142 => x"06",
          8143 => x"75",
          8144 => x"18",
          8145 => x"b4",
          8146 => x"2e",
          8147 => x"0b",
          8148 => x"71",
          8149 => x"7c",
          8150 => x"81",
          8151 => x"38",
          8152 => x"53",
          8153 => x"81",
          8154 => x"f6",
          8155 => x"bb",
          8156 => x"2e",
          8157 => x"59",
          8158 => x"b4",
          8159 => x"fc",
          8160 => x"82",
          8161 => x"06",
          8162 => x"05",
          8163 => x"82",
          8164 => x"90",
          8165 => x"2b",
          8166 => x"33",
          8167 => x"88",
          8168 => x"71",
          8169 => x"fe",
          8170 => x"84",
          8171 => x"41",
          8172 => x"5a",
          8173 => x"0d",
          8174 => x"b4",
          8175 => x"b8",
          8176 => x"81",
          8177 => x"5c",
          8178 => x"81",
          8179 => x"84",
          8180 => x"09",
          8181 => x"be",
          8182 => x"84",
          8183 => x"34",
          8184 => x"a8",
          8185 => x"84",
          8186 => x"5b",
          8187 => x"18",
          8188 => x"84",
          8189 => x"33",
          8190 => x"2e",
          8191 => x"fd",
          8192 => x"54",
          8193 => x"a0",
          8194 => x"53",
          8195 => x"17",
          8196 => x"98",
          8197 => x"fd",
          8198 => x"54",
          8199 => x"53",
          8200 => x"53",
          8201 => x"52",
          8202 => x"3f",
          8203 => x"08",
          8204 => x"81",
          8205 => x"38",
          8206 => x"08",
          8207 => x"b4",
          8208 => x"18",
          8209 => x"7c",
          8210 => x"27",
          8211 => x"17",
          8212 => x"82",
          8213 => x"38",
          8214 => x"08",
          8215 => x"39",
          8216 => x"17",
          8217 => x"17",
          8218 => x"18",
          8219 => x"f5",
          8220 => x"5a",
          8221 => x"08",
          8222 => x"81",
          8223 => x"38",
          8224 => x"08",
          8225 => x"b4",
          8226 => x"18",
          8227 => x"bb",
          8228 => x"5e",
          8229 => x"08",
          8230 => x"38",
          8231 => x"55",
          8232 => x"09",
          8233 => x"b8",
          8234 => x"b4",
          8235 => x"18",
          8236 => x"7b",
          8237 => x"33",
          8238 => x"3f",
          8239 => x"a0",
          8240 => x"b4",
          8241 => x"b8",
          8242 => x"81",
          8243 => x"5e",
          8244 => x"81",
          8245 => x"84",
          8246 => x"09",
          8247 => x"cb",
          8248 => x"84",
          8249 => x"34",
          8250 => x"a8",
          8251 => x"84",
          8252 => x"5b",
          8253 => x"18",
          8254 => x"91",
          8255 => x"33",
          8256 => x"2e",
          8257 => x"fb",
          8258 => x"54",
          8259 => x"a0",
          8260 => x"53",
          8261 => x"17",
          8262 => x"90",
          8263 => x"fa",
          8264 => x"54",
          8265 => x"a0",
          8266 => x"53",
          8267 => x"17",
          8268 => x"f8",
          8269 => x"39",
          8270 => x"f9",
          8271 => x"9f",
          8272 => x"0d",
          8273 => x"5d",
          8274 => x"58",
          8275 => x"9c",
          8276 => x"1a",
          8277 => x"38",
          8278 => x"74",
          8279 => x"38",
          8280 => x"81",
          8281 => x"81",
          8282 => x"38",
          8283 => x"84",
          8284 => x"0d",
          8285 => x"2a",
          8286 => x"05",
          8287 => x"b4",
          8288 => x"5c",
          8289 => x"86",
          8290 => x"19",
          8291 => x"5d",
          8292 => x"09",
          8293 => x"fa",
          8294 => x"77",
          8295 => x"52",
          8296 => x"51",
          8297 => x"84",
          8298 => x"80",
          8299 => x"ff",
          8300 => x"77",
          8301 => x"79",
          8302 => x"b0",
          8303 => x"83",
          8304 => x"05",
          8305 => x"ff",
          8306 => x"76",
          8307 => x"76",
          8308 => x"79",
          8309 => x"81",
          8310 => x"34",
          8311 => x"84",
          8312 => x"0d",
          8313 => x"2e",
          8314 => x"fe",
          8315 => x"87",
          8316 => x"08",
          8317 => x"0b",
          8318 => x"58",
          8319 => x"2e",
          8320 => x"83",
          8321 => x"5b",
          8322 => x"2e",
          8323 => x"84",
          8324 => x"54",
          8325 => x"19",
          8326 => x"33",
          8327 => x"3f",
          8328 => x"08",
          8329 => x"38",
          8330 => x"5a",
          8331 => x"0c",
          8332 => x"fe",
          8333 => x"82",
          8334 => x"06",
          8335 => x"11",
          8336 => x"70",
          8337 => x"0a",
          8338 => x"0a",
          8339 => x"57",
          8340 => x"7d",
          8341 => x"2a",
          8342 => x"1d",
          8343 => x"2a",
          8344 => x"1d",
          8345 => x"2a",
          8346 => x"1d",
          8347 => x"83",
          8348 => x"e8",
          8349 => x"2a",
          8350 => x"2a",
          8351 => x"05",
          8352 => x"59",
          8353 => x"78",
          8354 => x"80",
          8355 => x"33",
          8356 => x"5d",
          8357 => x"09",
          8358 => x"d4",
          8359 => x"77",
          8360 => x"52",
          8361 => x"51",
          8362 => x"84",
          8363 => x"80",
          8364 => x"ff",
          8365 => x"77",
          8366 => x"7b",
          8367 => x"ac",
          8368 => x"ff",
          8369 => x"05",
          8370 => x"81",
          8371 => x"57",
          8372 => x"80",
          8373 => x"7a",
          8374 => x"f0",
          8375 => x"8f",
          8376 => x"56",
          8377 => x"34",
          8378 => x"1a",
          8379 => x"2a",
          8380 => x"05",
          8381 => x"b4",
          8382 => x"5f",
          8383 => x"83",
          8384 => x"54",
          8385 => x"19",
          8386 => x"1a",
          8387 => x"f0",
          8388 => x"58",
          8389 => x"08",
          8390 => x"81",
          8391 => x"38",
          8392 => x"08",
          8393 => x"b4",
          8394 => x"a8",
          8395 => x"a0",
          8396 => x"bb",
          8397 => x"5c",
          8398 => x"7a",
          8399 => x"82",
          8400 => x"74",
          8401 => x"e4",
          8402 => x"75",
          8403 => x"81",
          8404 => x"ee",
          8405 => x"bb",
          8406 => x"2e",
          8407 => x"56",
          8408 => x"b4",
          8409 => x"fc",
          8410 => x"83",
          8411 => x"b8",
          8412 => x"2a",
          8413 => x"8f",
          8414 => x"2a",
          8415 => x"f0",
          8416 => x"06",
          8417 => x"74",
          8418 => x"0b",
          8419 => x"fc",
          8420 => x"54",
          8421 => x"19",
          8422 => x"1a",
          8423 => x"ef",
          8424 => x"5a",
          8425 => x"08",
          8426 => x"81",
          8427 => x"38",
          8428 => x"08",
          8429 => x"b4",
          8430 => x"a8",
          8431 => x"a0",
          8432 => x"bb",
          8433 => x"59",
          8434 => x"77",
          8435 => x"38",
          8436 => x"55",
          8437 => x"09",
          8438 => x"bd",
          8439 => x"76",
          8440 => x"52",
          8441 => x"51",
          8442 => x"7b",
          8443 => x"39",
          8444 => x"53",
          8445 => x"53",
          8446 => x"52",
          8447 => x"3f",
          8448 => x"bb",
          8449 => x"2e",
          8450 => x"fd",
          8451 => x"bb",
          8452 => x"1a",
          8453 => x"08",
          8454 => x"08",
          8455 => x"08",
          8456 => x"08",
          8457 => x"5f",
          8458 => x"fc",
          8459 => x"19",
          8460 => x"82",
          8461 => x"06",
          8462 => x"81",
          8463 => x"53",
          8464 => x"19",
          8465 => x"e4",
          8466 => x"fc",
          8467 => x"54",
          8468 => x"19",
          8469 => x"1a",
          8470 => x"ed",
          8471 => x"5a",
          8472 => x"08",
          8473 => x"81",
          8474 => x"38",
          8475 => x"08",
          8476 => x"b4",
          8477 => x"a8",
          8478 => x"a0",
          8479 => x"bb",
          8480 => x"5f",
          8481 => x"7d",
          8482 => x"38",
          8483 => x"55",
          8484 => x"09",
          8485 => x"fa",
          8486 => x"7c",
          8487 => x"52",
          8488 => x"51",
          8489 => x"7b",
          8490 => x"39",
          8491 => x"1c",
          8492 => x"81",
          8493 => x"ec",
          8494 => x"58",
          8495 => x"7b",
          8496 => x"fe",
          8497 => x"7c",
          8498 => x"06",
          8499 => x"76",
          8500 => x"76",
          8501 => x"79",
          8502 => x"f9",
          8503 => x"58",
          8504 => x"7b",
          8505 => x"83",
          8506 => x"05",
          8507 => x"11",
          8508 => x"2b",
          8509 => x"7f",
          8510 => x"07",
          8511 => x"5d",
          8512 => x"34",
          8513 => x"56",
          8514 => x"34",
          8515 => x"5a",
          8516 => x"34",
          8517 => x"5b",
          8518 => x"34",
          8519 => x"f6",
          8520 => x"7e",
          8521 => x"5c",
          8522 => x"8a",
          8523 => x"08",
          8524 => x"2e",
          8525 => x"76",
          8526 => x"27",
          8527 => x"94",
          8528 => x"56",
          8529 => x"2e",
          8530 => x"76",
          8531 => x"93",
          8532 => x"81",
          8533 => x"19",
          8534 => x"89",
          8535 => x"75",
          8536 => x"b2",
          8537 => x"79",
          8538 => x"3f",
          8539 => x"08",
          8540 => x"d0",
          8541 => x"84",
          8542 => x"81",
          8543 => x"84",
          8544 => x"09",
          8545 => x"72",
          8546 => x"70",
          8547 => x"51",
          8548 => x"82",
          8549 => x"77",
          8550 => x"06",
          8551 => x"73",
          8552 => x"bb",
          8553 => x"3d",
          8554 => x"57",
          8555 => x"84",
          8556 => x"58",
          8557 => x"52",
          8558 => x"a4",
          8559 => x"74",
          8560 => x"08",
          8561 => x"84",
          8562 => x"55",
          8563 => x"08",
          8564 => x"38",
          8565 => x"84",
          8566 => x"26",
          8567 => x"57",
          8568 => x"81",
          8569 => x"19",
          8570 => x"83",
          8571 => x"75",
          8572 => x"ef",
          8573 => x"58",
          8574 => x"08",
          8575 => x"a0",
          8576 => x"84",
          8577 => x"30",
          8578 => x"80",
          8579 => x"07",
          8580 => x"08",
          8581 => x"55",
          8582 => x"85",
          8583 => x"84",
          8584 => x"9a",
          8585 => x"08",
          8586 => x"27",
          8587 => x"73",
          8588 => x"27",
          8589 => x"73",
          8590 => x"fe",
          8591 => x"80",
          8592 => x"38",
          8593 => x"52",
          8594 => x"f5",
          8595 => x"84",
          8596 => x"84",
          8597 => x"84",
          8598 => x"07",
          8599 => x"58",
          8600 => x"c4",
          8601 => x"e3",
          8602 => x"1a",
          8603 => x"08",
          8604 => x"1a",
          8605 => x"74",
          8606 => x"38",
          8607 => x"1a",
          8608 => x"33",
          8609 => x"79",
          8610 => x"75",
          8611 => x"bb",
          8612 => x"3d",
          8613 => x"0b",
          8614 => x"0c",
          8615 => x"04",
          8616 => x"08",
          8617 => x"39",
          8618 => x"ff",
          8619 => x"53",
          8620 => x"51",
          8621 => x"84",
          8622 => x"55",
          8623 => x"84",
          8624 => x"84",
          8625 => x"8c",
          8626 => x"ff",
          8627 => x"2e",
          8628 => x"81",
          8629 => x"39",
          8630 => x"7a",
          8631 => x"59",
          8632 => x"f0",
          8633 => x"80",
          8634 => x"9f",
          8635 => x"80",
          8636 => x"90",
          8637 => x"18",
          8638 => x"80",
          8639 => x"33",
          8640 => x"26",
          8641 => x"73",
          8642 => x"82",
          8643 => x"22",
          8644 => x"79",
          8645 => x"ac",
          8646 => x"19",
          8647 => x"19",
          8648 => x"08",
          8649 => x"72",
          8650 => x"38",
          8651 => x"13",
          8652 => x"73",
          8653 => x"17",
          8654 => x"19",
          8655 => x"75",
          8656 => x"0c",
          8657 => x"04",
          8658 => x"bb",
          8659 => x"3d",
          8660 => x"17",
          8661 => x"80",
          8662 => x"38",
          8663 => x"70",
          8664 => x"59",
          8665 => x"a5",
          8666 => x"08",
          8667 => x"fe",
          8668 => x"80",
          8669 => x"27",
          8670 => x"17",
          8671 => x"29",
          8672 => x"05",
          8673 => x"98",
          8674 => x"91",
          8675 => x"77",
          8676 => x"3f",
          8677 => x"08",
          8678 => x"84",
          8679 => x"a4",
          8680 => x"84",
          8681 => x"27",
          8682 => x"9c",
          8683 => x"84",
          8684 => x"73",
          8685 => x"38",
          8686 => x"54",
          8687 => x"cd",
          8688 => x"39",
          8689 => x"bb",
          8690 => x"3d",
          8691 => x"3d",
          8692 => x"08",
          8693 => x"a0",
          8694 => x"57",
          8695 => x"7a",
          8696 => x"80",
          8697 => x"0c",
          8698 => x"55",
          8699 => x"80",
          8700 => x"79",
          8701 => x"5b",
          8702 => x"81",
          8703 => x"08",
          8704 => x"a9",
          8705 => x"2a",
          8706 => x"57",
          8707 => x"27",
          8708 => x"77",
          8709 => x"79",
          8710 => x"78",
          8711 => x"9c",
          8712 => x"56",
          8713 => x"84",
          8714 => x"0d",
          8715 => x"18",
          8716 => x"22",
          8717 => x"89",
          8718 => x"7b",
          8719 => x"52",
          8720 => x"9c",
          8721 => x"84",
          8722 => x"56",
          8723 => x"bb",
          8724 => x"d0",
          8725 => x"84",
          8726 => x"ff",
          8727 => x"9c",
          8728 => x"bb",
          8729 => x"82",
          8730 => x"80",
          8731 => x"38",
          8732 => x"52",
          8733 => x"a7",
          8734 => x"84",
          8735 => x"56",
          8736 => x"08",
          8737 => x"9c",
          8738 => x"84",
          8739 => x"81",
          8740 => x"38",
          8741 => x"bb",
          8742 => x"2e",
          8743 => x"84",
          8744 => x"83",
          8745 => x"58",
          8746 => x"38",
          8747 => x"1a",
          8748 => x"59",
          8749 => x"75",
          8750 => x"38",
          8751 => x"76",
          8752 => x"1b",
          8753 => x"5e",
          8754 => x"0c",
          8755 => x"84",
          8756 => x"55",
          8757 => x"81",
          8758 => x"ff",
          8759 => x"f4",
          8760 => x"8a",
          8761 => x"75",
          8762 => x"80",
          8763 => x"75",
          8764 => x"52",
          8765 => x"51",
          8766 => x"84",
          8767 => x"80",
          8768 => x"16",
          8769 => x"7a",
          8770 => x"84",
          8771 => x"84",
          8772 => x"0d",
          8773 => x"b4",
          8774 => x"b8",
          8775 => x"81",
          8776 => x"56",
          8777 => x"84",
          8778 => x"80",
          8779 => x"bb",
          8780 => x"1a",
          8781 => x"08",
          8782 => x"31",
          8783 => x"1a",
          8784 => x"e8",
          8785 => x"33",
          8786 => x"2e",
          8787 => x"fe",
          8788 => x"54",
          8789 => x"a0",
          8790 => x"53",
          8791 => x"19",
          8792 => x"c8",
          8793 => x"39",
          8794 => x"55",
          8795 => x"ff",
          8796 => x"76",
          8797 => x"06",
          8798 => x"94",
          8799 => x"1d",
          8800 => x"fe",
          8801 => x"80",
          8802 => x"27",
          8803 => x"8a",
          8804 => x"71",
          8805 => x"08",
          8806 => x"0c",
          8807 => x"39",
          8808 => x"bb",
          8809 => x"3d",
          8810 => x"3d",
          8811 => x"41",
          8812 => x"08",
          8813 => x"ff",
          8814 => x"08",
          8815 => x"75",
          8816 => x"d2",
          8817 => x"5f",
          8818 => x"58",
          8819 => x"76",
          8820 => x"38",
          8821 => x"78",
          8822 => x"78",
          8823 => x"06",
          8824 => x"81",
          8825 => x"b8",
          8826 => x"19",
          8827 => x"bd",
          8828 => x"84",
          8829 => x"85",
          8830 => x"81",
          8831 => x"1a",
          8832 => x"76",
          8833 => x"9c",
          8834 => x"33",
          8835 => x"80",
          8836 => x"38",
          8837 => x"bf",
          8838 => x"ff",
          8839 => x"60",
          8840 => x"76",
          8841 => x"70",
          8842 => x"32",
          8843 => x"80",
          8844 => x"25",
          8845 => x"45",
          8846 => x"93",
          8847 => x"df",
          8848 => x"61",
          8849 => x"bf",
          8850 => x"2e",
          8851 => x"81",
          8852 => x"52",
          8853 => x"f6",
          8854 => x"84",
          8855 => x"bb",
          8856 => x"b2",
          8857 => x"08",
          8858 => x"dc",
          8859 => x"bb",
          8860 => x"3d",
          8861 => x"54",
          8862 => x"53",
          8863 => x"19",
          8864 => x"a8",
          8865 => x"84",
          8866 => x"78",
          8867 => x"06",
          8868 => x"84",
          8869 => x"83",
          8870 => x"19",
          8871 => x"08",
          8872 => x"84",
          8873 => x"7a",
          8874 => x"27",
          8875 => x"82",
          8876 => x"60",
          8877 => x"81",
          8878 => x"38",
          8879 => x"19",
          8880 => x"08",
          8881 => x"52",
          8882 => x"51",
          8883 => x"77",
          8884 => x"39",
          8885 => x"09",
          8886 => x"e7",
          8887 => x"2a",
          8888 => x"7a",
          8889 => x"38",
          8890 => x"77",
          8891 => x"70",
          8892 => x"7f",
          8893 => x"59",
          8894 => x"7d",
          8895 => x"81",
          8896 => x"5d",
          8897 => x"81",
          8898 => x"2e",
          8899 => x"fe",
          8900 => x"39",
          8901 => x"0b",
          8902 => x"7a",
          8903 => x"0c",
          8904 => x"04",
          8905 => x"df",
          8906 => x"33",
          8907 => x"2e",
          8908 => x"cb",
          8909 => x"08",
          8910 => x"9a",
          8911 => x"88",
          8912 => x"56",
          8913 => x"b7",
          8914 => x"70",
          8915 => x"8d",
          8916 => x"51",
          8917 => x"58",
          8918 => x"84",
          8919 => x"05",
          8920 => x"71",
          8921 => x"2b",
          8922 => x"56",
          8923 => x"80",
          8924 => x"81",
          8925 => x"87",
          8926 => x"61",
          8927 => x"42",
          8928 => x"81",
          8929 => x"17",
          8930 => x"27",
          8931 => x"33",
          8932 => x"81",
          8933 => x"77",
          8934 => x"38",
          8935 => x"26",
          8936 => x"79",
          8937 => x"43",
          8938 => x"ff",
          8939 => x"ff",
          8940 => x"fd",
          8941 => x"83",
          8942 => x"ca",
          8943 => x"55",
          8944 => x"7c",
          8945 => x"55",
          8946 => x"81",
          8947 => x"80",
          8948 => x"70",
          8949 => x"33",
          8950 => x"70",
          8951 => x"ff",
          8952 => x"59",
          8953 => x"74",
          8954 => x"81",
          8955 => x"ac",
          8956 => x"84",
          8957 => x"94",
          8958 => x"ef",
          8959 => x"70",
          8960 => x"80",
          8961 => x"f5",
          8962 => x"bb",
          8963 => x"84",
          8964 => x"82",
          8965 => x"ff",
          8966 => x"ff",
          8967 => x"0c",
          8968 => x"98",
          8969 => x"80",
          8970 => x"08",
          8971 => x"cc",
          8972 => x"33",
          8973 => x"74",
          8974 => x"81",
          8975 => x"38",
          8976 => x"53",
          8977 => x"81",
          8978 => x"dc",
          8979 => x"bb",
          8980 => x"2e",
          8981 => x"56",
          8982 => x"b4",
          8983 => x"5a",
          8984 => x"38",
          8985 => x"70",
          8986 => x"76",
          8987 => x"99",
          8988 => x"33",
          8989 => x"81",
          8990 => x"58",
          8991 => x"34",
          8992 => x"2e",
          8993 => x"75",
          8994 => x"06",
          8995 => x"2e",
          8996 => x"74",
          8997 => x"75",
          8998 => x"e5",
          8999 => x"38",
          9000 => x"58",
          9001 => x"81",
          9002 => x"80",
          9003 => x"70",
          9004 => x"33",
          9005 => x"70",
          9006 => x"ff",
          9007 => x"5d",
          9008 => x"74",
          9009 => x"cd",
          9010 => x"33",
          9011 => x"76",
          9012 => x"0b",
          9013 => x"57",
          9014 => x"05",
          9015 => x"70",
          9016 => x"33",
          9017 => x"ff",
          9018 => x"42",
          9019 => x"2e",
          9020 => x"75",
          9021 => x"38",
          9022 => x"ff",
          9023 => x"0c",
          9024 => x"51",
          9025 => x"84",
          9026 => x"5a",
          9027 => x"08",
          9028 => x"8f",
          9029 => x"bb",
          9030 => x"3d",
          9031 => x"54",
          9032 => x"53",
          9033 => x"1b",
          9034 => x"80",
          9035 => x"84",
          9036 => x"78",
          9037 => x"06",
          9038 => x"84",
          9039 => x"83",
          9040 => x"1b",
          9041 => x"08",
          9042 => x"84",
          9043 => x"78",
          9044 => x"27",
          9045 => x"82",
          9046 => x"79",
          9047 => x"81",
          9048 => x"38",
          9049 => x"1b",
          9050 => x"08",
          9051 => x"52",
          9052 => x"51",
          9053 => x"77",
          9054 => x"39",
          9055 => x"e4",
          9056 => x"33",
          9057 => x"81",
          9058 => x"60",
          9059 => x"76",
          9060 => x"06",
          9061 => x"2e",
          9062 => x"19",
          9063 => x"bf",
          9064 => x"1f",
          9065 => x"05",
          9066 => x"5f",
          9067 => x"af",
          9068 => x"55",
          9069 => x"52",
          9070 => x"92",
          9071 => x"84",
          9072 => x"bb",
          9073 => x"2e",
          9074 => x"fe",
          9075 => x"80",
          9076 => x"38",
          9077 => x"ff",
          9078 => x"0c",
          9079 => x"8d",
          9080 => x"7e",
          9081 => x"81",
          9082 => x"8c",
          9083 => x"1a",
          9084 => x"33",
          9085 => x"07",
          9086 => x"76",
          9087 => x"78",
          9088 => x"06",
          9089 => x"05",
          9090 => x"77",
          9091 => x"e7",
          9092 => x"79",
          9093 => x"33",
          9094 => x"88",
          9095 => x"42",
          9096 => x"2e",
          9097 => x"79",
          9098 => x"ff",
          9099 => x"51",
          9100 => x"3f",
          9101 => x"08",
          9102 => x"05",
          9103 => x"43",
          9104 => x"56",
          9105 => x"3f",
          9106 => x"84",
          9107 => x"81",
          9108 => x"38",
          9109 => x"18",
          9110 => x"27",
          9111 => x"78",
          9112 => x"2a",
          9113 => x"59",
          9114 => x"92",
          9115 => x"2e",
          9116 => x"10",
          9117 => x"22",
          9118 => x"fe",
          9119 => x"1d",
          9120 => x"06",
          9121 => x"ae",
          9122 => x"84",
          9123 => x"93",
          9124 => x"76",
          9125 => x"2e",
          9126 => x"81",
          9127 => x"94",
          9128 => x"0d",
          9129 => x"70",
          9130 => x"81",
          9131 => x"5a",
          9132 => x"56",
          9133 => x"38",
          9134 => x"08",
          9135 => x"57",
          9136 => x"2e",
          9137 => x"1d",
          9138 => x"70",
          9139 => x"5d",
          9140 => x"95",
          9141 => x"5b",
          9142 => x"7b",
          9143 => x"75",
          9144 => x"57",
          9145 => x"81",
          9146 => x"ff",
          9147 => x"ef",
          9148 => x"db",
          9149 => x"81",
          9150 => x"76",
          9151 => x"aa",
          9152 => x"0b",
          9153 => x"81",
          9154 => x"40",
          9155 => x"08",
          9156 => x"8b",
          9157 => x"57",
          9158 => x"81",
          9159 => x"76",
          9160 => x"58",
          9161 => x"55",
          9162 => x"85",
          9163 => x"c2",
          9164 => x"22",
          9165 => x"80",
          9166 => x"74",
          9167 => x"56",
          9168 => x"81",
          9169 => x"07",
          9170 => x"70",
          9171 => x"06",
          9172 => x"81",
          9173 => x"56",
          9174 => x"2e",
          9175 => x"84",
          9176 => x"57",
          9177 => x"77",
          9178 => x"38",
          9179 => x"74",
          9180 => x"02",
          9181 => x"cf",
          9182 => x"76",
          9183 => x"06",
          9184 => x"27",
          9185 => x"15",
          9186 => x"34",
          9187 => x"19",
          9188 => x"59",
          9189 => x"e3",
          9190 => x"59",
          9191 => x"34",
          9192 => x"56",
          9193 => x"a0",
          9194 => x"55",
          9195 => x"98",
          9196 => x"56",
          9197 => x"88",
          9198 => x"1a",
          9199 => x"57",
          9200 => x"09",
          9201 => x"38",
          9202 => x"a0",
          9203 => x"26",
          9204 => x"3d",
          9205 => x"05",
          9206 => x"33",
          9207 => x"74",
          9208 => x"76",
          9209 => x"38",
          9210 => x"8f",
          9211 => x"84",
          9212 => x"81",
          9213 => x"e3",
          9214 => x"91",
          9215 => x"7a",
          9216 => x"82",
          9217 => x"bb",
          9218 => x"84",
          9219 => x"84",
          9220 => x"06",
          9221 => x"02",
          9222 => x"33",
          9223 => x"7d",
          9224 => x"05",
          9225 => x"33",
          9226 => x"81",
          9227 => x"5f",
          9228 => x"80",
          9229 => x"8d",
          9230 => x"51",
          9231 => x"3f",
          9232 => x"08",
          9233 => x"52",
          9234 => x"8c",
          9235 => x"84",
          9236 => x"bb",
          9237 => x"82",
          9238 => x"84",
          9239 => x"5e",
          9240 => x"08",
          9241 => x"b4",
          9242 => x"2e",
          9243 => x"83",
          9244 => x"7f",
          9245 => x"81",
          9246 => x"38",
          9247 => x"53",
          9248 => x"81",
          9249 => x"d4",
          9250 => x"bb",
          9251 => x"2e",
          9252 => x"56",
          9253 => x"b4",
          9254 => x"56",
          9255 => x"9c",
          9256 => x"33",
          9257 => x"81",
          9258 => x"c9",
          9259 => x"70",
          9260 => x"07",
          9261 => x"80",
          9262 => x"38",
          9263 => x"78",
          9264 => x"89",
          9265 => x"7d",
          9266 => x"3f",
          9267 => x"08",
          9268 => x"84",
          9269 => x"ff",
          9270 => x"58",
          9271 => x"81",
          9272 => x"58",
          9273 => x"38",
          9274 => x"7f",
          9275 => x"98",
          9276 => x"b4",
          9277 => x"2e",
          9278 => x"1c",
          9279 => x"40",
          9280 => x"38",
          9281 => x"53",
          9282 => x"81",
          9283 => x"d3",
          9284 => x"bb",
          9285 => x"2e",
          9286 => x"57",
          9287 => x"b4",
          9288 => x"58",
          9289 => x"38",
          9290 => x"1f",
          9291 => x"80",
          9292 => x"05",
          9293 => x"15",
          9294 => x"38",
          9295 => x"1f",
          9296 => x"58",
          9297 => x"81",
          9298 => x"77",
          9299 => x"59",
          9300 => x"55",
          9301 => x"9c",
          9302 => x"1f",
          9303 => x"5e",
          9304 => x"1b",
          9305 => x"83",
          9306 => x"56",
          9307 => x"84",
          9308 => x"0d",
          9309 => x"30",
          9310 => x"72",
          9311 => x"57",
          9312 => x"38",
          9313 => x"52",
          9314 => x"c2",
          9315 => x"84",
          9316 => x"bb",
          9317 => x"2e",
          9318 => x"fe",
          9319 => x"54",
          9320 => x"53",
          9321 => x"18",
          9322 => x"80",
          9323 => x"84",
          9324 => x"09",
          9325 => x"bf",
          9326 => x"84",
          9327 => x"34",
          9328 => x"a8",
          9329 => x"55",
          9330 => x"08",
          9331 => x"82",
          9332 => x"60",
          9333 => x"ac",
          9334 => x"84",
          9335 => x"9c",
          9336 => x"2b",
          9337 => x"71",
          9338 => x"7d",
          9339 => x"3f",
          9340 => x"08",
          9341 => x"84",
          9342 => x"38",
          9343 => x"84",
          9344 => x"8b",
          9345 => x"2a",
          9346 => x"29",
          9347 => x"81",
          9348 => x"57",
          9349 => x"81",
          9350 => x"19",
          9351 => x"76",
          9352 => x"81",
          9353 => x"1d",
          9354 => x"1e",
          9355 => x"56",
          9356 => x"77",
          9357 => x"83",
          9358 => x"7a",
          9359 => x"81",
          9360 => x"38",
          9361 => x"53",
          9362 => x"81",
          9363 => x"d0",
          9364 => x"bb",
          9365 => x"2e",
          9366 => x"57",
          9367 => x"b4",
          9368 => x"58",
          9369 => x"38",
          9370 => x"9c",
          9371 => x"81",
          9372 => x"5c",
          9373 => x"1c",
          9374 => x"8b",
          9375 => x"8c",
          9376 => x"9a",
          9377 => x"9b",
          9378 => x"8d",
          9379 => x"76",
          9380 => x"59",
          9381 => x"ff",
          9382 => x"78",
          9383 => x"22",
          9384 => x"58",
          9385 => x"84",
          9386 => x"05",
          9387 => x"70",
          9388 => x"34",
          9389 => x"56",
          9390 => x"76",
          9391 => x"ff",
          9392 => x"18",
          9393 => x"27",
          9394 => x"83",
          9395 => x"81",
          9396 => x"10",
          9397 => x"58",
          9398 => x"2e",
          9399 => x"7c",
          9400 => x"0b",
          9401 => x"80",
          9402 => x"e9",
          9403 => x"bb",
          9404 => x"84",
          9405 => x"fc",
          9406 => x"ff",
          9407 => x"fe",
          9408 => x"eb",
          9409 => x"b4",
          9410 => x"b8",
          9411 => x"81",
          9412 => x"59",
          9413 => x"81",
          9414 => x"84",
          9415 => x"38",
          9416 => x"08",
          9417 => x"b4",
          9418 => x"1d",
          9419 => x"bb",
          9420 => x"41",
          9421 => x"08",
          9422 => x"38",
          9423 => x"42",
          9424 => x"09",
          9425 => x"bc",
          9426 => x"b4",
          9427 => x"1d",
          9428 => x"78",
          9429 => x"33",
          9430 => x"3f",
          9431 => x"a4",
          9432 => x"1f",
          9433 => x"57",
          9434 => x"81",
          9435 => x"81",
          9436 => x"38",
          9437 => x"81",
          9438 => x"76",
          9439 => x"9f",
          9440 => x"39",
          9441 => x"07",
          9442 => x"39",
          9443 => x"1c",
          9444 => x"52",
          9445 => x"51",
          9446 => x"84",
          9447 => x"76",
          9448 => x"06",
          9449 => x"bb",
          9450 => x"1d",
          9451 => x"08",
          9452 => x"31",
          9453 => x"1d",
          9454 => x"38",
          9455 => x"5f",
          9456 => x"aa",
          9457 => x"84",
          9458 => x"f8",
          9459 => x"1c",
          9460 => x"80",
          9461 => x"38",
          9462 => x"75",
          9463 => x"e8",
          9464 => x"59",
          9465 => x"2e",
          9466 => x"fa",
          9467 => x"54",
          9468 => x"a0",
          9469 => x"53",
          9470 => x"1c",
          9471 => x"ac",
          9472 => x"39",
          9473 => x"18",
          9474 => x"08",
          9475 => x"52",
          9476 => x"51",
          9477 => x"f8",
          9478 => x"3d",
          9479 => x"71",
          9480 => x"5c",
          9481 => x"1e",
          9482 => x"08",
          9483 => x"b5",
          9484 => x"08",
          9485 => x"d9",
          9486 => x"71",
          9487 => x"08",
          9488 => x"58",
          9489 => x"72",
          9490 => x"38",
          9491 => x"14",
          9492 => x"1b",
          9493 => x"7a",
          9494 => x"80",
          9495 => x"70",
          9496 => x"06",
          9497 => x"8f",
          9498 => x"83",
          9499 => x"1a",
          9500 => x"22",
          9501 => x"5b",
          9502 => x"7a",
          9503 => x"25",
          9504 => x"06",
          9505 => x"7c",
          9506 => x"57",
          9507 => x"18",
          9508 => x"89",
          9509 => x"58",
          9510 => x"16",
          9511 => x"18",
          9512 => x"74",
          9513 => x"38",
          9514 => x"81",
          9515 => x"89",
          9516 => x"70",
          9517 => x"25",
          9518 => x"77",
          9519 => x"38",
          9520 => x"8b",
          9521 => x"70",
          9522 => x"34",
          9523 => x"74",
          9524 => x"05",
          9525 => x"18",
          9526 => x"27",
          9527 => x"7c",
          9528 => x"55",
          9529 => x"16",
          9530 => x"33",
          9531 => x"38",
          9532 => x"38",
          9533 => x"1e",
          9534 => x"7c",
          9535 => x"56",
          9536 => x"17",
          9537 => x"08",
          9538 => x"55",
          9539 => x"38",
          9540 => x"34",
          9541 => x"53",
          9542 => x"88",
          9543 => x"1c",
          9544 => x"83",
          9545 => x"12",
          9546 => x"2b",
          9547 => x"07",
          9548 => x"70",
          9549 => x"2b",
          9550 => x"07",
          9551 => x"97",
          9552 => x"17",
          9553 => x"2b",
          9554 => x"5b",
          9555 => x"5b",
          9556 => x"1e",
          9557 => x"33",
          9558 => x"71",
          9559 => x"5d",
          9560 => x"1e",
          9561 => x"0d",
          9562 => x"55",
          9563 => x"77",
          9564 => x"81",
          9565 => x"58",
          9566 => x"b5",
          9567 => x"2b",
          9568 => x"81",
          9569 => x"84",
          9570 => x"83",
          9571 => x"55",
          9572 => x"27",
          9573 => x"76",
          9574 => x"38",
          9575 => x"54",
          9576 => x"74",
          9577 => x"82",
          9578 => x"80",
          9579 => x"08",
          9580 => x"19",
          9581 => x"22",
          9582 => x"79",
          9583 => x"fd",
          9584 => x"30",
          9585 => x"78",
          9586 => x"72",
          9587 => x"58",
          9588 => x"80",
          9589 => x"7a",
          9590 => x"05",
          9591 => x"8c",
          9592 => x"5b",
          9593 => x"73",
          9594 => x"5a",
          9595 => x"80",
          9596 => x"38",
          9597 => x"7e",
          9598 => x"89",
          9599 => x"bf",
          9600 => x"78",
          9601 => x"38",
          9602 => x"8c",
          9603 => x"5b",
          9604 => x"b4",
          9605 => x"2a",
          9606 => x"06",
          9607 => x"2e",
          9608 => x"14",
          9609 => x"ff",
          9610 => x"73",
          9611 => x"05",
          9612 => x"16",
          9613 => x"19",
          9614 => x"33",
          9615 => x"56",
          9616 => x"b7",
          9617 => x"39",
          9618 => x"53",
          9619 => x"7b",
          9620 => x"25",
          9621 => x"06",
          9622 => x"58",
          9623 => x"ef",
          9624 => x"70",
          9625 => x"57",
          9626 => x"70",
          9627 => x"53",
          9628 => x"83",
          9629 => x"74",
          9630 => x"81",
          9631 => x"80",
          9632 => x"38",
          9633 => x"88",
          9634 => x"33",
          9635 => x"3d",
          9636 => x"9f",
          9637 => x"a7",
          9638 => x"8c",
          9639 => x"80",
          9640 => x"70",
          9641 => x"33",
          9642 => x"81",
          9643 => x"7f",
          9644 => x"2e",
          9645 => x"83",
          9646 => x"27",
          9647 => x"10",
          9648 => x"76",
          9649 => x"57",
          9650 => x"ff",
          9651 => x"32",
          9652 => x"73",
          9653 => x"25",
          9654 => x"5b",
          9655 => x"90",
          9656 => x"dc",
          9657 => x"38",
          9658 => x"26",
          9659 => x"e6",
          9660 => x"e6",
          9661 => x"81",
          9662 => x"54",
          9663 => x"2e",
          9664 => x"73",
          9665 => x"38",
          9666 => x"33",
          9667 => x"06",
          9668 => x"73",
          9669 => x"81",
          9670 => x"7a",
          9671 => x"76",
          9672 => x"80",
          9673 => x"10",
          9674 => x"7d",
          9675 => x"62",
          9676 => x"05",
          9677 => x"54",
          9678 => x"2e",
          9679 => x"80",
          9680 => x"73",
          9681 => x"70",
          9682 => x"25",
          9683 => x"55",
          9684 => x"80",
          9685 => x"81",
          9686 => x"54",
          9687 => x"54",
          9688 => x"2e",
          9689 => x"80",
          9690 => x"30",
          9691 => x"77",
          9692 => x"57",
          9693 => x"72",
          9694 => x"73",
          9695 => x"94",
          9696 => x"55",
          9697 => x"fe",
          9698 => x"39",
          9699 => x"73",
          9700 => x"ae",
          9701 => x"84",
          9702 => x"ff",
          9703 => x"fe",
          9704 => x"54",
          9705 => x"84",
          9706 => x"0d",
          9707 => x"a0",
          9708 => x"ff",
          9709 => x"7a",
          9710 => x"e3",
          9711 => x"ff",
          9712 => x"1d",
          9713 => x"7b",
          9714 => x"3f",
          9715 => x"08",
          9716 => x"0c",
          9717 => x"04",
          9718 => x"dc",
          9719 => x"70",
          9720 => x"07",
          9721 => x"56",
          9722 => x"a1",
          9723 => x"42",
          9724 => x"33",
          9725 => x"72",
          9726 => x"38",
          9727 => x"32",
          9728 => x"80",
          9729 => x"40",
          9730 => x"e1",
          9731 => x"0c",
          9732 => x"82",
          9733 => x"81",
          9734 => x"38",
          9735 => x"83",
          9736 => x"17",
          9737 => x"2e",
          9738 => x"17",
          9739 => x"05",
          9740 => x"a0",
          9741 => x"70",
          9742 => x"42",
          9743 => x"59",
          9744 => x"84",
          9745 => x"38",
          9746 => x"76",
          9747 => x"59",
          9748 => x"80",
          9749 => x"80",
          9750 => x"38",
          9751 => x"70",
          9752 => x"06",
          9753 => x"55",
          9754 => x"2e",
          9755 => x"73",
          9756 => x"06",
          9757 => x"2e",
          9758 => x"76",
          9759 => x"38",
          9760 => x"05",
          9761 => x"54",
          9762 => x"9d",
          9763 => x"18",
          9764 => x"ff",
          9765 => x"80",
          9766 => x"fe",
          9767 => x"5e",
          9768 => x"2e",
          9769 => x"eb",
          9770 => x"a0",
          9771 => x"a0",
          9772 => x"05",
          9773 => x"13",
          9774 => x"38",
          9775 => x"5e",
          9776 => x"70",
          9777 => x"59",
          9778 => x"74",
          9779 => x"ed",
          9780 => x"2e",
          9781 => x"74",
          9782 => x"30",
          9783 => x"55",
          9784 => x"77",
          9785 => x"38",
          9786 => x"38",
          9787 => x"7b",
          9788 => x"81",
          9789 => x"32",
          9790 => x"72",
          9791 => x"70",
          9792 => x"51",
          9793 => x"80",
          9794 => x"38",
          9795 => x"86",
          9796 => x"77",
          9797 => x"79",
          9798 => x"75",
          9799 => x"38",
          9800 => x"5b",
          9801 => x"2b",
          9802 => x"77",
          9803 => x"5d",
          9804 => x"22",
          9805 => x"56",
          9806 => x"95",
          9807 => x"33",
          9808 => x"e5",
          9809 => x"38",
          9810 => x"82",
          9811 => x"8c",
          9812 => x"8c",
          9813 => x"38",
          9814 => x"55",
          9815 => x"82",
          9816 => x"81",
          9817 => x"56",
          9818 => x"7d",
          9819 => x"7c",
          9820 => x"38",
          9821 => x"5a",
          9822 => x"81",
          9823 => x"80",
          9824 => x"79",
          9825 => x"79",
          9826 => x"7b",
          9827 => x"3f",
          9828 => x"08",
          9829 => x"56",
          9830 => x"84",
          9831 => x"81",
          9832 => x"bb",
          9833 => x"2e",
          9834 => x"fb",
          9835 => x"85",
          9836 => x"5a",
          9837 => x"84",
          9838 => x"82",
          9839 => x"59",
          9840 => x"38",
          9841 => x"55",
          9842 => x"8c",
          9843 => x"80",
          9844 => x"39",
          9845 => x"11",
          9846 => x"22",
          9847 => x"56",
          9848 => x"f0",
          9849 => x"2e",
          9850 => x"79",
          9851 => x"fd",
          9852 => x"18",
          9853 => x"ae",
          9854 => x"06",
          9855 => x"77",
          9856 => x"ae",
          9857 => x"06",
          9858 => x"76",
          9859 => x"80",
          9860 => x"0b",
          9861 => x"53",
          9862 => x"73",
          9863 => x"a0",
          9864 => x"70",
          9865 => x"34",
          9866 => x"8a",
          9867 => x"38",
          9868 => x"58",
          9869 => x"34",
          9870 => x"bf",
          9871 => x"84",
          9872 => x"33",
          9873 => x"bb",
          9874 => x"d6",
          9875 => x"2a",
          9876 => x"77",
          9877 => x"86",
          9878 => x"84",
          9879 => x"56",
          9880 => x"2e",
          9881 => x"90",
          9882 => x"ff",
          9883 => x"80",
          9884 => x"80",
          9885 => x"71",
          9886 => x"62",
          9887 => x"54",
          9888 => x"2e",
          9889 => x"74",
          9890 => x"7b",
          9891 => x"56",
          9892 => x"77",
          9893 => x"ae",
          9894 => x"38",
          9895 => x"76",
          9896 => x"fb",
          9897 => x"83",
          9898 => x"56",
          9899 => x"39",
          9900 => x"81",
          9901 => x"8c",
          9902 => x"77",
          9903 => x"81",
          9904 => x"38",
          9905 => x"5a",
          9906 => x"85",
          9907 => x"34",
          9908 => x"09",
          9909 => x"f6",
          9910 => x"ff",
          9911 => x"1d",
          9912 => x"84",
          9913 => x"93",
          9914 => x"74",
          9915 => x"9d",
          9916 => x"75",
          9917 => x"38",
          9918 => x"78",
          9919 => x"f7",
          9920 => x"07",
          9921 => x"57",
          9922 => x"a4",
          9923 => x"07",
          9924 => x"52",
          9925 => x"85",
          9926 => x"bb",
          9927 => x"ff",
          9928 => x"87",
          9929 => x"5a",
          9930 => x"2e",
          9931 => x"80",
          9932 => x"e7",
          9933 => x"56",
          9934 => x"ff",
          9935 => x"38",
          9936 => x"81",
          9937 => x"e6",
          9938 => x"e6",
          9939 => x"81",
          9940 => x"54",
          9941 => x"2e",
          9942 => x"73",
          9943 => x"38",
          9944 => x"33",
          9945 => x"06",
          9946 => x"73",
          9947 => x"81",
          9948 => x"78",
          9949 => x"ff",
          9950 => x"73",
          9951 => x"38",
          9952 => x"70",
          9953 => x"5f",
          9954 => x"15",
          9955 => x"26",
          9956 => x"81",
          9957 => x"ff",
          9958 => x"70",
          9959 => x"06",
          9960 => x"53",
          9961 => x"05",
          9962 => x"34",
          9963 => x"75",
          9964 => x"fc",
          9965 => x"fa",
          9966 => x"e6",
          9967 => x"81",
          9968 => x"53",
          9969 => x"ff",
          9970 => x"df",
          9971 => x"7d",
          9972 => x"5b",
          9973 => x"79",
          9974 => x"5b",
          9975 => x"cd",
          9976 => x"cc",
          9977 => x"98",
          9978 => x"2b",
          9979 => x"88",
          9980 => x"57",
          9981 => x"7b",
          9982 => x"75",
          9983 => x"54",
          9984 => x"81",
          9985 => x"a0",
          9986 => x"74",
          9987 => x"1b",
          9988 => x"39",
          9989 => x"a0",
          9990 => x"5a",
          9991 => x"2e",
          9992 => x"fa",
          9993 => x"a3",
          9994 => x"2a",
          9995 => x"7b",
          9996 => x"85",
          9997 => x"84",
          9998 => x"0d",
          9999 => x"0d",
         10000 => x"88",
         10001 => x"05",
         10002 => x"5e",
         10003 => x"ff",
         10004 => x"59",
         10005 => x"80",
         10006 => x"38",
         10007 => x"05",
         10008 => x"9f",
         10009 => x"75",
         10010 => x"d0",
         10011 => x"38",
         10012 => x"85",
         10013 => x"e2",
         10014 => x"80",
         10015 => x"b2",
         10016 => x"10",
         10017 => x"05",
         10018 => x"5a",
         10019 => x"80",
         10020 => x"38",
         10021 => x"7f",
         10022 => x"77",
         10023 => x"7b",
         10024 => x"38",
         10025 => x"51",
         10026 => x"3f",
         10027 => x"08",
         10028 => x"70",
         10029 => x"58",
         10030 => x"86",
         10031 => x"77",
         10032 => x"5d",
         10033 => x"1d",
         10034 => x"34",
         10035 => x"17",
         10036 => x"bb",
         10037 => x"bb",
         10038 => x"ff",
         10039 => x"06",
         10040 => x"58",
         10041 => x"38",
         10042 => x"8d",
         10043 => x"2a",
         10044 => x"8a",
         10045 => x"b1",
         10046 => x"7a",
         10047 => x"ff",
         10048 => x"0c",
         10049 => x"55",
         10050 => x"53",
         10051 => x"53",
         10052 => x"52",
         10053 => x"95",
         10054 => x"84",
         10055 => x"85",
         10056 => x"81",
         10057 => x"18",
         10058 => x"78",
         10059 => x"b7",
         10060 => x"b6",
         10061 => x"88",
         10062 => x"56",
         10063 => x"82",
         10064 => x"85",
         10065 => x"81",
         10066 => x"84",
         10067 => x"33",
         10068 => x"bf",
         10069 => x"75",
         10070 => x"cd",
         10071 => x"75",
         10072 => x"c5",
         10073 => x"17",
         10074 => x"18",
         10075 => x"2b",
         10076 => x"7c",
         10077 => x"09",
         10078 => x"ad",
         10079 => x"17",
         10080 => x"18",
         10081 => x"2b",
         10082 => x"75",
         10083 => x"dc",
         10084 => x"33",
         10085 => x"71",
         10086 => x"88",
         10087 => x"14",
         10088 => x"07",
         10089 => x"33",
         10090 => x"5a",
         10091 => x"5f",
         10092 => x"18",
         10093 => x"17",
         10094 => x"34",
         10095 => x"33",
         10096 => x"81",
         10097 => x"40",
         10098 => x"7c",
         10099 => x"d9",
         10100 => x"ff",
         10101 => x"29",
         10102 => x"33",
         10103 => x"77",
         10104 => x"77",
         10105 => x"2e",
         10106 => x"ff",
         10107 => x"42",
         10108 => x"38",
         10109 => x"33",
         10110 => x"33",
         10111 => x"07",
         10112 => x"88",
         10113 => x"75",
         10114 => x"5a",
         10115 => x"82",
         10116 => x"cc",
         10117 => x"cb",
         10118 => x"88",
         10119 => x"5c",
         10120 => x"80",
         10121 => x"11",
         10122 => x"33",
         10123 => x"71",
         10124 => x"81",
         10125 => x"72",
         10126 => x"75",
         10127 => x"53",
         10128 => x"42",
         10129 => x"c7",
         10130 => x"c6",
         10131 => x"88",
         10132 => x"58",
         10133 => x"80",
         10134 => x"38",
         10135 => x"84",
         10136 => x"79",
         10137 => x"c1",
         10138 => x"74",
         10139 => x"fd",
         10140 => x"84",
         10141 => x"56",
         10142 => x"08",
         10143 => x"a9",
         10144 => x"84",
         10145 => x"ff",
         10146 => x"83",
         10147 => x"75",
         10148 => x"26",
         10149 => x"5d",
         10150 => x"26",
         10151 => x"81",
         10152 => x"70",
         10153 => x"7b",
         10154 => x"7b",
         10155 => x"1a",
         10156 => x"b0",
         10157 => x"59",
         10158 => x"8a",
         10159 => x"17",
         10160 => x"58",
         10161 => x"80",
         10162 => x"16",
         10163 => x"78",
         10164 => x"82",
         10165 => x"78",
         10166 => x"81",
         10167 => x"06",
         10168 => x"83",
         10169 => x"2a",
         10170 => x"78",
         10171 => x"26",
         10172 => x"0b",
         10173 => x"ff",
         10174 => x"0c",
         10175 => x"84",
         10176 => x"83",
         10177 => x"38",
         10178 => x"84",
         10179 => x"81",
         10180 => x"84",
         10181 => x"7c",
         10182 => x"84",
         10183 => x"8c",
         10184 => x"0b",
         10185 => x"80",
         10186 => x"bb",
         10187 => x"3d",
         10188 => x"0b",
         10189 => x"0c",
         10190 => x"04",
         10191 => x"11",
         10192 => x"06",
         10193 => x"74",
         10194 => x"38",
         10195 => x"81",
         10196 => x"05",
         10197 => x"7a",
         10198 => x"38",
         10199 => x"83",
         10200 => x"40",
         10201 => x"7f",
         10202 => x"70",
         10203 => x"33",
         10204 => x"05",
         10205 => x"9f",
         10206 => x"56",
         10207 => x"89",
         10208 => x"70",
         10209 => x"57",
         10210 => x"17",
         10211 => x"26",
         10212 => x"17",
         10213 => x"06",
         10214 => x"30",
         10215 => x"59",
         10216 => x"2e",
         10217 => x"85",
         10218 => x"be",
         10219 => x"32",
         10220 => x"72",
         10221 => x"7a",
         10222 => x"55",
         10223 => x"87",
         10224 => x"1c",
         10225 => x"5c",
         10226 => x"ff",
         10227 => x"56",
         10228 => x"78",
         10229 => x"cf",
         10230 => x"2a",
         10231 => x"8a",
         10232 => x"c5",
         10233 => x"fe",
         10234 => x"78",
         10235 => x"75",
         10236 => x"09",
         10237 => x"38",
         10238 => x"81",
         10239 => x"30",
         10240 => x"7b",
         10241 => x"5c",
         10242 => x"38",
         10243 => x"2e",
         10244 => x"93",
         10245 => x"5a",
         10246 => x"fa",
         10247 => x"59",
         10248 => x"2e",
         10249 => x"81",
         10250 => x"80",
         10251 => x"90",
         10252 => x"2b",
         10253 => x"19",
         10254 => x"07",
         10255 => x"fe",
         10256 => x"07",
         10257 => x"40",
         10258 => x"7a",
         10259 => x"5c",
         10260 => x"90",
         10261 => x"78",
         10262 => x"be",
         10263 => x"f9",
         10264 => x"30",
         10265 => x"72",
         10266 => x"3d",
         10267 => x"05",
         10268 => x"b6",
         10269 => x"52",
         10270 => x"78",
         10271 => x"56",
         10272 => x"80",
         10273 => x"0b",
         10274 => x"ff",
         10275 => x"0c",
         10276 => x"56",
         10277 => x"a5",
         10278 => x"7a",
         10279 => x"52",
         10280 => x"51",
         10281 => x"3f",
         10282 => x"08",
         10283 => x"38",
         10284 => x"56",
         10285 => x"0c",
         10286 => x"bf",
         10287 => x"33",
         10288 => x"88",
         10289 => x"5e",
         10290 => x"82",
         10291 => x"09",
         10292 => x"38",
         10293 => x"18",
         10294 => x"75",
         10295 => x"82",
         10296 => x"81",
         10297 => x"30",
         10298 => x"7a",
         10299 => x"42",
         10300 => x"75",
         10301 => x"b6",
         10302 => x"77",
         10303 => x"56",
         10304 => x"ba",
         10305 => x"5d",
         10306 => x"2e",
         10307 => x"83",
         10308 => x"81",
         10309 => x"bd",
         10310 => x"2e",
         10311 => x"81",
         10312 => x"5a",
         10313 => x"27",
         10314 => x"f8",
         10315 => x"0b",
         10316 => x"83",
         10317 => x"5d",
         10318 => x"81",
         10319 => x"7e",
         10320 => x"40",
         10321 => x"31",
         10322 => x"52",
         10323 => x"80",
         10324 => x"38",
         10325 => x"e1",
         10326 => x"81",
         10327 => x"e6",
         10328 => x"58",
         10329 => x"05",
         10330 => x"70",
         10331 => x"33",
         10332 => x"ff",
         10333 => x"42",
         10334 => x"2e",
         10335 => x"75",
         10336 => x"38",
         10337 => x"f3",
         10338 => x"7c",
         10339 => x"77",
         10340 => x"0c",
         10341 => x"04",
         10342 => x"80",
         10343 => x"38",
         10344 => x"8a",
         10345 => x"b8",
         10346 => x"ff",
         10347 => x"0b",
         10348 => x"0c",
         10349 => x"04",
         10350 => x"ee",
         10351 => x"b4",
         10352 => x"78",
         10353 => x"5a",
         10354 => x"81",
         10355 => x"71",
         10356 => x"1b",
         10357 => x"5f",
         10358 => x"83",
         10359 => x"80",
         10360 => x"85",
         10361 => x"18",
         10362 => x"5c",
         10363 => x"70",
         10364 => x"33",
         10365 => x"05",
         10366 => x"71",
         10367 => x"5b",
         10368 => x"77",
         10369 => x"91",
         10370 => x"2e",
         10371 => x"3d",
         10372 => x"83",
         10373 => x"39",
         10374 => x"c6",
         10375 => x"17",
         10376 => x"18",
         10377 => x"2b",
         10378 => x"75",
         10379 => x"81",
         10380 => x"38",
         10381 => x"80",
         10382 => x"08",
         10383 => x"38",
         10384 => x"5b",
         10385 => x"09",
         10386 => x"9b",
         10387 => x"77",
         10388 => x"52",
         10389 => x"51",
         10390 => x"3f",
         10391 => x"08",
         10392 => x"38",
         10393 => x"5a",
         10394 => x"0c",
         10395 => x"38",
         10396 => x"34",
         10397 => x"33",
         10398 => x"33",
         10399 => x"07",
         10400 => x"82",
         10401 => x"09",
         10402 => x"fc",
         10403 => x"83",
         10404 => x"12",
         10405 => x"2b",
         10406 => x"07",
         10407 => x"70",
         10408 => x"2b",
         10409 => x"07",
         10410 => x"45",
         10411 => x"77",
         10412 => x"a4",
         10413 => x"81",
         10414 => x"38",
         10415 => x"83",
         10416 => x"12",
         10417 => x"2b",
         10418 => x"07",
         10419 => x"70",
         10420 => x"2b",
         10421 => x"07",
         10422 => x"5b",
         10423 => x"60",
         10424 => x"e4",
         10425 => x"81",
         10426 => x"38",
         10427 => x"83",
         10428 => x"12",
         10429 => x"2b",
         10430 => x"07",
         10431 => x"70",
         10432 => x"2b",
         10433 => x"07",
         10434 => x"5d",
         10435 => x"83",
         10436 => x"12",
         10437 => x"2b",
         10438 => x"07",
         10439 => x"70",
         10440 => x"2b",
         10441 => x"07",
         10442 => x"0c",
         10443 => x"46",
         10444 => x"45",
         10445 => x"7c",
         10446 => x"e2",
         10447 => x"05",
         10448 => x"e2",
         10449 => x"86",
         10450 => x"e2",
         10451 => x"18",
         10452 => x"98",
         10453 => x"cf",
         10454 => x"24",
         10455 => x"7b",
         10456 => x"56",
         10457 => x"75",
         10458 => x"08",
         10459 => x"70",
         10460 => x"33",
         10461 => x"af",
         10462 => x"bb",
         10463 => x"2e",
         10464 => x"81",
         10465 => x"bb",
         10466 => x"18",
         10467 => x"08",
         10468 => x"31",
         10469 => x"18",
         10470 => x"38",
         10471 => x"41",
         10472 => x"81",
         10473 => x"bb",
         10474 => x"fd",
         10475 => x"56",
         10476 => x"f3",
         10477 => x"0b",
         10478 => x"83",
         10479 => x"5a",
         10480 => x"39",
         10481 => x"33",
         10482 => x"33",
         10483 => x"07",
         10484 => x"58",
         10485 => x"38",
         10486 => x"42",
         10487 => x"38",
         10488 => x"83",
         10489 => x"12",
         10490 => x"2b",
         10491 => x"07",
         10492 => x"70",
         10493 => x"2b",
         10494 => x"07",
         10495 => x"5a",
         10496 => x"5a",
         10497 => x"59",
         10498 => x"39",
         10499 => x"80",
         10500 => x"38",
         10501 => x"e3",
         10502 => x"2e",
         10503 => x"93",
         10504 => x"5a",
         10505 => x"f2",
         10506 => x"79",
         10507 => x"fc",
         10508 => x"54",
         10509 => x"a0",
         10510 => x"53",
         10511 => x"17",
         10512 => x"ad",
         10513 => x"85",
         10514 => x"0d",
         10515 => x"05",
         10516 => x"43",
         10517 => x"57",
         10518 => x"5a",
         10519 => x"2e",
         10520 => x"78",
         10521 => x"5a",
         10522 => x"26",
         10523 => x"ba",
         10524 => x"38",
         10525 => x"74",
         10526 => x"d9",
         10527 => x"e0",
         10528 => x"74",
         10529 => x"38",
         10530 => x"84",
         10531 => x"70",
         10532 => x"73",
         10533 => x"38",
         10534 => x"62",
         10535 => x"2e",
         10536 => x"74",
         10537 => x"73",
         10538 => x"54",
         10539 => x"92",
         10540 => x"93",
         10541 => x"84",
         10542 => x"81",
         10543 => x"84",
         10544 => x"84",
         10545 => x"92",
         10546 => x"8b",
         10547 => x"84",
         10548 => x"0d",
         10549 => x"d0",
         10550 => x"ff",
         10551 => x"57",
         10552 => x"91",
         10553 => x"77",
         10554 => x"d0",
         10555 => x"77",
         10556 => x"f7",
         10557 => x"08",
         10558 => x"5e",
         10559 => x"08",
         10560 => x"79",
         10561 => x"5b",
         10562 => x"81",
         10563 => x"ff",
         10564 => x"57",
         10565 => x"26",
         10566 => x"15",
         10567 => x"06",
         10568 => x"9f",
         10569 => x"99",
         10570 => x"e0",
         10571 => x"ff",
         10572 => x"74",
         10573 => x"2a",
         10574 => x"76",
         10575 => x"06",
         10576 => x"ff",
         10577 => x"79",
         10578 => x"70",
         10579 => x"2a",
         10580 => x"57",
         10581 => x"2e",
         10582 => x"1b",
         10583 => x"5b",
         10584 => x"ff",
         10585 => x"54",
         10586 => x"7a",
         10587 => x"38",
         10588 => x"0c",
         10589 => x"39",
         10590 => x"6c",
         10591 => x"80",
         10592 => x"56",
         10593 => x"79",
         10594 => x"38",
         10595 => x"70",
         10596 => x"cc",
         10597 => x"3d",
         10598 => x"59",
         10599 => x"84",
         10600 => x"57",
         10601 => x"08",
         10602 => x"38",
         10603 => x"76",
         10604 => x"bb",
         10605 => x"3d",
         10606 => x"40",
         10607 => x"3d",
         10608 => x"e1",
         10609 => x"bb",
         10610 => x"84",
         10611 => x"80",
         10612 => x"38",
         10613 => x"5d",
         10614 => x"81",
         10615 => x"80",
         10616 => x"38",
         10617 => x"84",
         10618 => x"88",
         10619 => x"ff",
         10620 => x"83",
         10621 => x"58",
         10622 => x"81",
         10623 => x"9b",
         10624 => x"12",
         10625 => x"2b",
         10626 => x"33",
         10627 => x"5e",
         10628 => x"2e",
         10629 => x"80",
         10630 => x"34",
         10631 => x"17",
         10632 => x"90",
         10633 => x"cc",
         10634 => x"34",
         10635 => x"0b",
         10636 => x"7e",
         10637 => x"80",
         10638 => x"34",
         10639 => x"17",
         10640 => x"5d",
         10641 => x"85",
         10642 => x"58",
         10643 => x"19",
         10644 => x"9d",
         10645 => x"0b",
         10646 => x"80",
         10647 => x"34",
         10648 => x"0b",
         10649 => x"7a",
         10650 => x"e2",
         10651 => x"11",
         10652 => x"08",
         10653 => x"57",
         10654 => x"89",
         10655 => x"08",
         10656 => x"ec",
         10657 => x"80",
         10658 => x"a3",
         10659 => x"e7",
         10660 => x"98",
         10661 => x"7a",
         10662 => x"b8",
         10663 => x"9c",
         10664 => x"7c",
         10665 => x"76",
         10666 => x"02",
         10667 => x"33",
         10668 => x"81",
         10669 => x"7b",
         10670 => x"78",
         10671 => x"06",
         10672 => x"2e",
         10673 => x"81",
         10674 => x"82",
         10675 => x"83",
         10676 => x"56",
         10677 => x"86",
         10678 => x"c0",
         10679 => x"b4",
         10680 => x"1c",
         10681 => x"1c",
         10682 => x"11",
         10683 => x"33",
         10684 => x"07",
         10685 => x"5b",
         10686 => x"7b",
         10687 => x"fb",
         10688 => x"1b",
         10689 => x"83",
         10690 => x"12",
         10691 => x"2b",
         10692 => x"07",
         10693 => x"70",
         10694 => x"2b",
         10695 => x"07",
         10696 => x"0c",
         10697 => x"0c",
         10698 => x"59",
         10699 => x"22",
         10700 => x"78",
         10701 => x"80",
         10702 => x"34",
         10703 => x"1b",
         10704 => x"94",
         10705 => x"1a",
         10706 => x"7c",
         10707 => x"76",
         10708 => x"58",
         10709 => x"55",
         10710 => x"78",
         10711 => x"06",
         10712 => x"2e",
         10713 => x"8c",
         10714 => x"74",
         10715 => x"bf",
         10716 => x"1b",
         10717 => x"22",
         10718 => x"88",
         10719 => x"59",
         10720 => x"76",
         10721 => x"07",
         10722 => x"55",
         10723 => x"83",
         10724 => x"70",
         10725 => x"5b",
         10726 => x"83",
         10727 => x"52",
         10728 => x"ac",
         10729 => x"bb",
         10730 => x"84",
         10731 => x"81",
         10732 => x"82",
         10733 => x"84",
         10734 => x"b6",
         10735 => x"31",
         10736 => x"02",
         10737 => x"33",
         10738 => x"7d",
         10739 => x"82",
         10740 => x"55",
         10741 => x"fc",
         10742 => x"57",
         10743 => x"fb",
         10744 => x"57",
         10745 => x"fb",
         10746 => x"57",
         10747 => x"fb",
         10748 => x"76",
         10749 => x"57",
         10750 => x"95",
         10751 => x"17",
         10752 => x"2b",
         10753 => x"07",
         10754 => x"1d",
         10755 => x"83",
         10756 => x"12",
         10757 => x"2b",
         10758 => x"07",
         10759 => x"70",
         10760 => x"2b",
         10761 => x"07",
         10762 => x"0c",
         10763 => x"0c",
         10764 => x"5b",
         10765 => x"86",
         10766 => x"1b",
         10767 => x"1b",
         10768 => x"91",
         10769 => x"0b",
         10770 => x"80",
         10771 => x"0c",
         10772 => x"84",
         10773 => x"55",
         10774 => x"7b",
         10775 => x"3f",
         10776 => x"08",
         10777 => x"5a",
         10778 => x"c0",
         10779 => x"39",
         10780 => x"51",
         10781 => x"3f",
         10782 => x"08",
         10783 => x"84",
         10784 => x"80",
         10785 => x"bb",
         10786 => x"2e",
         10787 => x"84",
         10788 => x"ff",
         10789 => x"38",
         10790 => x"52",
         10791 => x"b1",
         10792 => x"bb",
         10793 => x"8f",
         10794 => x"08",
         10795 => x"18",
         10796 => x"58",
         10797 => x"90",
         10798 => x"94",
         10799 => x"16",
         10800 => x"55",
         10801 => x"34",
         10802 => x"7d",
         10803 => x"38",
         10804 => x"72",
         10805 => x"5d",
         10806 => x"7e",
         10807 => x"83",
         10808 => x"77",
         10809 => x"81",
         10810 => x"38",
         10811 => x"53",
         10812 => x"81",
         10813 => x"ff",
         10814 => x"84",
         10815 => x"80",
         10816 => x"ff",
         10817 => x"76",
         10818 => x"7e",
         10819 => x"1c",
         10820 => x"57",
         10821 => x"fb",
         10822 => x"7a",
         10823 => x"39",
         10824 => x"17",
         10825 => x"95",
         10826 => x"9e",
         10827 => x"33",
         10828 => x"71",
         10829 => x"90",
         10830 => x"07",
         10831 => x"80",
         10832 => x"34",
         10833 => x"17",
         10834 => x"90",
         10835 => x"cc",
         10836 => x"34",
         10837 => x"0b",
         10838 => x"7e",
         10839 => x"80",
         10840 => x"34",
         10841 => x"17",
         10842 => x"5d",
         10843 => x"09",
         10844 => x"d6",
         10845 => x"39",
         10846 => x"0c",
         10847 => x"38",
         10848 => x"06",
         10849 => x"2e",
         10850 => x"7e",
         10851 => x"12",
         10852 => x"40",
         10853 => x"7e",
         10854 => x"38",
         10855 => x"78",
         10856 => x"1b",
         10857 => x"5b",
         10858 => x"f9",
         10859 => x"89",
         10860 => x"9c",
         10861 => x"81",
         10862 => x"7b",
         10863 => x"33",
         10864 => x"e9",
         10865 => x"84",
         10866 => x"f7",
         10867 => x"57",
         10868 => x"f7",
         10869 => x"54",
         10870 => x"53",
         10871 => x"53",
         10872 => x"52",
         10873 => x"c4",
         10874 => x"84",
         10875 => x"09",
         10876 => x"ce",
         10877 => x"84",
         10878 => x"34",
         10879 => x"a8",
         10880 => x"84",
         10881 => x"5d",
         10882 => x"17",
         10883 => x"dc",
         10884 => x"33",
         10885 => x"2e",
         10886 => x"fd",
         10887 => x"54",
         10888 => x"a0",
         10889 => x"53",
         10890 => x"16",
         10891 => x"a1",
         10892 => x"5c",
         10893 => x"84",
         10894 => x"57",
         10895 => x"f6",
         10896 => x"5c",
         10897 => x"f2",
         10898 => x"63",
         10899 => x"40",
         10900 => x"7e",
         10901 => x"78",
         10902 => x"38",
         10903 => x"75",
         10904 => x"38",
         10905 => x"74",
         10906 => x"38",
         10907 => x"84",
         10908 => x"5b",
         10909 => x"83",
         10910 => x"55",
         10911 => x"55",
         10912 => x"38",
         10913 => x"55",
         10914 => x"38",
         10915 => x"81",
         10916 => x"56",
         10917 => x"81",
         10918 => x"19",
         10919 => x"08",
         10920 => x"56",
         10921 => x"81",
         10922 => x"80",
         10923 => x"38",
         10924 => x"06",
         10925 => x"99",
         10926 => x"11",
         10927 => x"77",
         10928 => x"5d",
         10929 => x"38",
         10930 => x"38",
         10931 => x"55",
         10932 => x"83",
         10933 => x"ff",
         10934 => x"38",
         10935 => x"0c",
         10936 => x"19",
         10937 => x"9c",
         10938 => x"05",
         10939 => x"7b",
         10940 => x"38",
         10941 => x"70",
         10942 => x"1a",
         10943 => x"56",
         10944 => x"83",
         10945 => x"15",
         10946 => x"5c",
         10947 => x"2e",
         10948 => x"7a",
         10949 => x"75",
         10950 => x"75",
         10951 => x"7a",
         10952 => x"7c",
         10953 => x"33",
         10954 => x"81",
         10955 => x"84",
         10956 => x"38",
         10957 => x"70",
         10958 => x"56",
         10959 => x"82",
         10960 => x"89",
         10961 => x"77",
         10962 => x"18",
         10963 => x"1e",
         10964 => x"19",
         10965 => x"1c",
         10966 => x"79",
         10967 => x"80",
         10968 => x"bb",
         10969 => x"3d",
         10970 => x"84",
         10971 => x"90",
         10972 => x"74",
         10973 => x"39",
         10974 => x"56",
         10975 => x"80",
         10976 => x"19",
         10977 => x"2b",
         10978 => x"5d",
         10979 => x"25",
         10980 => x"54",
         10981 => x"52",
         10982 => x"51",
         10983 => x"3f",
         10984 => x"08",
         10985 => x"90",
         10986 => x"ff",
         10987 => x"90",
         10988 => x"58",
         10989 => x"53",
         10990 => x"18",
         10991 => x"9d",
         10992 => x"bb",
         10993 => x"c1",
         10994 => x"1a",
         10995 => x"08",
         10996 => x"ff",
         10997 => x"71",
         10998 => x"79",
         10999 => x"38",
         11000 => x"7d",
         11001 => x"05",
         11002 => x"76",
         11003 => x"d6",
         11004 => x"81",
         11005 => x"78",
         11006 => x"5a",
         11007 => x"56",
         11008 => x"fe",
         11009 => x"70",
         11010 => x"33",
         11011 => x"05",
         11012 => x"16",
         11013 => x"38",
         11014 => x"98",
         11015 => x"78",
         11016 => x"bc",
         11017 => x"84",
         11018 => x"a4",
         11019 => x"33",
         11020 => x"a7",
         11021 => x"84",
         11022 => x"55",
         11023 => x"38",
         11024 => x"56",
         11025 => x"39",
         11026 => x"77",
         11027 => x"7b",
         11028 => x"38",
         11029 => x"71",
         11030 => x"1b",
         11031 => x"75",
         11032 => x"57",
         11033 => x"81",
         11034 => x"ff",
         11035 => x"80",
         11036 => x"38",
         11037 => x"05",
         11038 => x"70",
         11039 => x"34",
         11040 => x"74",
         11041 => x"ba",
         11042 => x"91",
         11043 => x"0b",
         11044 => x"0c",
         11045 => x"04",
         11046 => x"1a",
         11047 => x"84",
         11048 => x"90",
         11049 => x"f1",
         11050 => x"64",
         11051 => x"41",
         11052 => x"7f",
         11053 => x"78",
         11054 => x"38",
         11055 => x"75",
         11056 => x"38",
         11057 => x"74",
         11058 => x"38",
         11059 => x"84",
         11060 => x"5a",
         11061 => x"84",
         11062 => x"55",
         11063 => x"55",
         11064 => x"38",
         11065 => x"55",
         11066 => x"38",
         11067 => x"70",
         11068 => x"06",
         11069 => x"56",
         11070 => x"82",
         11071 => x"19",
         11072 => x"5d",
         11073 => x"27",
         11074 => x"09",
         11075 => x"2e",
         11076 => x"76",
         11077 => x"5d",
         11078 => x"38",
         11079 => x"22",
         11080 => x"89",
         11081 => x"58",
         11082 => x"76",
         11083 => x"88",
         11084 => x"74",
         11085 => x"8c",
         11086 => x"2e",
         11087 => x"74",
         11088 => x"d8",
         11089 => x"1a",
         11090 => x"08",
         11091 => x"88",
         11092 => x"58",
         11093 => x"70",
         11094 => x"57",
         11095 => x"82",
         11096 => x"19",
         11097 => x"9c",
         11098 => x"05",
         11099 => x"7c",
         11100 => x"38",
         11101 => x"70",
         11102 => x"1a",
         11103 => x"56",
         11104 => x"83",
         11105 => x"15",
         11106 => x"5b",
         11107 => x"2e",
         11108 => x"79",
         11109 => x"75",
         11110 => x"75",
         11111 => x"79",
         11112 => x"7d",
         11113 => x"33",
         11114 => x"80",
         11115 => x"84",
         11116 => x"38",
         11117 => x"7c",
         11118 => x"7a",
         11119 => x"84",
         11120 => x"1a",
         11121 => x"60",
         11122 => x"55",
         11123 => x"05",
         11124 => x"70",
         11125 => x"34",
         11126 => x"74",
         11127 => x"19",
         11128 => x"06",
         11129 => x"1a",
         11130 => x"2b",
         11131 => x"31",
         11132 => x"60",
         11133 => x"94",
         11134 => x"70",
         11135 => x"0c",
         11136 => x"59",
         11137 => x"5b",
         11138 => x"83",
         11139 => x"74",
         11140 => x"7a",
         11141 => x"90",
         11142 => x"77",
         11143 => x"5b",
         11144 => x"34",
         11145 => x"84",
         11146 => x"91",
         11147 => x"74",
         11148 => x"0c",
         11149 => x"04",
         11150 => x"7c",
         11151 => x"94",
         11152 => x"76",
         11153 => x"27",
         11154 => x"54",
         11155 => x"19",
         11156 => x"33",
         11157 => x"d5",
         11158 => x"84",
         11159 => x"38",
         11160 => x"57",
         11161 => x"0c",
         11162 => x"06",
         11163 => x"31",
         11164 => x"78",
         11165 => x"7a",
         11166 => x"16",
         11167 => x"59",
         11168 => x"80",
         11169 => x"76",
         11170 => x"58",
         11171 => x"81",
         11172 => x"ff",
         11173 => x"ef",
         11174 => x"33",
         11175 => x"5a",
         11176 => x"34",
         11177 => x"98",
         11178 => x"78",
         11179 => x"ef",
         11180 => x"84",
         11181 => x"bb",
         11182 => x"fd",
         11183 => x"33",
         11184 => x"39",
         11185 => x"51",
         11186 => x"3f",
         11187 => x"08",
         11188 => x"84",
         11189 => x"38",
         11190 => x"54",
         11191 => x"53",
         11192 => x"81",
         11193 => x"ff",
         11194 => x"84",
         11195 => x"ac",
         11196 => x"33",
         11197 => x"56",
         11198 => x"34",
         11199 => x"e2",
         11200 => x"33",
         11201 => x"d3",
         11202 => x"84",
         11203 => x"55",
         11204 => x"38",
         11205 => x"56",
         11206 => x"39",
         11207 => x"1a",
         11208 => x"84",
         11209 => x"91",
         11210 => x"82",
         11211 => x"34",
         11212 => x"bb",
         11213 => x"3d",
         11214 => x"3d",
         11215 => x"89",
         11216 => x"2e",
         11217 => x"08",
         11218 => x"2e",
         11219 => x"33",
         11220 => x"2e",
         11221 => x"16",
         11222 => x"22",
         11223 => x"79",
         11224 => x"38",
         11225 => x"5c",
         11226 => x"81",
         11227 => x"18",
         11228 => x"2a",
         11229 => x"57",
         11230 => x"81",
         11231 => x"98",
         11232 => x"76",
         11233 => x"38",
         11234 => x"08",
         11235 => x"16",
         11236 => x"b8",
         11237 => x"83",
         11238 => x"5b",
         11239 => x"7a",
         11240 => x"06",
         11241 => x"81",
         11242 => x"b8",
         11243 => x"16",
         11244 => x"95",
         11245 => x"bb",
         11246 => x"2e",
         11247 => x"57",
         11248 => x"b4",
         11249 => x"56",
         11250 => x"38",
         11251 => x"8b",
         11252 => x"07",
         11253 => x"8b",
         11254 => x"08",
         11255 => x"70",
         11256 => x"06",
         11257 => x"7a",
         11258 => x"7a",
         11259 => x"79",
         11260 => x"9c",
         11261 => x"96",
         11262 => x"5b",
         11263 => x"81",
         11264 => x"18",
         11265 => x"7b",
         11266 => x"2a",
         11267 => x"18",
         11268 => x"2a",
         11269 => x"18",
         11270 => x"2a",
         11271 => x"18",
         11272 => x"34",
         11273 => x"18",
         11274 => x"98",
         11275 => x"cc",
         11276 => x"34",
         11277 => x"18",
         11278 => x"93",
         11279 => x"5b",
         11280 => x"1c",
         11281 => x"ff",
         11282 => x"84",
         11283 => x"90",
         11284 => x"bf",
         11285 => x"79",
         11286 => x"75",
         11287 => x"bb",
         11288 => x"3d",
         11289 => x"54",
         11290 => x"53",
         11291 => x"53",
         11292 => x"52",
         11293 => x"b4",
         11294 => x"84",
         11295 => x"7a",
         11296 => x"06",
         11297 => x"84",
         11298 => x"83",
         11299 => x"16",
         11300 => x"08",
         11301 => x"84",
         11302 => x"74",
         11303 => x"27",
         11304 => x"82",
         11305 => x"74",
         11306 => x"81",
         11307 => x"38",
         11308 => x"16",
         11309 => x"08",
         11310 => x"52",
         11311 => x"51",
         11312 => x"3f",
         11313 => x"df",
         11314 => x"2a",
         11315 => x"18",
         11316 => x"2a",
         11317 => x"18",
         11318 => x"08",
         11319 => x"34",
         11320 => x"5b",
         11321 => x"34",
         11322 => x"56",
         11323 => x"34",
         11324 => x"59",
         11325 => x"34",
         11326 => x"80",
         11327 => x"34",
         11328 => x"18",
         11329 => x"0b",
         11330 => x"80",
         11331 => x"34",
         11332 => x"18",
         11333 => x"81",
         11334 => x"34",
         11335 => x"96",
         11336 => x"bb",
         11337 => x"19",
         11338 => x"06",
         11339 => x"90",
         11340 => x"a7",
         11341 => x"33",
         11342 => x"9f",
         11343 => x"84",
         11344 => x"55",
         11345 => x"38",
         11346 => x"56",
         11347 => x"39",
         11348 => x"18",
         11349 => x"18",
         11350 => x"11",
         11351 => x"ff",
         11352 => x"81",
         11353 => x"84",
         11354 => x"38",
         11355 => x"80",
         11356 => x"78",
         11357 => x"7b",
         11358 => x"58",
         11359 => x"08",
         11360 => x"81",
         11361 => x"38",
         11362 => x"f9",
         11363 => x"70",
         11364 => x"a6",
         11365 => x"84",
         11366 => x"bb",
         11367 => x"38",
         11368 => x"80",
         11369 => x"74",
         11370 => x"80",
         11371 => x"72",
         11372 => x"80",
         11373 => x"86",
         11374 => x"16",
         11375 => x"71",
         11376 => x"38",
         11377 => x"58",
         11378 => x"84",
         11379 => x"0c",
         11380 => x"84",
         11381 => x"0d",
         11382 => x"33",
         11383 => x"fb",
         11384 => x"84",
         11385 => x"53",
         11386 => x"73",
         11387 => x"56",
         11388 => x"3d",
         11389 => x"70",
         11390 => x"75",
         11391 => x"38",
         11392 => x"05",
         11393 => x"9f",
         11394 => x"71",
         11395 => x"38",
         11396 => x"71",
         11397 => x"38",
         11398 => x"33",
         11399 => x"24",
         11400 => x"84",
         11401 => x"80",
         11402 => x"84",
         11403 => x"0d",
         11404 => x"84",
         11405 => x"8c",
         11406 => x"78",
         11407 => x"70",
         11408 => x"53",
         11409 => x"89",
         11410 => x"82",
         11411 => x"ff",
         11412 => x"59",
         11413 => x"2e",
         11414 => x"80",
         11415 => x"f4",
         11416 => x"08",
         11417 => x"76",
         11418 => x"58",
         11419 => x"81",
         11420 => x"ff",
         11421 => x"54",
         11422 => x"26",
         11423 => x"12",
         11424 => x"06",
         11425 => x"9f",
         11426 => x"99",
         11427 => x"e0",
         11428 => x"ff",
         11429 => x"71",
         11430 => x"2a",
         11431 => x"73",
         11432 => x"06",
         11433 => x"ff",
         11434 => x"76",
         11435 => x"70",
         11436 => x"2a",
         11437 => x"52",
         11438 => x"2e",
         11439 => x"18",
         11440 => x"58",
         11441 => x"ff",
         11442 => x"51",
         11443 => x"77",
         11444 => x"38",
         11445 => x"51",
         11446 => x"ea",
         11447 => x"53",
         11448 => x"05",
         11449 => x"51",
         11450 => x"84",
         11451 => x"55",
         11452 => x"08",
         11453 => x"38",
         11454 => x"84",
         11455 => x"0d",
         11456 => x"68",
         11457 => x"d0",
         11458 => x"d3",
         11459 => x"84",
         11460 => x"bb",
         11461 => x"c6",
         11462 => x"d7",
         11463 => x"98",
         11464 => x"80",
         11465 => x"e2",
         11466 => x"05",
         11467 => x"2a",
         11468 => x"59",
         11469 => x"b2",
         11470 => x"9b",
         11471 => x"12",
         11472 => x"2b",
         11473 => x"5e",
         11474 => x"58",
         11475 => x"a4",
         11476 => x"19",
         11477 => x"bb",
         11478 => x"3d",
         11479 => x"bb",
         11480 => x"2e",
         11481 => x"ff",
         11482 => x"0b",
         11483 => x"0c",
         11484 => x"04",
         11485 => x"94",
         11486 => x"98",
         11487 => x"2b",
         11488 => x"98",
         11489 => x"54",
         11490 => x"7e",
         11491 => x"58",
         11492 => x"84",
         11493 => x"0d",
         11494 => x"3d",
         11495 => x"3d",
         11496 => x"3d",
         11497 => x"80",
         11498 => x"53",
         11499 => x"fd",
         11500 => x"80",
         11501 => x"d1",
         11502 => x"bb",
         11503 => x"84",
         11504 => x"83",
         11505 => x"80",
         11506 => x"7f",
         11507 => x"08",
         11508 => x"0c",
         11509 => x"3d",
         11510 => x"79",
         11511 => x"cc",
         11512 => x"3d",
         11513 => x"5b",
         11514 => x"51",
         11515 => x"3f",
         11516 => x"08",
         11517 => x"84",
         11518 => x"38",
         11519 => x"3d",
         11520 => x"b4",
         11521 => x"2e",
         11522 => x"bb",
         11523 => x"17",
         11524 => x"7d",
         11525 => x"81",
         11526 => x"b8",
         11527 => x"16",
         11528 => x"8d",
         11529 => x"bb",
         11530 => x"2e",
         11531 => x"57",
         11532 => x"b4",
         11533 => x"82",
         11534 => x"df",
         11535 => x"11",
         11536 => x"33",
         11537 => x"07",
         11538 => x"5d",
         11539 => x"56",
         11540 => x"82",
         11541 => x"80",
         11542 => x"80",
         11543 => x"ff",
         11544 => x"84",
         11545 => x"59",
         11546 => x"08",
         11547 => x"80",
         11548 => x"ff",
         11549 => x"84",
         11550 => x"59",
         11551 => x"08",
         11552 => x"df",
         11553 => x"11",
         11554 => x"33",
         11555 => x"07",
         11556 => x"42",
         11557 => x"56",
         11558 => x"81",
         11559 => x"7a",
         11560 => x"84",
         11561 => x"52",
         11562 => x"a6",
         11563 => x"bb",
         11564 => x"84",
         11565 => x"80",
         11566 => x"38",
         11567 => x"83",
         11568 => x"81",
         11569 => x"e4",
         11570 => x"05",
         11571 => x"ff",
         11572 => x"78",
         11573 => x"33",
         11574 => x"80",
         11575 => x"82",
         11576 => x"17",
         11577 => x"33",
         11578 => x"7c",
         11579 => x"17",
         11580 => x"26",
         11581 => x"76",
         11582 => x"38",
         11583 => x"05",
         11584 => x"80",
         11585 => x"11",
         11586 => x"19",
         11587 => x"58",
         11588 => x"34",
         11589 => x"ff",
         11590 => x"3d",
         11591 => x"58",
         11592 => x"80",
         11593 => x"5a",
         11594 => x"38",
         11595 => x"82",
         11596 => x"0b",
         11597 => x"33",
         11598 => x"83",
         11599 => x"70",
         11600 => x"43",
         11601 => x"5a",
         11602 => x"8d",
         11603 => x"70",
         11604 => x"57",
         11605 => x"f5",
         11606 => x"5b",
         11607 => x"ab",
         11608 => x"76",
         11609 => x"38",
         11610 => x"7e",
         11611 => x"81",
         11612 => x"81",
         11613 => x"77",
         11614 => x"ba",
         11615 => x"05",
         11616 => x"ff",
         11617 => x"06",
         11618 => x"91",
         11619 => x"34",
         11620 => x"84",
         11621 => x"3d",
         11622 => x"16",
         11623 => x"33",
         11624 => x"71",
         11625 => x"79",
         11626 => x"5e",
         11627 => x"95",
         11628 => x"17",
         11629 => x"2b",
         11630 => x"07",
         11631 => x"dd",
         11632 => x"5d",
         11633 => x"51",
         11634 => x"3f",
         11635 => x"08",
         11636 => x"84",
         11637 => x"fd",
         11638 => x"b1",
         11639 => x"b4",
         11640 => x"b8",
         11641 => x"81",
         11642 => x"5e",
         11643 => x"3f",
         11644 => x"bb",
         11645 => x"be",
         11646 => x"84",
         11647 => x"34",
         11648 => x"a8",
         11649 => x"84",
         11650 => x"5a",
         11651 => x"17",
         11652 => x"83",
         11653 => x"33",
         11654 => x"2e",
         11655 => x"fb",
         11656 => x"54",
         11657 => x"a0",
         11658 => x"53",
         11659 => x"16",
         11660 => x"89",
         11661 => x"59",
         11662 => x"ff",
         11663 => x"3d",
         11664 => x"58",
         11665 => x"80",
         11666 => x"e0",
         11667 => x"10",
         11668 => x"05",
         11669 => x"33",
         11670 => x"5e",
         11671 => x"2e",
         11672 => x"fd",
         11673 => x"f1",
         11674 => x"3d",
         11675 => x"19",
         11676 => x"33",
         11677 => x"05",
         11678 => x"60",
         11679 => x"38",
         11680 => x"08",
         11681 => x"59",
         11682 => x"7c",
         11683 => x"5e",
         11684 => x"26",
         11685 => x"f5",
         11686 => x"80",
         11687 => x"84",
         11688 => x"80",
         11689 => x"04",
         11690 => x"7d",
         11691 => x"89",
         11692 => x"2e",
         11693 => x"08",
         11694 => x"2e",
         11695 => x"33",
         11696 => x"2e",
         11697 => x"16",
         11698 => x"22",
         11699 => x"7a",
         11700 => x"38",
         11701 => x"5c",
         11702 => x"82",
         11703 => x"17",
         11704 => x"82",
         11705 => x"17",
         11706 => x"78",
         11707 => x"38",
         11708 => x"56",
         11709 => x"7a",
         11710 => x"38",
         11711 => x"22",
         11712 => x"52",
         11713 => x"7a",
         11714 => x"38",
         11715 => x"19",
         11716 => x"93",
         11717 => x"84",
         11718 => x"79",
         11719 => x"57",
         11720 => x"83",
         11721 => x"84",
         11722 => x"82",
         11723 => x"30",
         11724 => x"94",
         11725 => x"71",
         11726 => x"08",
         11727 => x"75",
         11728 => x"92",
         11729 => x"27",
         11730 => x"78",
         11731 => x"18",
         11732 => x"19",
         11733 => x"33",
         11734 => x"81",
         11735 => x"59",
         11736 => x"82",
         11737 => x"52",
         11738 => x"9b",
         11739 => x"bb",
         11740 => x"84",
         11741 => x"80",
         11742 => x"75",
         11743 => x"d1",
         11744 => x"27",
         11745 => x"7b",
         11746 => x"16",
         11747 => x"f8",
         11748 => x"18",
         11749 => x"39",
         11750 => x"08",
         11751 => x"08",
         11752 => x"0c",
         11753 => x"06",
         11754 => x"2e",
         11755 => x"fe",
         11756 => x"08",
         11757 => x"57",
         11758 => x"27",
         11759 => x"8a",
         11760 => x"71",
         11761 => x"08",
         11762 => x"2a",
         11763 => x"55",
         11764 => x"82",
         11765 => x"17",
         11766 => x"17",
         11767 => x"76",
         11768 => x"75",
         11769 => x"90",
         11770 => x"c0",
         11771 => x"90",
         11772 => x"83",
         11773 => x"7a",
         11774 => x"ab",
         11775 => x"08",
         11776 => x"2e",
         11777 => x"90",
         11778 => x"98",
         11779 => x"5a",
         11780 => x"80",
         11781 => x"81",
         11782 => x"77",
         11783 => x"11",
         11784 => x"ff",
         11785 => x"84",
         11786 => x"a5",
         11787 => x"33",
         11788 => x"55",
         11789 => x"34",
         11790 => x"53",
         11791 => x"81",
         11792 => x"58",
         11793 => x"3f",
         11794 => x"08",
         11795 => x"d3",
         11796 => x"91",
         11797 => x"55",
         11798 => x"84",
         11799 => x"0d",
         11800 => x"33",
         11801 => x"81",
         11802 => x"75",
         11803 => x"77",
         11804 => x"57",
         11805 => x"78",
         11806 => x"81",
         11807 => x"38",
         11808 => x"0c",
         11809 => x"80",
         11810 => x"0c",
         11811 => x"56",
         11812 => x"80",
         11813 => x"98",
         11814 => x"80",
         11815 => x"38",
         11816 => x"79",
         11817 => x"80",
         11818 => x"84",
         11819 => x"0d",
         11820 => x"76",
         11821 => x"a8",
         11822 => x"84",
         11823 => x"bb",
         11824 => x"33",
         11825 => x"93",
         11826 => x"84",
         11827 => x"55",
         11828 => x"38",
         11829 => x"56",
         11830 => x"39",
         11831 => x"51",
         11832 => x"3f",
         11833 => x"08",
         11834 => x"84",
         11835 => x"98",
         11836 => x"84",
         11837 => x"fe",
         11838 => x"bb",
         11839 => x"18",
         11840 => x"18",
         11841 => x"39",
         11842 => x"18",
         11843 => x"84",
         11844 => x"8d",
         11845 => x"f6",
         11846 => x"56",
         11847 => x"80",
         11848 => x"80",
         11849 => x"fc",
         11850 => x"3d",
         11851 => x"c6",
         11852 => x"bb",
         11853 => x"84",
         11854 => x"80",
         11855 => x"80",
         11856 => x"54",
         11857 => x"84",
         11858 => x"0d",
         11859 => x"0c",
         11860 => x"51",
         11861 => x"3f",
         11862 => x"08",
         11863 => x"84",
         11864 => x"38",
         11865 => x"70",
         11866 => x"59",
         11867 => x"af",
         11868 => x"33",
         11869 => x"81",
         11870 => x"79",
         11871 => x"c5",
         11872 => x"08",
         11873 => x"9a",
         11874 => x"88",
         11875 => x"70",
         11876 => x"5a",
         11877 => x"83",
         11878 => x"77",
         11879 => x"7a",
         11880 => x"22",
         11881 => x"74",
         11882 => x"ff",
         11883 => x"84",
         11884 => x"55",
         11885 => x"8d",
         11886 => x"2e",
         11887 => x"80",
         11888 => x"fe",
         11889 => x"80",
         11890 => x"f6",
         11891 => x"33",
         11892 => x"71",
         11893 => x"90",
         11894 => x"07",
         11895 => x"5a",
         11896 => x"39",
         11897 => x"78",
         11898 => x"74",
         11899 => x"38",
         11900 => x"72",
         11901 => x"38",
         11902 => x"71",
         11903 => x"38",
         11904 => x"84",
         11905 => x"52",
         11906 => x"94",
         11907 => x"71",
         11908 => x"38",
         11909 => x"73",
         11910 => x"0c",
         11911 => x"04",
         11912 => x"51",
         11913 => x"3f",
         11914 => x"08",
         11915 => x"71",
         11916 => x"75",
         11917 => x"d7",
         11918 => x"0d",
         11919 => x"55",
         11920 => x"80",
         11921 => x"74",
         11922 => x"80",
         11923 => x"73",
         11924 => x"80",
         11925 => x"86",
         11926 => x"16",
         11927 => x"72",
         11928 => x"97",
         11929 => x"72",
         11930 => x"75",
         11931 => x"76",
         11932 => x"f3",
         11933 => x"74",
         11934 => x"ae",
         11935 => x"84",
         11936 => x"bb",
         11937 => x"2e",
         11938 => x"bb",
         11939 => x"38",
         11940 => x"51",
         11941 => x"3f",
         11942 => x"51",
         11943 => x"3f",
         11944 => x"08",
         11945 => x"30",
         11946 => x"9f",
         11947 => x"84",
         11948 => x"57",
         11949 => x"bb",
         11950 => x"3d",
         11951 => x"77",
         11952 => x"53",
         11953 => x"3f",
         11954 => x"51",
         11955 => x"3f",
         11956 => x"08",
         11957 => x"30",
         11958 => x"9f",
         11959 => x"84",
         11960 => x"57",
         11961 => x"75",
         11962 => x"ff",
         11963 => x"84",
         11964 => x"84",
         11965 => x"8a",
         11966 => x"81",
         11967 => x"fe",
         11968 => x"84",
         11969 => x"81",
         11970 => x"fe",
         11971 => x"75",
         11972 => x"fe",
         11973 => x"3d",
         11974 => x"80",
         11975 => x"70",
         11976 => x"52",
         11977 => x"3f",
         11978 => x"08",
         11979 => x"84",
         11980 => x"8a",
         11981 => x"bb",
         11982 => x"3d",
         11983 => x"52",
         11984 => x"b6",
         11985 => x"bb",
         11986 => x"84",
         11987 => x"e5",
         11988 => x"cb",
         11989 => x"98",
         11990 => x"80",
         11991 => x"38",
         11992 => x"d1",
         11993 => x"75",
         11994 => x"ae",
         11995 => x"bb",
         11996 => x"3d",
         11997 => x"0b",
         11998 => x"0c",
         11999 => x"04",
         12000 => x"66",
         12001 => x"80",
         12002 => x"ec",
         12003 => x"3d",
         12004 => x"3f",
         12005 => x"08",
         12006 => x"84",
         12007 => x"7f",
         12008 => x"08",
         12009 => x"fe",
         12010 => x"08",
         12011 => x"57",
         12012 => x"8d",
         12013 => x"0c",
         12014 => x"84",
         12015 => x"0d",
         12016 => x"84",
         12017 => x"5a",
         12018 => x"2e",
         12019 => x"77",
         12020 => x"84",
         12021 => x"5a",
         12022 => x"80",
         12023 => x"81",
         12024 => x"5d",
         12025 => x"08",
         12026 => x"ef",
         12027 => x"33",
         12028 => x"7c",
         12029 => x"81",
         12030 => x"b8",
         12031 => x"17",
         12032 => x"fd",
         12033 => x"bb",
         12034 => x"2e",
         12035 => x"5a",
         12036 => x"b4",
         12037 => x"7e",
         12038 => x"80",
         12039 => x"33",
         12040 => x"2e",
         12041 => x"77",
         12042 => x"83",
         12043 => x"12",
         12044 => x"2b",
         12045 => x"07",
         12046 => x"70",
         12047 => x"2b",
         12048 => x"80",
         12049 => x"80",
         12050 => x"30",
         12051 => x"63",
         12052 => x"05",
         12053 => x"62",
         12054 => x"41",
         12055 => x"52",
         12056 => x"5e",
         12057 => x"f2",
         12058 => x"0c",
         12059 => x"0c",
         12060 => x"81",
         12061 => x"84",
         12062 => x"84",
         12063 => x"95",
         12064 => x"81",
         12065 => x"08",
         12066 => x"70",
         12067 => x"33",
         12068 => x"fd",
         12069 => x"5e",
         12070 => x"08",
         12071 => x"84",
         12072 => x"83",
         12073 => x"17",
         12074 => x"08",
         12075 => x"84",
         12076 => x"74",
         12077 => x"27",
         12078 => x"82",
         12079 => x"74",
         12080 => x"81",
         12081 => x"38",
         12082 => x"17",
         12083 => x"08",
         12084 => x"52",
         12085 => x"51",
         12086 => x"3f",
         12087 => x"97",
         12088 => x"42",
         12089 => x"56",
         12090 => x"51",
         12091 => x"3f",
         12092 => x"08",
         12093 => x"e8",
         12094 => x"84",
         12095 => x"80",
         12096 => x"bb",
         12097 => x"70",
         12098 => x"08",
         12099 => x"7c",
         12100 => x"62",
         12101 => x"5c",
         12102 => x"76",
         12103 => x"7a",
         12104 => x"94",
         12105 => x"17",
         12106 => x"58",
         12107 => x"34",
         12108 => x"77",
         12109 => x"81",
         12110 => x"33",
         12111 => x"07",
         12112 => x"80",
         12113 => x"1d",
         12114 => x"ff",
         12115 => x"5f",
         12116 => x"55",
         12117 => x"38",
         12118 => x"77",
         12119 => x"39",
         12120 => x"5a",
         12121 => x"7a",
         12122 => x"84",
         12123 => x"07",
         12124 => x"18",
         12125 => x"39",
         12126 => x"5a",
         12127 => x"3d",
         12128 => x"89",
         12129 => x"2e",
         12130 => x"08",
         12131 => x"2e",
         12132 => x"33",
         12133 => x"2e",
         12134 => x"16",
         12135 => x"22",
         12136 => x"79",
         12137 => x"38",
         12138 => x"5b",
         12139 => x"38",
         12140 => x"57",
         12141 => x"38",
         12142 => x"70",
         12143 => x"06",
         12144 => x"56",
         12145 => x"80",
         12146 => x"18",
         12147 => x"8c",
         12148 => x"80",
         12149 => x"81",
         12150 => x"18",
         12151 => x"58",
         12152 => x"27",
         12153 => x"17",
         12154 => x"80",
         12155 => x"57",
         12156 => x"19",
         12157 => x"08",
         12158 => x"78",
         12159 => x"55",
         12160 => x"34",
         12161 => x"74",
         12162 => x"79",
         12163 => x"38",
         12164 => x"18",
         12165 => x"18",
         12166 => x"11",
         12167 => x"fe",
         12168 => x"84",
         12169 => x"80",
         12170 => x"38",
         12171 => x"91",
         12172 => x"56",
         12173 => x"84",
         12174 => x"0d",
         12175 => x"79",
         12176 => x"ff",
         12177 => x"77",
         12178 => x"94",
         12179 => x"84",
         12180 => x"bb",
         12181 => x"2e",
         12182 => x"84",
         12183 => x"81",
         12184 => x"38",
         12185 => x"08",
         12186 => x"f5",
         12187 => x"74",
         12188 => x"ff",
         12189 => x"84",
         12190 => x"82",
         12191 => x"17",
         12192 => x"94",
         12193 => x"56",
         12194 => x"27",
         12195 => x"81",
         12196 => x"0c",
         12197 => x"81",
         12198 => x"84",
         12199 => x"55",
         12200 => x"ff",
         12201 => x"39",
         12202 => x"51",
         12203 => x"3f",
         12204 => x"08",
         12205 => x"74",
         12206 => x"74",
         12207 => x"57",
         12208 => x"80",
         12209 => x"33",
         12210 => x"57",
         12211 => x"19",
         12212 => x"39",
         12213 => x"52",
         12214 => x"fe",
         12215 => x"bb",
         12216 => x"2e",
         12217 => x"84",
         12218 => x"81",
         12219 => x"38",
         12220 => x"38",
         12221 => x"bb",
         12222 => x"1a",
         12223 => x"a1",
         12224 => x"84",
         12225 => x"08",
         12226 => x"57",
         12227 => x"84",
         12228 => x"27",
         12229 => x"84",
         12230 => x"9c",
         12231 => x"81",
         12232 => x"80",
         12233 => x"ff",
         12234 => x"76",
         12235 => x"91",
         12236 => x"84",
         12237 => x"bb",
         12238 => x"e3",
         12239 => x"77",
         12240 => x"9c",
         12241 => x"84",
         12242 => x"bb",
         12243 => x"2e",
         12244 => x"84",
         12245 => x"81",
         12246 => x"38",
         12247 => x"08",
         12248 => x"8f",
         12249 => x"74",
         12250 => x"ff",
         12251 => x"84",
         12252 => x"80",
         12253 => x"17",
         12254 => x"94",
         12255 => x"56",
         12256 => x"27",
         12257 => x"16",
         12258 => x"84",
         12259 => x"07",
         12260 => x"18",
         12261 => x"78",
         12262 => x"a1",
         12263 => x"75",
         12264 => x"33",
         12265 => x"39",
         12266 => x"bb",
         12267 => x"90",
         12268 => x"57",
         12269 => x"82",
         12270 => x"90",
         12271 => x"ff",
         12272 => x"90",
         12273 => x"56",
         12274 => x"82",
         12275 => x"33",
         12276 => x"f6",
         12277 => x"84",
         12278 => x"33",
         12279 => x"ea",
         12280 => x"90",
         12281 => x"55",
         12282 => x"84",
         12283 => x"57",
         12284 => x"81",
         12285 => x"39",
         12286 => x"82",
         12287 => x"ff",
         12288 => x"a8",
         12289 => x"b8",
         12290 => x"bb",
         12291 => x"84",
         12292 => x"80",
         12293 => x"75",
         12294 => x"0c",
         12295 => x"04",
         12296 => x"3d",
         12297 => x"3d",
         12298 => x"ff",
         12299 => x"84",
         12300 => x"56",
         12301 => x"08",
         12302 => x"81",
         12303 => x"70",
         12304 => x"06",
         12305 => x"56",
         12306 => x"76",
         12307 => x"80",
         12308 => x"38",
         12309 => x"05",
         12310 => x"06",
         12311 => x"56",
         12312 => x"38",
         12313 => x"08",
         12314 => x"9a",
         12315 => x"88",
         12316 => x"33",
         12317 => x"57",
         12318 => x"2e",
         12319 => x"76",
         12320 => x"06",
         12321 => x"2e",
         12322 => x"87",
         12323 => x"08",
         12324 => x"83",
         12325 => x"7a",
         12326 => x"84",
         12327 => x"3d",
         12328 => x"ff",
         12329 => x"84",
         12330 => x"56",
         12331 => x"08",
         12332 => x"84",
         12333 => x"52",
         12334 => x"91",
         12335 => x"bb",
         12336 => x"84",
         12337 => x"a0",
         12338 => x"84",
         12339 => x"a7",
         12340 => x"95",
         12341 => x"17",
         12342 => x"2b",
         12343 => x"07",
         12344 => x"5d",
         12345 => x"39",
         12346 => x"08",
         12347 => x"38",
         12348 => x"08",
         12349 => x"78",
         12350 => x"3d",
         12351 => x"57",
         12352 => x"80",
         12353 => x"52",
         12354 => x"8b",
         12355 => x"bb",
         12356 => x"84",
         12357 => x"80",
         12358 => x"75",
         12359 => x"07",
         12360 => x"5a",
         12361 => x"9a",
         12362 => x"2e",
         12363 => x"79",
         12364 => x"81",
         12365 => x"38",
         12366 => x"7b",
         12367 => x"38",
         12368 => x"fd",
         12369 => x"51",
         12370 => x"3f",
         12371 => x"08",
         12372 => x"0c",
         12373 => x"04",
         12374 => x"98",
         12375 => x"80",
         12376 => x"08",
         12377 => x"b9",
         12378 => x"33",
         12379 => x"74",
         12380 => x"81",
         12381 => x"38",
         12382 => x"53",
         12383 => x"81",
         12384 => x"fe",
         12385 => x"84",
         12386 => x"80",
         12387 => x"ff",
         12388 => x"75",
         12389 => x"77",
         12390 => x"38",
         12391 => x"58",
         12392 => x"81",
         12393 => x"34",
         12394 => x"7c",
         12395 => x"38",
         12396 => x"51",
         12397 => x"3f",
         12398 => x"08",
         12399 => x"84",
         12400 => x"ff",
         12401 => x"84",
         12402 => x"06",
         12403 => x"82",
         12404 => x"39",
         12405 => x"17",
         12406 => x"52",
         12407 => x"51",
         12408 => x"3f",
         12409 => x"bb",
         12410 => x"2e",
         12411 => x"ff",
         12412 => x"bb",
         12413 => x"18",
         12414 => x"08",
         12415 => x"31",
         12416 => x"08",
         12417 => x"a0",
         12418 => x"fe",
         12419 => x"17",
         12420 => x"82",
         12421 => x"06",
         12422 => x"81",
         12423 => x"08",
         12424 => x"05",
         12425 => x"81",
         12426 => x"fe",
         12427 => x"79",
         12428 => x"39",
         12429 => x"78",
         12430 => x"38",
         12431 => x"51",
         12432 => x"3f",
         12433 => x"08",
         12434 => x"84",
         12435 => x"80",
         12436 => x"bb",
         12437 => x"2e",
         12438 => x"84",
         12439 => x"ff",
         12440 => x"38",
         12441 => x"52",
         12442 => x"fd",
         12443 => x"bb",
         12444 => x"38",
         12445 => x"fe",
         12446 => x"08",
         12447 => x"75",
         12448 => x"b0",
         12449 => x"94",
         12450 => x"17",
         12451 => x"5c",
         12452 => x"34",
         12453 => x"7a",
         12454 => x"38",
         12455 => x"a2",
         12456 => x"fd",
         12457 => x"bb",
         12458 => x"fd",
         12459 => x"56",
         12460 => x"e3",
         12461 => x"53",
         12462 => x"bc",
         12463 => x"3d",
         12464 => x"f9",
         12465 => x"84",
         12466 => x"bb",
         12467 => x"2e",
         12468 => x"84",
         12469 => x"9f",
         12470 => x"7d",
         12471 => x"93",
         12472 => x"5a",
         12473 => x"3f",
         12474 => x"08",
         12475 => x"84",
         12476 => x"88",
         12477 => x"84",
         12478 => x"0d",
         12479 => x"84",
         12480 => x"09",
         12481 => x"38",
         12482 => x"05",
         12483 => x"2a",
         12484 => x"58",
         12485 => x"ff",
         12486 => x"5f",
         12487 => x"3d",
         12488 => x"ff",
         12489 => x"84",
         12490 => x"75",
         12491 => x"bb",
         12492 => x"38",
         12493 => x"bb",
         12494 => x"2e",
         12495 => x"84",
         12496 => x"ff",
         12497 => x"38",
         12498 => x"38",
         12499 => x"84",
         12500 => x"33",
         12501 => x"7a",
         12502 => x"fe",
         12503 => x"08",
         12504 => x"56",
         12505 => x"79",
         12506 => x"8a",
         12507 => x"71",
         12508 => x"08",
         12509 => x"7a",
         12510 => x"b8",
         12511 => x"80",
         12512 => x"80",
         12513 => x"05",
         12514 => x"15",
         12515 => x"38",
         12516 => x"17",
         12517 => x"75",
         12518 => x"38",
         12519 => x"1b",
         12520 => x"81",
         12521 => x"fe",
         12522 => x"84",
         12523 => x"81",
         12524 => x"18",
         12525 => x"82",
         12526 => x"39",
         12527 => x"17",
         12528 => x"17",
         12529 => x"18",
         12530 => x"fe",
         12531 => x"81",
         12532 => x"84",
         12533 => x"84",
         12534 => x"83",
         12535 => x"17",
         12536 => x"08",
         12537 => x"a0",
         12538 => x"fe",
         12539 => x"17",
         12540 => x"82",
         12541 => x"06",
         12542 => x"75",
         12543 => x"08",
         12544 => x"05",
         12545 => x"81",
         12546 => x"fe",
         12547 => x"fe",
         12548 => x"56",
         12549 => x"58",
         12550 => x"27",
         12551 => x"7b",
         12552 => x"27",
         12553 => x"74",
         12554 => x"fe",
         12555 => x"84",
         12556 => x"5a",
         12557 => x"08",
         12558 => x"96",
         12559 => x"84",
         12560 => x"fd",
         12561 => x"bb",
         12562 => x"2e",
         12563 => x"80",
         12564 => x"76",
         12565 => x"e9",
         12566 => x"84",
         12567 => x"38",
         12568 => x"fe",
         12569 => x"08",
         12570 => x"77",
         12571 => x"38",
         12572 => x"18",
         12573 => x"33",
         12574 => x"7b",
         12575 => x"79",
         12576 => x"26",
         12577 => x"75",
         12578 => x"0c",
         12579 => x"04",
         12580 => x"55",
         12581 => x"ff",
         12582 => x"56",
         12583 => x"09",
         12584 => x"f0",
         12585 => x"b8",
         12586 => x"a0",
         12587 => x"05",
         12588 => x"16",
         12589 => x"38",
         12590 => x"0b",
         12591 => x"7d",
         12592 => x"80",
         12593 => x"7d",
         12594 => x"ce",
         12595 => x"80",
         12596 => x"a1",
         12597 => x"1a",
         12598 => x"0b",
         12599 => x"34",
         12600 => x"ff",
         12601 => x"56",
         12602 => x"17",
         12603 => x"2a",
         12604 => x"d3",
         12605 => x"33",
         12606 => x"2e",
         12607 => x"7d",
         12608 => x"80",
         12609 => x"1b",
         12610 => x"74",
         12611 => x"56",
         12612 => x"81",
         12613 => x"ff",
         12614 => x"ef",
         12615 => x"ae",
         12616 => x"17",
         12617 => x"71",
         12618 => x"06",
         12619 => x"78",
         12620 => x"34",
         12621 => x"5b",
         12622 => x"17",
         12623 => x"55",
         12624 => x"80",
         12625 => x"5b",
         12626 => x"1c",
         12627 => x"ff",
         12628 => x"84",
         12629 => x"56",
         12630 => x"08",
         12631 => x"69",
         12632 => x"84",
         12633 => x"34",
         12634 => x"08",
         12635 => x"a1",
         12636 => x"34",
         12637 => x"99",
         12638 => x"6a",
         12639 => x"9a",
         12640 => x"88",
         12641 => x"9b",
         12642 => x"33",
         12643 => x"2e",
         12644 => x"69",
         12645 => x"8b",
         12646 => x"57",
         12647 => x"18",
         12648 => x"fe",
         12649 => x"84",
         12650 => x"56",
         12651 => x"84",
         12652 => x"0d",
         12653 => x"2a",
         12654 => x"ec",
         12655 => x"88",
         12656 => x"80",
         12657 => x"fe",
         12658 => x"90",
         12659 => x"80",
         12660 => x"7a",
         12661 => x"74",
         12662 => x"34",
         12663 => x"0b",
         12664 => x"b8",
         12665 => x"56",
         12666 => x"7b",
         12667 => x"77",
         12668 => x"77",
         12669 => x"7b",
         12670 => x"69",
         12671 => x"8b",
         12672 => x"57",
         12673 => x"18",
         12674 => x"fe",
         12675 => x"84",
         12676 => x"56",
         12677 => x"d1",
         12678 => x"3d",
         12679 => x"70",
         12680 => x"79",
         12681 => x"38",
         12682 => x"05",
         12683 => x"9f",
         12684 => x"75",
         12685 => x"b8",
         12686 => x"38",
         12687 => x"81",
         12688 => x"53",
         12689 => x"fc",
         12690 => x"3d",
         12691 => x"ed",
         12692 => x"84",
         12693 => x"bb",
         12694 => x"2e",
         12695 => x"84",
         12696 => x"b1",
         12697 => x"7f",
         12698 => x"b2",
         12699 => x"a5",
         12700 => x"59",
         12701 => x"3f",
         12702 => x"08",
         12703 => x"84",
         12704 => x"02",
         12705 => x"33",
         12706 => x"5d",
         12707 => x"ce",
         12708 => x"92",
         12709 => x"08",
         12710 => x"75",
         12711 => x"57",
         12712 => x"81",
         12713 => x"ff",
         12714 => x"ef",
         12715 => x"58",
         12716 => x"58",
         12717 => x"70",
         12718 => x"33",
         12719 => x"05",
         12720 => x"15",
         12721 => x"38",
         12722 => x"52",
         12723 => x"9f",
         12724 => x"bb",
         12725 => x"84",
         12726 => x"85",
         12727 => x"a8",
         12728 => x"81",
         12729 => x"0b",
         12730 => x"0c",
         12731 => x"04",
         12732 => x"11",
         12733 => x"06",
         12734 => x"74",
         12735 => x"38",
         12736 => x"81",
         12737 => x"05",
         12738 => x"7a",
         12739 => x"38",
         12740 => x"83",
         12741 => x"08",
         12742 => x"5f",
         12743 => x"70",
         12744 => x"33",
         12745 => x"05",
         12746 => x"9f",
         12747 => x"56",
         12748 => x"89",
         12749 => x"70",
         12750 => x"57",
         12751 => x"17",
         12752 => x"26",
         12753 => x"17",
         12754 => x"06",
         12755 => x"30",
         12756 => x"59",
         12757 => x"2e",
         12758 => x"85",
         12759 => x"be",
         12760 => x"32",
         12761 => x"72",
         12762 => x"7a",
         12763 => x"55",
         12764 => x"95",
         12765 => x"84",
         12766 => x"7b",
         12767 => x"c2",
         12768 => x"7e",
         12769 => x"96",
         12770 => x"24",
         12771 => x"79",
         12772 => x"53",
         12773 => x"fc",
         12774 => x"3d",
         12775 => x"9d",
         12776 => x"84",
         12777 => x"bb",
         12778 => x"b2",
         12779 => x"39",
         12780 => x"08",
         12781 => x"06",
         12782 => x"77",
         12783 => x"e1",
         12784 => x"84",
         12785 => x"bb",
         12786 => x"92",
         12787 => x"93",
         12788 => x"02",
         12789 => x"cd",
         12790 => x"5a",
         12791 => x"05",
         12792 => x"70",
         12793 => x"34",
         12794 => x"79",
         12795 => x"80",
         12796 => x"8b",
         12797 => x"18",
         12798 => x"2a",
         12799 => x"56",
         12800 => x"75",
         12801 => x"76",
         12802 => x"7f",
         12803 => x"83",
         12804 => x"18",
         12805 => x"2a",
         12806 => x"5c",
         12807 => x"81",
         12808 => x"3d",
         12809 => x"81",
         12810 => x"9b",
         12811 => x"1a",
         12812 => x"2b",
         12813 => x"41",
         12814 => x"7d",
         12815 => x"e0",
         12816 => x"9c",
         12817 => x"05",
         12818 => x"7d",
         12819 => x"38",
         12820 => x"76",
         12821 => x"19",
         12822 => x"5e",
         12823 => x"82",
         12824 => x"7a",
         12825 => x"17",
         12826 => x"aa",
         12827 => x"33",
         12828 => x"bc",
         12829 => x"75",
         12830 => x"52",
         12831 => x"51",
         12832 => x"3f",
         12833 => x"08",
         12834 => x"38",
         12835 => x"5c",
         12836 => x"0c",
         12837 => x"80",
         12838 => x"56",
         12839 => x"38",
         12840 => x"5a",
         12841 => x"09",
         12842 => x"38",
         12843 => x"ff",
         12844 => x"56",
         12845 => x"18",
         12846 => x"2a",
         12847 => x"f3",
         12848 => x"33",
         12849 => x"2e",
         12850 => x"93",
         12851 => x"2a",
         12852 => x"ec",
         12853 => x"88",
         12854 => x"80",
         12855 => x"7f",
         12856 => x"83",
         12857 => x"08",
         12858 => x"b2",
         12859 => x"5c",
         12860 => x"2e",
         12861 => x"52",
         12862 => x"fb",
         12863 => x"bb",
         12864 => x"84",
         12865 => x"80",
         12866 => x"16",
         12867 => x"08",
         12868 => x"b4",
         12869 => x"2e",
         12870 => x"16",
         12871 => x"5f",
         12872 => x"09",
         12873 => x"a8",
         12874 => x"76",
         12875 => x"52",
         12876 => x"51",
         12877 => x"3f",
         12878 => x"08",
         12879 => x"38",
         12880 => x"58",
         12881 => x"0c",
         12882 => x"aa",
         12883 => x"08",
         12884 => x"34",
         12885 => x"17",
         12886 => x"08",
         12887 => x"38",
         12888 => x"51",
         12889 => x"3f",
         12890 => x"08",
         12891 => x"84",
         12892 => x"ff",
         12893 => x"56",
         12894 => x"f9",
         12895 => x"56",
         12896 => x"38",
         12897 => x"e5",
         12898 => x"bb",
         12899 => x"bb",
         12900 => x"3d",
         12901 => x"0b",
         12902 => x"0c",
         12903 => x"04",
         12904 => x"94",
         12905 => x"98",
         12906 => x"2b",
         12907 => x"58",
         12908 => x"8d",
         12909 => x"84",
         12910 => x"fb",
         12911 => x"bb",
         12912 => x"2e",
         12913 => x"75",
         12914 => x"0c",
         12915 => x"04",
         12916 => x"16",
         12917 => x"52",
         12918 => x"51",
         12919 => x"3f",
         12920 => x"bb",
         12921 => x"2e",
         12922 => x"fe",
         12923 => x"bb",
         12924 => x"17",
         12925 => x"08",
         12926 => x"31",
         12927 => x"08",
         12928 => x"a0",
         12929 => x"fe",
         12930 => x"16",
         12931 => x"82",
         12932 => x"06",
         12933 => x"81",
         12934 => x"08",
         12935 => x"05",
         12936 => x"81",
         12937 => x"fe",
         12938 => x"79",
         12939 => x"39",
         12940 => x"17",
         12941 => x"17",
         12942 => x"18",
         12943 => x"fe",
         12944 => x"81",
         12945 => x"84",
         12946 => x"38",
         12947 => x"08",
         12948 => x"b4",
         12949 => x"18",
         12950 => x"bb",
         12951 => x"55",
         12952 => x"08",
         12953 => x"38",
         12954 => x"5d",
         12955 => x"09",
         12956 => x"81",
         12957 => x"b4",
         12958 => x"18",
         12959 => x"7a",
         12960 => x"33",
         12961 => x"a4",
         12962 => x"fb",
         12963 => x"3d",
         12964 => x"df",
         12965 => x"84",
         12966 => x"05",
         12967 => x"82",
         12968 => x"cc",
         12969 => x"3d",
         12970 => x"91",
         12971 => x"84",
         12972 => x"bb",
         12973 => x"2e",
         12974 => x"84",
         12975 => x"96",
         12976 => x"78",
         12977 => x"96",
         12978 => x"51",
         12979 => x"3f",
         12980 => x"08",
         12981 => x"84",
         12982 => x"02",
         12983 => x"33",
         12984 => x"54",
         12985 => x"d2",
         12986 => x"06",
         12987 => x"8b",
         12988 => x"06",
         12989 => x"07",
         12990 => x"55",
         12991 => x"34",
         12992 => x"0b",
         12993 => x"78",
         12994 => x"d3",
         12995 => x"84",
         12996 => x"84",
         12997 => x"0d",
         12998 => x"0d",
         12999 => x"53",
         13000 => x"05",
         13001 => x"51",
         13002 => x"3f",
         13003 => x"08",
         13004 => x"84",
         13005 => x"8a",
         13006 => x"bb",
         13007 => x"3d",
         13008 => x"5a",
         13009 => x"3d",
         13010 => x"ff",
         13011 => x"84",
         13012 => x"55",
         13013 => x"08",
         13014 => x"80",
         13015 => x"81",
         13016 => x"86",
         13017 => x"38",
         13018 => x"22",
         13019 => x"71",
         13020 => x"59",
         13021 => x"96",
         13022 => x"88",
         13023 => x"97",
         13024 => x"90",
         13025 => x"98",
         13026 => x"98",
         13027 => x"99",
         13028 => x"57",
         13029 => x"18",
         13030 => x"fe",
         13031 => x"84",
         13032 => x"84",
         13033 => x"96",
         13034 => x"e8",
         13035 => x"6d",
         13036 => x"53",
         13037 => x"05",
         13038 => x"51",
         13039 => x"3f",
         13040 => x"08",
         13041 => x"08",
         13042 => x"bb",
         13043 => x"80",
         13044 => x"57",
         13045 => x"8b",
         13046 => x"76",
         13047 => x"78",
         13048 => x"76",
         13049 => x"07",
         13050 => x"5b",
         13051 => x"81",
         13052 => x"70",
         13053 => x"58",
         13054 => x"81",
         13055 => x"a4",
         13056 => x"56",
         13057 => x"16",
         13058 => x"82",
         13059 => x"16",
         13060 => x"55",
         13061 => x"09",
         13062 => x"98",
         13063 => x"76",
         13064 => x"52",
         13065 => x"51",
         13066 => x"3f",
         13067 => x"08",
         13068 => x"38",
         13069 => x"59",
         13070 => x"0c",
         13071 => x"bd",
         13072 => x"33",
         13073 => x"c3",
         13074 => x"2e",
         13075 => x"e4",
         13076 => x"2e",
         13077 => x"56",
         13078 => x"05",
         13079 => x"82",
         13080 => x"90",
         13081 => x"2b",
         13082 => x"33",
         13083 => x"88",
         13084 => x"71",
         13085 => x"5f",
         13086 => x"59",
         13087 => x"bb",
         13088 => x"3d",
         13089 => x"5e",
         13090 => x"52",
         13091 => x"52",
         13092 => x"c4",
         13093 => x"84",
         13094 => x"bb",
         13095 => x"2e",
         13096 => x"76",
         13097 => x"81",
         13098 => x"38",
         13099 => x"80",
         13100 => x"39",
         13101 => x"16",
         13102 => x"16",
         13103 => x"17",
         13104 => x"fe",
         13105 => x"77",
         13106 => x"84",
         13107 => x"09",
         13108 => x"e8",
         13109 => x"84",
         13110 => x"34",
         13111 => x"a8",
         13112 => x"84",
         13113 => x"5a",
         13114 => x"17",
         13115 => x"ad",
         13116 => x"33",
         13117 => x"2e",
         13118 => x"fe",
         13119 => x"54",
         13120 => x"a0",
         13121 => x"53",
         13122 => x"16",
         13123 => x"dc",
         13124 => x"59",
         13125 => x"53",
         13126 => x"81",
         13127 => x"fe",
         13128 => x"84",
         13129 => x"80",
         13130 => x"38",
         13131 => x"75",
         13132 => x"fe",
         13133 => x"84",
         13134 => x"57",
         13135 => x"08",
         13136 => x"84",
         13137 => x"84",
         13138 => x"66",
         13139 => x"79",
         13140 => x"7c",
         13141 => x"56",
         13142 => x"34",
         13143 => x"8a",
         13144 => x"38",
         13145 => x"57",
         13146 => x"34",
         13147 => x"fc",
         13148 => x"18",
         13149 => x"33",
         13150 => x"79",
         13151 => x"38",
         13152 => x"79",
         13153 => x"39",
         13154 => x"82",
         13155 => x"ff",
         13156 => x"a2",
         13157 => x"9d",
         13158 => x"bb",
         13159 => x"84",
         13160 => x"82",
         13161 => x"3d",
         13162 => x"57",
         13163 => x"70",
         13164 => x"34",
         13165 => x"74",
         13166 => x"a3",
         13167 => x"33",
         13168 => x"06",
         13169 => x"5a",
         13170 => x"81",
         13171 => x"3d",
         13172 => x"5c",
         13173 => x"06",
         13174 => x"55",
         13175 => x"38",
         13176 => x"74",
         13177 => x"26",
         13178 => x"74",
         13179 => x"3f",
         13180 => x"84",
         13181 => x"51",
         13182 => x"84",
         13183 => x"83",
         13184 => x"57",
         13185 => x"81",
         13186 => x"e8",
         13187 => x"e8",
         13188 => x"81",
         13189 => x"56",
         13190 => x"2e",
         13191 => x"74",
         13192 => x"2e",
         13193 => x"18",
         13194 => x"81",
         13195 => x"57",
         13196 => x"2e",
         13197 => x"77",
         13198 => x"06",
         13199 => x"81",
         13200 => x"78",
         13201 => x"81",
         13202 => x"81",
         13203 => x"89",
         13204 => x"38",
         13205 => x"27",
         13206 => x"88",
         13207 => x"7b",
         13208 => x"5d",
         13209 => x"5a",
         13210 => x"81",
         13211 => x"81",
         13212 => x"08",
         13213 => x"81",
         13214 => x"58",
         13215 => x"9f",
         13216 => x"38",
         13217 => x"57",
         13218 => x"81",
         13219 => x"38",
         13220 => x"99",
         13221 => x"05",
         13222 => x"70",
         13223 => x"7a",
         13224 => x"81",
         13225 => x"ff",
         13226 => x"ed",
         13227 => x"80",
         13228 => x"95",
         13229 => x"56",
         13230 => x"3f",
         13231 => x"08",
         13232 => x"84",
         13233 => x"b4",
         13234 => x"75",
         13235 => x"0c",
         13236 => x"04",
         13237 => x"74",
         13238 => x"3f",
         13239 => x"08",
         13240 => x"06",
         13241 => x"f8",
         13242 => x"75",
         13243 => x"0c",
         13244 => x"04",
         13245 => x"33",
         13246 => x"39",
         13247 => x"51",
         13248 => x"3f",
         13249 => x"08",
         13250 => x"84",
         13251 => x"38",
         13252 => x"82",
         13253 => x"6c",
         13254 => x"55",
         13255 => x"05",
         13256 => x"70",
         13257 => x"34",
         13258 => x"74",
         13259 => x"5d",
         13260 => x"1e",
         13261 => x"fe",
         13262 => x"84",
         13263 => x"55",
         13264 => x"87",
         13265 => x"27",
         13266 => x"86",
         13267 => x"39",
         13268 => x"08",
         13269 => x"81",
         13270 => x"38",
         13271 => x"75",
         13272 => x"38",
         13273 => x"53",
         13274 => x"fe",
         13275 => x"84",
         13276 => x"57",
         13277 => x"08",
         13278 => x"81",
         13279 => x"38",
         13280 => x"08",
         13281 => x"5a",
         13282 => x"57",
         13283 => x"18",
         13284 => x"b2",
         13285 => x"33",
         13286 => x"2e",
         13287 => x"81",
         13288 => x"54",
         13289 => x"18",
         13290 => x"33",
         13291 => x"fd",
         13292 => x"84",
         13293 => x"85",
         13294 => x"81",
         13295 => x"19",
         13296 => x"78",
         13297 => x"9c",
         13298 => x"33",
         13299 => x"74",
         13300 => x"81",
         13301 => x"30",
         13302 => x"78",
         13303 => x"74",
         13304 => x"d7",
         13305 => x"5a",
         13306 => x"a5",
         13307 => x"75",
         13308 => x"da",
         13309 => x"84",
         13310 => x"bb",
         13311 => x"2e",
         13312 => x"87",
         13313 => x"2e",
         13314 => x"76",
         13315 => x"b9",
         13316 => x"57",
         13317 => x"70",
         13318 => x"34",
         13319 => x"74",
         13320 => x"56",
         13321 => x"17",
         13322 => x"7e",
         13323 => x"76",
         13324 => x"58",
         13325 => x"81",
         13326 => x"ff",
         13327 => x"80",
         13328 => x"38",
         13329 => x"05",
         13330 => x"70",
         13331 => x"34",
         13332 => x"74",
         13333 => x"d6",
         13334 => x"e5",
         13335 => x"5d",
         13336 => x"1e",
         13337 => x"fe",
         13338 => x"84",
         13339 => x"55",
         13340 => x"81",
         13341 => x"39",
         13342 => x"18",
         13343 => x"52",
         13344 => x"51",
         13345 => x"3f",
         13346 => x"08",
         13347 => x"81",
         13348 => x"38",
         13349 => x"08",
         13350 => x"b4",
         13351 => x"19",
         13352 => x"7b",
         13353 => x"27",
         13354 => x"18",
         13355 => x"82",
         13356 => x"84",
         13357 => x"59",
         13358 => x"74",
         13359 => x"75",
         13360 => x"8a",
         13361 => x"84",
         13362 => x"bb",
         13363 => x"2e",
         13364 => x"fe",
         13365 => x"70",
         13366 => x"80",
         13367 => x"38",
         13368 => x"81",
         13369 => x"08",
         13370 => x"05",
         13371 => x"81",
         13372 => x"fe",
         13373 => x"fd",
         13374 => x"3d",
         13375 => x"02",
         13376 => x"cb",
         13377 => x"5b",
         13378 => x"76",
         13379 => x"38",
         13380 => x"74",
         13381 => x"38",
         13382 => x"73",
         13383 => x"38",
         13384 => x"84",
         13385 => x"59",
         13386 => x"81",
         13387 => x"54",
         13388 => x"81",
         13389 => x"17",
         13390 => x"81",
         13391 => x"80",
         13392 => x"38",
         13393 => x"81",
         13394 => x"17",
         13395 => x"2a",
         13396 => x"5d",
         13397 => x"81",
         13398 => x"8a",
         13399 => x"89",
         13400 => x"7c",
         13401 => x"59",
         13402 => x"3f",
         13403 => x"06",
         13404 => x"72",
         13405 => x"84",
         13406 => x"05",
         13407 => x"79",
         13408 => x"55",
         13409 => x"27",
         13410 => x"19",
         13411 => x"83",
         13412 => x"77",
         13413 => x"80",
         13414 => x"76",
         13415 => x"c0",
         13416 => x"7f",
         13417 => x"14",
         13418 => x"83",
         13419 => x"84",
         13420 => x"81",
         13421 => x"38",
         13422 => x"08",
         13423 => x"d8",
         13424 => x"84",
         13425 => x"38",
         13426 => x"78",
         13427 => x"38",
         13428 => x"09",
         13429 => x"38",
         13430 => x"54",
         13431 => x"84",
         13432 => x"0d",
         13433 => x"84",
         13434 => x"90",
         13435 => x"81",
         13436 => x"fe",
         13437 => x"84",
         13438 => x"81",
         13439 => x"fe",
         13440 => x"77",
         13441 => x"fe",
         13442 => x"80",
         13443 => x"38",
         13444 => x"58",
         13445 => x"ab",
         13446 => x"54",
         13447 => x"80",
         13448 => x"53",
         13449 => x"51",
         13450 => x"3f",
         13451 => x"08",
         13452 => x"84",
         13453 => x"38",
         13454 => x"ff",
         13455 => x"5e",
         13456 => x"7e",
         13457 => x"0c",
         13458 => x"2e",
         13459 => x"7a",
         13460 => x"79",
         13461 => x"90",
         13462 => x"c0",
         13463 => x"90",
         13464 => x"15",
         13465 => x"94",
         13466 => x"5a",
         13467 => x"fe",
         13468 => x"7d",
         13469 => x"0c",
         13470 => x"81",
         13471 => x"84",
         13472 => x"54",
         13473 => x"ff",
         13474 => x"39",
         13475 => x"59",
         13476 => x"82",
         13477 => x"39",
         13478 => x"c0",
         13479 => x"5e",
         13480 => x"84",
         13481 => x"e3",
         13482 => x"3d",
         13483 => x"08",
         13484 => x"81",
         13485 => x"44",
         13486 => x"0b",
         13487 => x"70",
         13488 => x"79",
         13489 => x"8a",
         13490 => x"81",
         13491 => x"70",
         13492 => x"56",
         13493 => x"85",
         13494 => x"ed",
         13495 => x"2e",
         13496 => x"84",
         13497 => x"56",
         13498 => x"84",
         13499 => x"10",
         13500 => x"cc",
         13501 => x"56",
         13502 => x"2e",
         13503 => x"75",
         13504 => x"84",
         13505 => x"33",
         13506 => x"12",
         13507 => x"5d",
         13508 => x"51",
         13509 => x"3f",
         13510 => x"08",
         13511 => x"70",
         13512 => x"56",
         13513 => x"84",
         13514 => x"82",
         13515 => x"40",
         13516 => x"84",
         13517 => x"3d",
         13518 => x"83",
         13519 => x"fe",
         13520 => x"84",
         13521 => x"84",
         13522 => x"55",
         13523 => x"84",
         13524 => x"82",
         13525 => x"84",
         13526 => x"15",
         13527 => x"74",
         13528 => x"7e",
         13529 => x"38",
         13530 => x"26",
         13531 => x"7e",
         13532 => x"26",
         13533 => x"ff",
         13534 => x"55",
         13535 => x"38",
         13536 => x"a6",
         13537 => x"2a",
         13538 => x"77",
         13539 => x"5b",
         13540 => x"85",
         13541 => x"30",
         13542 => x"77",
         13543 => x"91",
         13544 => x"b0",
         13545 => x"2e",
         13546 => x"81",
         13547 => x"60",
         13548 => x"fe",
         13549 => x"81",
         13550 => x"84",
         13551 => x"38",
         13552 => x"05",
         13553 => x"fe",
         13554 => x"88",
         13555 => x"56",
         13556 => x"82",
         13557 => x"09",
         13558 => x"f8",
         13559 => x"29",
         13560 => x"b2",
         13561 => x"58",
         13562 => x"82",
         13563 => x"b6",
         13564 => x"33",
         13565 => x"71",
         13566 => x"88",
         13567 => x"14",
         13568 => x"07",
         13569 => x"33",
         13570 => x"ba",
         13571 => x"33",
         13572 => x"71",
         13573 => x"88",
         13574 => x"14",
         13575 => x"07",
         13576 => x"33",
         13577 => x"a2",
         13578 => x"a3",
         13579 => x"3d",
         13580 => x"54",
         13581 => x"41",
         13582 => x"4d",
         13583 => x"ff",
         13584 => x"90",
         13585 => x"7a",
         13586 => x"82",
         13587 => x"81",
         13588 => x"06",
         13589 => x"80",
         13590 => x"38",
         13591 => x"45",
         13592 => x"89",
         13593 => x"06",
         13594 => x"f4",
         13595 => x"70",
         13596 => x"43",
         13597 => x"83",
         13598 => x"38",
         13599 => x"78",
         13600 => x"81",
         13601 => x"a8",
         13602 => x"74",
         13603 => x"38",
         13604 => x"98",
         13605 => x"a8",
         13606 => x"82",
         13607 => x"57",
         13608 => x"80",
         13609 => x"76",
         13610 => x"38",
         13611 => x"51",
         13612 => x"3f",
         13613 => x"08",
         13614 => x"55",
         13615 => x"08",
         13616 => x"96",
         13617 => x"84",
         13618 => x"10",
         13619 => x"08",
         13620 => x"72",
         13621 => x"57",
         13622 => x"ff",
         13623 => x"5d",
         13624 => x"47",
         13625 => x"11",
         13626 => x"11",
         13627 => x"6b",
         13628 => x"58",
         13629 => x"62",
         13630 => x"b8",
         13631 => x"5d",
         13632 => x"16",
         13633 => x"56",
         13634 => x"26",
         13635 => x"78",
         13636 => x"31",
         13637 => x"68",
         13638 => x"fc",
         13639 => x"84",
         13640 => x"40",
         13641 => x"89",
         13642 => x"82",
         13643 => x"06",
         13644 => x"83",
         13645 => x"84",
         13646 => x"27",
         13647 => x"7a",
         13648 => x"77",
         13649 => x"80",
         13650 => x"ef",
         13651 => x"fe",
         13652 => x"57",
         13653 => x"84",
         13654 => x"0d",
         13655 => x"0c",
         13656 => x"fb",
         13657 => x"0b",
         13658 => x"0c",
         13659 => x"84",
         13660 => x"04",
         13661 => x"11",
         13662 => x"06",
         13663 => x"74",
         13664 => x"38",
         13665 => x"81",
         13666 => x"05",
         13667 => x"7a",
         13668 => x"38",
         13669 => x"e6",
         13670 => x"7d",
         13671 => x"5b",
         13672 => x"05",
         13673 => x"70",
         13674 => x"33",
         13675 => x"45",
         13676 => x"99",
         13677 => x"e0",
         13678 => x"ff",
         13679 => x"ff",
         13680 => x"64",
         13681 => x"38",
         13682 => x"81",
         13683 => x"46",
         13684 => x"9f",
         13685 => x"76",
         13686 => x"81",
         13687 => x"78",
         13688 => x"75",
         13689 => x"30",
         13690 => x"9f",
         13691 => x"5d",
         13692 => x"80",
         13693 => x"38",
         13694 => x"1f",
         13695 => x"7c",
         13696 => x"38",
         13697 => x"e0",
         13698 => x"f8",
         13699 => x"52",
         13700 => x"cb",
         13701 => x"57",
         13702 => x"08",
         13703 => x"61",
         13704 => x"06",
         13705 => x"08",
         13706 => x"83",
         13707 => x"6c",
         13708 => x"7e",
         13709 => x"9c",
         13710 => x"31",
         13711 => x"39",
         13712 => x"d2",
         13713 => x"24",
         13714 => x"7b",
         13715 => x"0c",
         13716 => x"39",
         13717 => x"48",
         13718 => x"80",
         13719 => x"38",
         13720 => x"30",
         13721 => x"fc",
         13722 => x"bb",
         13723 => x"f5",
         13724 => x"7a",
         13725 => x"18",
         13726 => x"7b",
         13727 => x"38",
         13728 => x"84",
         13729 => x"9f",
         13730 => x"bb",
         13731 => x"80",
         13732 => x"2e",
         13733 => x"9f",
         13734 => x"8b",
         13735 => x"06",
         13736 => x"7a",
         13737 => x"84",
         13738 => x"55",
         13739 => x"81",
         13740 => x"ff",
         13741 => x"f4",
         13742 => x"83",
         13743 => x"57",
         13744 => x"81",
         13745 => x"76",
         13746 => x"58",
         13747 => x"55",
         13748 => x"60",
         13749 => x"74",
         13750 => x"61",
         13751 => x"77",
         13752 => x"34",
         13753 => x"ff",
         13754 => x"61",
         13755 => x"6a",
         13756 => x"7b",
         13757 => x"34",
         13758 => x"05",
         13759 => x"32",
         13760 => x"48",
         13761 => x"05",
         13762 => x"2a",
         13763 => x"68",
         13764 => x"34",
         13765 => x"83",
         13766 => x"86",
         13767 => x"83",
         13768 => x"55",
         13769 => x"05",
         13770 => x"2a",
         13771 => x"94",
         13772 => x"61",
         13773 => x"bf",
         13774 => x"34",
         13775 => x"05",
         13776 => x"9a",
         13777 => x"61",
         13778 => x"7e",
         13779 => x"34",
         13780 => x"48",
         13781 => x"05",
         13782 => x"2a",
         13783 => x"9e",
         13784 => x"98",
         13785 => x"90",
         13786 => x"90",
         13787 => x"05",
         13788 => x"2e",
         13789 => x"80",
         13790 => x"34",
         13791 => x"05",
         13792 => x"a9",
         13793 => x"cc",
         13794 => x"34",
         13795 => x"ff",
         13796 => x"61",
         13797 => x"74",
         13798 => x"6a",
         13799 => x"34",
         13800 => x"a4",
         13801 => x"61",
         13802 => x"93",
         13803 => x"83",
         13804 => x"57",
         13805 => x"81",
         13806 => x"76",
         13807 => x"58",
         13808 => x"55",
         13809 => x"60",
         13810 => x"49",
         13811 => x"34",
         13812 => x"05",
         13813 => x"6b",
         13814 => x"7e",
         13815 => x"79",
         13816 => x"c8",
         13817 => x"84",
         13818 => x"fa",
         13819 => x"17",
         13820 => x"2e",
         13821 => x"69",
         13822 => x"80",
         13823 => x"05",
         13824 => x"15",
         13825 => x"38",
         13826 => x"5b",
         13827 => x"86",
         13828 => x"ff",
         13829 => x"62",
         13830 => x"38",
         13831 => x"61",
         13832 => x"2a",
         13833 => x"74",
         13834 => x"05",
         13835 => x"90",
         13836 => x"64",
         13837 => x"46",
         13838 => x"2a",
         13839 => x"34",
         13840 => x"59",
         13841 => x"83",
         13842 => x"78",
         13843 => x"60",
         13844 => x"fe",
         13845 => x"84",
         13846 => x"85",
         13847 => x"80",
         13848 => x"80",
         13849 => x"05",
         13850 => x"15",
         13851 => x"38",
         13852 => x"7a",
         13853 => x"76",
         13854 => x"81",
         13855 => x"80",
         13856 => x"38",
         13857 => x"83",
         13858 => x"66",
         13859 => x"75",
         13860 => x"38",
         13861 => x"54",
         13862 => x"52",
         13863 => x"c5",
         13864 => x"bb",
         13865 => x"9b",
         13866 => x"76",
         13867 => x"5b",
         13868 => x"8c",
         13869 => x"2e",
         13870 => x"58",
         13871 => x"ff",
         13872 => x"84",
         13873 => x"2e",
         13874 => x"58",
         13875 => x"38",
         13876 => x"81",
         13877 => x"81",
         13878 => x"80",
         13879 => x"80",
         13880 => x"05",
         13881 => x"19",
         13882 => x"38",
         13883 => x"34",
         13884 => x"34",
         13885 => x"05",
         13886 => x"34",
         13887 => x"05",
         13888 => x"82",
         13889 => x"67",
         13890 => x"77",
         13891 => x"34",
         13892 => x"fd",
         13893 => x"1f",
         13894 => x"8b",
         13895 => x"85",
         13896 => x"bb",
         13897 => x"2a",
         13898 => x"76",
         13899 => x"34",
         13900 => x"08",
         13901 => x"34",
         13902 => x"c6",
         13903 => x"61",
         13904 => x"34",
         13905 => x"c8",
         13906 => x"bb",
         13907 => x"83",
         13908 => x"62",
         13909 => x"05",
         13910 => x"2a",
         13911 => x"83",
         13912 => x"62",
         13913 => x"77",
         13914 => x"05",
         13915 => x"2a",
         13916 => x"83",
         13917 => x"81",
         13918 => x"60",
         13919 => x"fe",
         13920 => x"81",
         13921 => x"84",
         13922 => x"38",
         13923 => x"52",
         13924 => x"c4",
         13925 => x"57",
         13926 => x"08",
         13927 => x"84",
         13928 => x"84",
         13929 => x"9f",
         13930 => x"bb",
         13931 => x"62",
         13932 => x"39",
         13933 => x"16",
         13934 => x"c4",
         13935 => x"38",
         13936 => x"57",
         13937 => x"e8",
         13938 => x"58",
         13939 => x"9d",
         13940 => x"26",
         13941 => x"e8",
         13942 => x"10",
         13943 => x"22",
         13944 => x"74",
         13945 => x"38",
         13946 => x"ee",
         13947 => x"78",
         13948 => x"b3",
         13949 => x"84",
         13950 => x"84",
         13951 => x"89",
         13952 => x"a0",
         13953 => x"84",
         13954 => x"fc",
         13955 => x"58",
         13956 => x"f0",
         13957 => x"f5",
         13958 => x"57",
         13959 => x"84",
         13960 => x"83",
         13961 => x"f8",
         13962 => x"f8",
         13963 => x"81",
         13964 => x"f4",
         13965 => x"57",
         13966 => x"68",
         13967 => x"63",
         13968 => x"af",
         13969 => x"f4",
         13970 => x"61",
         13971 => x"75",
         13972 => x"68",
         13973 => x"34",
         13974 => x"5b",
         13975 => x"05",
         13976 => x"2a",
         13977 => x"a3",
         13978 => x"c6",
         13979 => x"80",
         13980 => x"80",
         13981 => x"05",
         13982 => x"80",
         13983 => x"80",
         13984 => x"c6",
         13985 => x"61",
         13986 => x"7c",
         13987 => x"7b",
         13988 => x"34",
         13989 => x"59",
         13990 => x"05",
         13991 => x"2a",
         13992 => x"a7",
         13993 => x"61",
         13994 => x"80",
         13995 => x"34",
         13996 => x"05",
         13997 => x"af",
         13998 => x"61",
         13999 => x"80",
         14000 => x"34",
         14001 => x"05",
         14002 => x"b3",
         14003 => x"80",
         14004 => x"05",
         14005 => x"80",
         14006 => x"93",
         14007 => x"05",
         14008 => x"59",
         14009 => x"70",
         14010 => x"33",
         14011 => x"05",
         14012 => x"15",
         14013 => x"2e",
         14014 => x"76",
         14015 => x"58",
         14016 => x"81",
         14017 => x"ff",
         14018 => x"da",
         14019 => x"39",
         14020 => x"53",
         14021 => x"51",
         14022 => x"3f",
         14023 => x"bb",
         14024 => x"b0",
         14025 => x"29",
         14026 => x"77",
         14027 => x"05",
         14028 => x"84",
         14029 => x"53",
         14030 => x"51",
         14031 => x"3f",
         14032 => x"81",
         14033 => x"84",
         14034 => x"0d",
         14035 => x"0c",
         14036 => x"34",
         14037 => x"6a",
         14038 => x"4c",
         14039 => x"70",
         14040 => x"34",
         14041 => x"ff",
         14042 => x"34",
         14043 => x"05",
         14044 => x"86",
         14045 => x"61",
         14046 => x"ff",
         14047 => x"34",
         14048 => x"05",
         14049 => x"8a",
         14050 => x"65",
         14051 => x"f9",
         14052 => x"54",
         14053 => x"60",
         14054 => x"fe",
         14055 => x"84",
         14056 => x"57",
         14057 => x"81",
         14058 => x"ff",
         14059 => x"f4",
         14060 => x"80",
         14061 => x"81",
         14062 => x"7b",
         14063 => x"75",
         14064 => x"57",
         14065 => x"75",
         14066 => x"57",
         14067 => x"75",
         14068 => x"61",
         14069 => x"34",
         14070 => x"83",
         14071 => x"80",
         14072 => x"e6",
         14073 => x"e1",
         14074 => x"05",
         14075 => x"05",
         14076 => x"83",
         14077 => x"7a",
         14078 => x"78",
         14079 => x"05",
         14080 => x"2a",
         14081 => x"83",
         14082 => x"7a",
         14083 => x"7f",
         14084 => x"05",
         14085 => x"83",
         14086 => x"76",
         14087 => x"05",
         14088 => x"83",
         14089 => x"76",
         14090 => x"05",
         14091 => x"69",
         14092 => x"6b",
         14093 => x"87",
         14094 => x"52",
         14095 => x"bd",
         14096 => x"54",
         14097 => x"60",
         14098 => x"fe",
         14099 => x"69",
         14100 => x"f7",
         14101 => x"3d",
         14102 => x"5b",
         14103 => x"61",
         14104 => x"57",
         14105 => x"25",
         14106 => x"3d",
         14107 => x"f8",
         14108 => x"53",
         14109 => x"51",
         14110 => x"3f",
         14111 => x"09",
         14112 => x"38",
         14113 => x"55",
         14114 => x"90",
         14115 => x"70",
         14116 => x"34",
         14117 => x"74",
         14118 => x"38",
         14119 => x"cd",
         14120 => x"34",
         14121 => x"83",
         14122 => x"74",
         14123 => x"0c",
         14124 => x"04",
         14125 => x"7b",
         14126 => x"b3",
         14127 => x"57",
         14128 => x"80",
         14129 => x"17",
         14130 => x"76",
         14131 => x"88",
         14132 => x"17",
         14133 => x"59",
         14134 => x"81",
         14135 => x"bb",
         14136 => x"74",
         14137 => x"81",
         14138 => x"0c",
         14139 => x"04",
         14140 => x"05",
         14141 => x"8c",
         14142 => x"08",
         14143 => x"a7",
         14144 => x"32",
         14145 => x"72",
         14146 => x"70",
         14147 => x"0c",
         14148 => x"1b",
         14149 => x"56",
         14150 => x"52",
         14151 => x"94",
         14152 => x"39",
         14153 => x"02",
         14154 => x"33",
         14155 => x"58",
         14156 => x"57",
         14157 => x"70",
         14158 => x"34",
         14159 => x"74",
         14160 => x"3d",
         14161 => x"77",
         14162 => x"f7",
         14163 => x"80",
         14164 => x"c0",
         14165 => x"17",
         14166 => x"59",
         14167 => x"81",
         14168 => x"bb",
         14169 => x"74",
         14170 => x"81",
         14171 => x"0c",
         14172 => x"75",
         14173 => x"9f",
         14174 => x"11",
         14175 => x"c0",
         14176 => x"08",
         14177 => x"9f",
         14178 => x"84",
         14179 => x"7c",
         14180 => x"38",
         14181 => x"bb",
         14182 => x"3d",
         14183 => x"3d",
         14184 => x"55",
         14185 => x"05",
         14186 => x"51",
         14187 => x"3f",
         14188 => x"70",
         14189 => x"07",
         14190 => x"30",
         14191 => x"56",
         14192 => x"8d",
         14193 => x"fd",
         14194 => x"81",
         14195 => x"bb",
         14196 => x"3d",
         14197 => x"3d",
         14198 => x"84",
         14199 => x"22",
         14200 => x"52",
         14201 => x"26",
         14202 => x"83",
         14203 => x"52",
         14204 => x"84",
         14205 => x"0d",
         14206 => x"ff",
         14207 => x"70",
         14208 => x"09",
         14209 => x"38",
         14210 => x"e4",
         14211 => x"c8",
         14212 => x"71",
         14213 => x"81",
         14214 => x"ff",
         14215 => x"54",
         14216 => x"26",
         14217 => x"10",
         14218 => x"05",
         14219 => x"51",
         14220 => x"80",
         14221 => x"ff",
         14222 => x"84",
         14223 => x"3d",
         14224 => x"3d",
         14225 => x"05",
         14226 => x"05",
         14227 => x"53",
         14228 => x"70",
         14229 => x"8c",
         14230 => x"72",
         14231 => x"0c",
         14232 => x"04",
         14233 => x"2e",
         14234 => x"ef",
         14235 => x"ff",
         14236 => x"70",
         14237 => x"c8",
         14238 => x"84",
         14239 => x"51",
         14240 => x"04",
         14241 => x"77",
         14242 => x"ff",
         14243 => x"e1",
         14244 => x"ff",
         14245 => x"ea",
         14246 => x"75",
         14247 => x"80",
         14248 => x"70",
         14249 => x"22",
         14250 => x"70",
         14251 => x"7a",
         14252 => x"56",
         14253 => x"b7",
         14254 => x"82",
         14255 => x"72",
         14256 => x"54",
         14257 => x"06",
         14258 => x"54",
         14259 => x"b1",
         14260 => x"38",
         14261 => x"70",
         14262 => x"52",
         14263 => x"30",
         14264 => x"75",
         14265 => x"53",
         14266 => x"80",
         14267 => x"75",
         14268 => x"bb",
         14269 => x"3d",
         14270 => x"ee",
         14271 => x"a2",
         14272 => x"26",
         14273 => x"10",
         14274 => x"f0",
         14275 => x"08",
         14276 => x"16",
         14277 => x"ff",
         14278 => x"75",
         14279 => x"ff",
         14280 => x"83",
         14281 => x"57",
         14282 => x"88",
         14283 => x"ff",
         14284 => x"51",
         14285 => x"16",
         14286 => x"ff",
         14287 => x"db",
         14288 => x"70",
         14289 => x"06",
         14290 => x"39",
         14291 => x"83",
         14292 => x"57",
         14293 => x"f0",
         14294 => x"ff",
         14295 => x"51",
         14296 => x"75",
         14297 => x"06",
         14298 => x"70",
         14299 => x"06",
         14300 => x"ff",
         14301 => x"73",
         14302 => x"05",
         14303 => x"52",
         14304 => x"00",
         14305 => x"ff",
         14306 => x"00",
         14307 => x"ff",
         14308 => x"ff",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"00",
         14747 => x"00",
         14748 => x"00",
         14749 => x"00",
         14750 => x"00",
         14751 => x"00",
         14752 => x"00",
         14753 => x"00",
         14754 => x"00",
         14755 => x"00",
         14756 => x"00",
         14757 => x"00",
         14758 => x"00",
         14759 => x"00",
         14760 => x"00",
         14761 => x"00",
         14762 => x"00",
         14763 => x"00",
         14764 => x"00",
         14765 => x"00",
         14766 => x"00",
         14767 => x"00",
         14768 => x"00",
         14769 => x"00",
         14770 => x"00",
         14771 => x"00",
         14772 => x"00",
         14773 => x"00",
         14774 => x"00",
         14775 => x"00",
         14776 => x"00",
         14777 => x"00",
         14778 => x"00",
         14779 => x"00",
         14780 => x"00",
         14781 => x"00",
         14782 => x"69",
         14783 => x"00",
         14784 => x"69",
         14785 => x"6c",
         14786 => x"69",
         14787 => x"00",
         14788 => x"6c",
         14789 => x"00",
         14790 => x"65",
         14791 => x"00",
         14792 => x"63",
         14793 => x"72",
         14794 => x"63",
         14795 => x"00",
         14796 => x"64",
         14797 => x"00",
         14798 => x"64",
         14799 => x"00",
         14800 => x"65",
         14801 => x"65",
         14802 => x"65",
         14803 => x"69",
         14804 => x"69",
         14805 => x"66",
         14806 => x"66",
         14807 => x"61",
         14808 => x"00",
         14809 => x"6d",
         14810 => x"65",
         14811 => x"72",
         14812 => x"65",
         14813 => x"00",
         14814 => x"6e",
         14815 => x"00",
         14816 => x"65",
         14817 => x"00",
         14818 => x"6c",
         14819 => x"38",
         14820 => x"62",
         14821 => x"63",
         14822 => x"62",
         14823 => x"63",
         14824 => x"69",
         14825 => x"00",
         14826 => x"64",
         14827 => x"6e",
         14828 => x"77",
         14829 => x"72",
         14830 => x"2e",
         14831 => x"61",
         14832 => x"65",
         14833 => x"73",
         14834 => x"63",
         14835 => x"65",
         14836 => x"00",
         14837 => x"6f",
         14838 => x"61",
         14839 => x"6f",
         14840 => x"20",
         14841 => x"65",
         14842 => x"00",
         14843 => x"6e",
         14844 => x"66",
         14845 => x"65",
         14846 => x"6d",
         14847 => x"72",
         14848 => x"00",
         14849 => x"69",
         14850 => x"69",
         14851 => x"6f",
         14852 => x"64",
         14853 => x"69",
         14854 => x"75",
         14855 => x"6f",
         14856 => x"61",
         14857 => x"6e",
         14858 => x"6e",
         14859 => x"6c",
         14860 => x"00",
         14861 => x"6f",
         14862 => x"74",
         14863 => x"6f",
         14864 => x"64",
         14865 => x"6f",
         14866 => x"6d",
         14867 => x"69",
         14868 => x"20",
         14869 => x"65",
         14870 => x"74",
         14871 => x"66",
         14872 => x"64",
         14873 => x"20",
         14874 => x"6b",
         14875 => x"69",
         14876 => x"6e",
         14877 => x"65",
         14878 => x"6c",
         14879 => x"00",
         14880 => x"72",
         14881 => x"20",
         14882 => x"62",
         14883 => x"69",
         14884 => x"6e",
         14885 => x"69",
         14886 => x"00",
         14887 => x"44",
         14888 => x"20",
         14889 => x"74",
         14890 => x"72",
         14891 => x"63",
         14892 => x"2e",
         14893 => x"69",
         14894 => x"68",
         14895 => x"6c",
         14896 => x"6e",
         14897 => x"69",
         14898 => x"00",
         14899 => x"69",
         14900 => x"61",
         14901 => x"61",
         14902 => x"65",
         14903 => x"74",
         14904 => x"00",
         14905 => x"63",
         14906 => x"73",
         14907 => x"6e",
         14908 => x"2e",
         14909 => x"6e",
         14910 => x"69",
         14911 => x"69",
         14912 => x"61",
         14913 => x"00",
         14914 => x"6f",
         14915 => x"74",
         14916 => x"6f",
         14917 => x"2e",
         14918 => x"6f",
         14919 => x"6c",
         14920 => x"6f",
         14921 => x"2e",
         14922 => x"69",
         14923 => x"6e",
         14924 => x"72",
         14925 => x"79",
         14926 => x"6e",
         14927 => x"6e",
         14928 => x"65",
         14929 => x"72",
         14930 => x"69",
         14931 => x"45",
         14932 => x"72",
         14933 => x"75",
         14934 => x"73",
         14935 => x"00",
         14936 => x"25",
         14937 => x"62",
         14938 => x"73",
         14939 => x"20",
         14940 => x"25",
         14941 => x"62",
         14942 => x"73",
         14943 => x"63",
         14944 => x"00",
         14945 => x"65",
         14946 => x"00",
         14947 => x"30",
         14948 => x"00",
         14949 => x"20",
         14950 => x"30",
         14951 => x"00",
         14952 => x"7c",
         14953 => x"00",
         14954 => x"20",
         14955 => x"30",
         14956 => x"00",
         14957 => x"20",
         14958 => x"20",
         14959 => x"00",
         14960 => x"4f",
         14961 => x"2a",
         14962 => x"20",
         14963 => x"35",
         14964 => x"2f",
         14965 => x"31",
         14966 => x"31",
         14967 => x"00",
         14968 => x"5a",
         14969 => x"20",
         14970 => x"20",
         14971 => x"78",
         14972 => x"73",
         14973 => x"20",
         14974 => x"0a",
         14975 => x"53",
         14976 => x"20",
         14977 => x"61",
         14978 => x"41",
         14979 => x"65",
         14980 => x"20",
         14981 => x"20",
         14982 => x"20",
         14983 => x"3d",
         14984 => x"38",
         14985 => x"00",
         14986 => x"20",
         14987 => x"70",
         14988 => x"64",
         14989 => x"73",
         14990 => x"20",
         14991 => x"20",
         14992 => x"20",
         14993 => x"3d",
         14994 => x"38",
         14995 => x"00",
         14996 => x"50",
         14997 => x"6e",
         14998 => x"72",
         14999 => x"20",
         15000 => x"64",
         15001 => x"00",
         15002 => x"41",
         15003 => x"20",
         15004 => x"69",
         15005 => x"72",
         15006 => x"74",
         15007 => x"41",
         15008 => x"20",
         15009 => x"69",
         15010 => x"72",
         15011 => x"74",
         15012 => x"41",
         15013 => x"20",
         15014 => x"69",
         15015 => x"72",
         15016 => x"74",
         15017 => x"41",
         15018 => x"20",
         15019 => x"69",
         15020 => x"72",
         15021 => x"74",
         15022 => x"4f",
         15023 => x"20",
         15024 => x"69",
         15025 => x"72",
         15026 => x"74",
         15027 => x"4f",
         15028 => x"20",
         15029 => x"69",
         15030 => x"72",
         15031 => x"74",
         15032 => x"53",
         15033 => x"6e",
         15034 => x"72",
         15035 => x"00",
         15036 => x"69",
         15037 => x"20",
         15038 => x"65",
         15039 => x"70",
         15040 => x"65",
         15041 => x"6e",
         15042 => x"70",
         15043 => x"6d",
         15044 => x"2e",
         15045 => x"6e",
         15046 => x"69",
         15047 => x"74",
         15048 => x"72",
         15049 => x"00",
         15050 => x"75",
         15051 => x"78",
         15052 => x"62",
         15053 => x"00",
         15054 => x"4f",
         15055 => x"70",
         15056 => x"73",
         15057 => x"61",
         15058 => x"64",
         15059 => x"20",
         15060 => x"74",
         15061 => x"69",
         15062 => x"73",
         15063 => x"61",
         15064 => x"30",
         15065 => x"6c",
         15066 => x"65",
         15067 => x"69",
         15068 => x"61",
         15069 => x"6c",
         15070 => x"00",
         15071 => x"20",
         15072 => x"64",
         15073 => x"73",
         15074 => x"3a",
         15075 => x"61",
         15076 => x"6f",
         15077 => x"6e",
         15078 => x"00",
         15079 => x"50",
         15080 => x"69",
         15081 => x"64",
         15082 => x"73",
         15083 => x"2e",
         15084 => x"00",
         15085 => x"6f",
         15086 => x"72",
         15087 => x"6f",
         15088 => x"67",
         15089 => x"00",
         15090 => x"65",
         15091 => x"72",
         15092 => x"67",
         15093 => x"70",
         15094 => x"61",
         15095 => x"6e",
         15096 => x"00",
         15097 => x"61",
         15098 => x"6e",
         15099 => x"6f",
         15100 => x"40",
         15101 => x"38",
         15102 => x"2e",
         15103 => x"00",
         15104 => x"61",
         15105 => x"72",
         15106 => x"72",
         15107 => x"20",
         15108 => x"65",
         15109 => x"64",
         15110 => x"00",
         15111 => x"78",
         15112 => x"74",
         15113 => x"20",
         15114 => x"65",
         15115 => x"25",
         15116 => x"78",
         15117 => x"2e",
         15118 => x"30",
         15119 => x"20",
         15120 => x"6c",
         15121 => x"00",
         15122 => x"30",
         15123 => x"20",
         15124 => x"58",
         15125 => x"6f",
         15126 => x"72",
         15127 => x"2e",
         15128 => x"00",
         15129 => x"30",
         15130 => x"28",
         15131 => x"78",
         15132 => x"25",
         15133 => x"78",
         15134 => x"38",
         15135 => x"00",
         15136 => x"6f",
         15137 => x"6e",
         15138 => x"2e",
         15139 => x"30",
         15140 => x"20",
         15141 => x"58",
         15142 => x"6c",
         15143 => x"69",
         15144 => x"2e",
         15145 => x"00",
         15146 => x"75",
         15147 => x"4d",
         15148 => x"72",
         15149 => x"43",
         15150 => x"6c",
         15151 => x"2e",
         15152 => x"64",
         15153 => x"73",
         15154 => x"00",
         15155 => x"65",
         15156 => x"79",
         15157 => x"68",
         15158 => x"74",
         15159 => x"20",
         15160 => x"6e",
         15161 => x"70",
         15162 => x"65",
         15163 => x"63",
         15164 => x"61",
         15165 => x"00",
         15166 => x"3f",
         15167 => x"64",
         15168 => x"2f",
         15169 => x"25",
         15170 => x"64",
         15171 => x"2e",
         15172 => x"64",
         15173 => x"6f",
         15174 => x"6f",
         15175 => x"67",
         15176 => x"74",
         15177 => x"00",
         15178 => x"0a",
         15179 => x"69",
         15180 => x"20",
         15181 => x"6c",
         15182 => x"6e",
         15183 => x"3a",
         15184 => x"64",
         15185 => x"73",
         15186 => x"3a",
         15187 => x"20",
         15188 => x"50",
         15189 => x"65",
         15190 => x"20",
         15191 => x"74",
         15192 => x"41",
         15193 => x"65",
         15194 => x"3d",
         15195 => x"38",
         15196 => x"00",
         15197 => x"20",
         15198 => x"50",
         15199 => x"65",
         15200 => x"79",
         15201 => x"61",
         15202 => x"41",
         15203 => x"65",
         15204 => x"3d",
         15205 => x"38",
         15206 => x"00",
         15207 => x"20",
         15208 => x"74",
         15209 => x"20",
         15210 => x"72",
         15211 => x"64",
         15212 => x"73",
         15213 => x"20",
         15214 => x"3d",
         15215 => x"38",
         15216 => x"00",
         15217 => x"69",
         15218 => x"00",
         15219 => x"20",
         15220 => x"50",
         15221 => x"64",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"20",
         15226 => x"3d",
         15227 => x"34",
         15228 => x"00",
         15229 => x"20",
         15230 => x"79",
         15231 => x"6d",
         15232 => x"6f",
         15233 => x"46",
         15234 => x"20",
         15235 => x"20",
         15236 => x"3d",
         15237 => x"2e",
         15238 => x"64",
         15239 => x"0a",
         15240 => x"20",
         15241 => x"69",
         15242 => x"6f",
         15243 => x"53",
         15244 => x"4d",
         15245 => x"6f",
         15246 => x"46",
         15247 => x"3d",
         15248 => x"2e",
         15249 => x"64",
         15250 => x"0a",
         15251 => x"20",
         15252 => x"44",
         15253 => x"20",
         15254 => x"63",
         15255 => x"72",
         15256 => x"20",
         15257 => x"20",
         15258 => x"3d",
         15259 => x"2e",
         15260 => x"64",
         15261 => x"0a",
         15262 => x"20",
         15263 => x"50",
         15264 => x"20",
         15265 => x"53",
         15266 => x"20",
         15267 => x"4f",
         15268 => x"00",
         15269 => x"20",
         15270 => x"42",
         15271 => x"43",
         15272 => x"20",
         15273 => x"49",
         15274 => x"4f",
         15275 => x"42",
         15276 => x"00",
         15277 => x"20",
         15278 => x"4e",
         15279 => x"43",
         15280 => x"20",
         15281 => x"61",
         15282 => x"6c",
         15283 => x"30",
         15284 => x"2e",
         15285 => x"20",
         15286 => x"49",
         15287 => x"31",
         15288 => x"20",
         15289 => x"6d",
         15290 => x"20",
         15291 => x"30",
         15292 => x"2e",
         15293 => x"20",
         15294 => x"44",
         15295 => x"52",
         15296 => x"20",
         15297 => x"76",
         15298 => x"73",
         15299 => x"30",
         15300 => x"2e",
         15301 => x"20",
         15302 => x"41",
         15303 => x"20",
         15304 => x"20",
         15305 => x"38",
         15306 => x"30",
         15307 => x"2e",
         15308 => x"20",
         15309 => x"52",
         15310 => x"20",
         15311 => x"20",
         15312 => x"38",
         15313 => x"30",
         15314 => x"2e",
         15315 => x"20",
         15316 => x"4e",
         15317 => x"42",
         15318 => x"20",
         15319 => x"38",
         15320 => x"30",
         15321 => x"2e",
         15322 => x"20",
         15323 => x"44",
         15324 => x"20",
         15325 => x"20",
         15326 => x"38",
         15327 => x"30",
         15328 => x"2e",
         15329 => x"20",
         15330 => x"42",
         15331 => x"52",
         15332 => x"20",
         15333 => x"38",
         15334 => x"30",
         15335 => x"2e",
         15336 => x"28",
         15337 => x"6d",
         15338 => x"43",
         15339 => x"6e",
         15340 => x"29",
         15341 => x"6e",
         15342 => x"77",
         15343 => x"56",
         15344 => x"00",
         15345 => x"6d",
         15346 => x"00",
         15347 => x"65",
         15348 => x"6d",
         15349 => x"6c",
         15350 => x"00",
         15351 => x"56",
         15352 => x"00",
         15353 => x"00",
         15354 => x"00",
         15355 => x"00",
         15356 => x"00",
         15357 => x"00",
         15358 => x"00",
         15359 => x"00",
         15360 => x"00",
         15361 => x"00",
         15362 => x"00",
         15363 => x"00",
         15364 => x"00",
         15365 => x"00",
         15366 => x"00",
         15367 => x"00",
         15368 => x"00",
         15369 => x"00",
         15370 => x"00",
         15371 => x"00",
         15372 => x"00",
         15373 => x"00",
         15374 => x"00",
         15375 => x"00",
         15376 => x"00",
         15377 => x"00",
         15378 => x"00",
         15379 => x"00",
         15380 => x"00",
         15381 => x"00",
         15382 => x"00",
         15383 => x"00",
         15384 => x"00",
         15385 => x"00",
         15386 => x"00",
         15387 => x"00",
         15388 => x"00",
         15389 => x"00",
         15390 => x"00",
         15391 => x"00",
         15392 => x"00",
         15393 => x"00",
         15394 => x"00",
         15395 => x"00",
         15396 => x"00",
         15397 => x"00",
         15398 => x"00",
         15399 => x"00",
         15400 => x"00",
         15401 => x"00",
         15402 => x"00",
         15403 => x"00",
         15404 => x"00",
         15405 => x"00",
         15406 => x"00",
         15407 => x"00",
         15408 => x"00",
         15409 => x"00",
         15410 => x"00",
         15411 => x"00",
         15412 => x"00",
         15413 => x"00",
         15414 => x"00",
         15415 => x"00",
         15416 => x"00",
         15417 => x"00",
         15418 => x"5b",
         15419 => x"5b",
         15420 => x"5b",
         15421 => x"5b",
         15422 => x"5b",
         15423 => x"5b",
         15424 => x"5b",
         15425 => x"30",
         15426 => x"5b",
         15427 => x"5b",
         15428 => x"5b",
         15429 => x"00",
         15430 => x"00",
         15431 => x"00",
         15432 => x"00",
         15433 => x"00",
         15434 => x"00",
         15435 => x"00",
         15436 => x"00",
         15437 => x"00",
         15438 => x"00",
         15439 => x"00",
         15440 => x"69",
         15441 => x"72",
         15442 => x"65",
         15443 => x"25",
         15444 => x"78",
         15445 => x"61",
         15446 => x"74",
         15447 => x"65",
         15448 => x"72",
         15449 => x"65",
         15450 => x"73",
         15451 => x"79",
         15452 => x"6c",
         15453 => x"64",
         15454 => x"62",
         15455 => x"67",
         15456 => x"69",
         15457 => x"72",
         15458 => x"69",
         15459 => x"00",
         15460 => x"00",
         15461 => x"69",
         15462 => x"72",
         15463 => x"75",
         15464 => x"72",
         15465 => x"38",
         15466 => x"00",
         15467 => x"30",
         15468 => x"20",
         15469 => x"0a",
         15470 => x"61",
         15471 => x"64",
         15472 => x"20",
         15473 => x"65",
         15474 => x"68",
         15475 => x"69",
         15476 => x"72",
         15477 => x"69",
         15478 => x"74",
         15479 => x"4f",
         15480 => x"00",
         15481 => x"25",
         15482 => x"00",
         15483 => x"5b",
         15484 => x"00",
         15485 => x"5b",
         15486 => x"5b",
         15487 => x"5b",
         15488 => x"5b",
         15489 => x"5b",
         15490 => x"00",
         15491 => x"5b",
         15492 => x"00",
         15493 => x"5b",
         15494 => x"00",
         15495 => x"5b",
         15496 => x"00",
         15497 => x"5b",
         15498 => x"00",
         15499 => x"5b",
         15500 => x"00",
         15501 => x"5b",
         15502 => x"00",
         15503 => x"5b",
         15504 => x"00",
         15505 => x"5b",
         15506 => x"00",
         15507 => x"5b",
         15508 => x"00",
         15509 => x"5b",
         15510 => x"00",
         15511 => x"5b",
         15512 => x"00",
         15513 => x"5b",
         15514 => x"5b",
         15515 => x"00",
         15516 => x"5b",
         15517 => x"00",
         15518 => x"3a",
         15519 => x"25",
         15520 => x"64",
         15521 => x"2c",
         15522 => x"25",
         15523 => x"30",
         15524 => x"00",
         15525 => x"3a",
         15526 => x"25",
         15527 => x"64",
         15528 => x"3a",
         15529 => x"25",
         15530 => x"64",
         15531 => x"64",
         15532 => x"3a",
         15533 => x"00",
         15534 => x"30",
         15535 => x"00",
         15536 => x"63",
         15537 => x"3b",
         15538 => x"00",
         15539 => x"65",
         15540 => x"74",
         15541 => x"72",
         15542 => x"3a",
         15543 => x"70",
         15544 => x"32",
         15545 => x"30",
         15546 => x"00",
         15547 => x"77",
         15548 => x"32",
         15549 => x"30",
         15550 => x"00",
         15551 => x"64",
         15552 => x"32",
         15553 => x"00",
         15554 => x"6f",
         15555 => x"73",
         15556 => x"65",
         15557 => x"65",
         15558 => x"00",
         15559 => x"44",
         15560 => x"2a",
         15561 => x"3f",
         15562 => x"00",
         15563 => x"2c",
         15564 => x"5d",
         15565 => x"41",
         15566 => x"41",
         15567 => x"00",
         15568 => x"fe",
         15569 => x"44",
         15570 => x"2e",
         15571 => x"4f",
         15572 => x"4d",
         15573 => x"20",
         15574 => x"54",
         15575 => x"20",
         15576 => x"4f",
         15577 => x"4d",
         15578 => x"20",
         15579 => x"54",
         15580 => x"20",
         15581 => x"00",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"03",
         15586 => x"0e",
         15587 => x"16",
         15588 => x"00",
         15589 => x"9a",
         15590 => x"41",
         15591 => x"45",
         15592 => x"49",
         15593 => x"92",
         15594 => x"4f",
         15595 => x"99",
         15596 => x"9d",
         15597 => x"49",
         15598 => x"a5",
         15599 => x"a9",
         15600 => x"ad",
         15601 => x"b1",
         15602 => x"b5",
         15603 => x"b9",
         15604 => x"bd",
         15605 => x"c1",
         15606 => x"c5",
         15607 => x"c9",
         15608 => x"cd",
         15609 => x"d1",
         15610 => x"d5",
         15611 => x"d9",
         15612 => x"dd",
         15613 => x"e1",
         15614 => x"e5",
         15615 => x"e9",
         15616 => x"ed",
         15617 => x"f1",
         15618 => x"f5",
         15619 => x"f9",
         15620 => x"fd",
         15621 => x"2e",
         15622 => x"5b",
         15623 => x"22",
         15624 => x"3e",
         15625 => x"00",
         15626 => x"01",
         15627 => x"10",
         15628 => x"00",
         15629 => x"00",
         15630 => x"01",
         15631 => x"04",
         15632 => x"10",
         15633 => x"00",
         15634 => x"c7",
         15635 => x"e9",
         15636 => x"e4",
         15637 => x"e5",
         15638 => x"ea",
         15639 => x"e8",
         15640 => x"ee",
         15641 => x"c4",
         15642 => x"c9",
         15643 => x"c6",
         15644 => x"f6",
         15645 => x"fb",
         15646 => x"ff",
         15647 => x"dc",
         15648 => x"a3",
         15649 => x"a7",
         15650 => x"e1",
         15651 => x"f3",
         15652 => x"f1",
         15653 => x"aa",
         15654 => x"bf",
         15655 => x"ac",
         15656 => x"bc",
         15657 => x"ab",
         15658 => x"91",
         15659 => x"93",
         15660 => x"24",
         15661 => x"62",
         15662 => x"55",
         15663 => x"51",
         15664 => x"5d",
         15665 => x"5b",
         15666 => x"14",
         15667 => x"2c",
         15668 => x"00",
         15669 => x"5e",
         15670 => x"5a",
         15671 => x"69",
         15672 => x"60",
         15673 => x"6c",
         15674 => x"68",
         15675 => x"65",
         15676 => x"58",
         15677 => x"53",
         15678 => x"6a",
         15679 => x"0c",
         15680 => x"84",
         15681 => x"90",
         15682 => x"b1",
         15683 => x"93",
         15684 => x"a3",
         15685 => x"b5",
         15686 => x"a6",
         15687 => x"a9",
         15688 => x"1e",
         15689 => x"b5",
         15690 => x"61",
         15691 => x"65",
         15692 => x"20",
         15693 => x"f7",
         15694 => x"b0",
         15695 => x"b7",
         15696 => x"7f",
         15697 => x"a0",
         15698 => x"61",
         15699 => x"e0",
         15700 => x"f8",
         15701 => x"ff",
         15702 => x"78",
         15703 => x"30",
         15704 => x"06",
         15705 => x"10",
         15706 => x"2e",
         15707 => x"06",
         15708 => x"4d",
         15709 => x"81",
         15710 => x"82",
         15711 => x"84",
         15712 => x"87",
         15713 => x"89",
         15714 => x"8b",
         15715 => x"8d",
         15716 => x"8f",
         15717 => x"91",
         15718 => x"93",
         15719 => x"f6",
         15720 => x"97",
         15721 => x"98",
         15722 => x"9b",
         15723 => x"9d",
         15724 => x"9f",
         15725 => x"a0",
         15726 => x"a2",
         15727 => x"a4",
         15728 => x"a7",
         15729 => x"a9",
         15730 => x"ab",
         15731 => x"ac",
         15732 => x"af",
         15733 => x"b1",
         15734 => x"b3",
         15735 => x"b5",
         15736 => x"b7",
         15737 => x"b8",
         15738 => x"bb",
         15739 => x"bc",
         15740 => x"f7",
         15741 => x"c1",
         15742 => x"c3",
         15743 => x"c5",
         15744 => x"c7",
         15745 => x"c7",
         15746 => x"cb",
         15747 => x"cd",
         15748 => x"dd",
         15749 => x"8e",
         15750 => x"12",
         15751 => x"03",
         15752 => x"f4",
         15753 => x"f8",
         15754 => x"22",
         15755 => x"3a",
         15756 => x"65",
         15757 => x"3b",
         15758 => x"66",
         15759 => x"40",
         15760 => x"41",
         15761 => x"0a",
         15762 => x"40",
         15763 => x"86",
         15764 => x"89",
         15765 => x"58",
         15766 => x"5a",
         15767 => x"5c",
         15768 => x"5e",
         15769 => x"93",
         15770 => x"62",
         15771 => x"64",
         15772 => x"66",
         15773 => x"97",
         15774 => x"6a",
         15775 => x"6c",
         15776 => x"6e",
         15777 => x"70",
         15778 => x"9d",
         15779 => x"74",
         15780 => x"76",
         15781 => x"78",
         15782 => x"7a",
         15783 => x"7c",
         15784 => x"7e",
         15785 => x"a6",
         15786 => x"82",
         15787 => x"84",
         15788 => x"86",
         15789 => x"ae",
         15790 => x"b1",
         15791 => x"45",
         15792 => x"8e",
         15793 => x"90",
         15794 => x"b7",
         15795 => x"03",
         15796 => x"fe",
         15797 => x"ac",
         15798 => x"86",
         15799 => x"89",
         15800 => x"b1",
         15801 => x"c2",
         15802 => x"a3",
         15803 => x"c4",
         15804 => x"cc",
         15805 => x"8c",
         15806 => x"8f",
         15807 => x"18",
         15808 => x"0a",
         15809 => x"f3",
         15810 => x"f5",
         15811 => x"f7",
         15812 => x"f9",
         15813 => x"fa",
         15814 => x"20",
         15815 => x"10",
         15816 => x"22",
         15817 => x"36",
         15818 => x"0e",
         15819 => x"01",
         15820 => x"d0",
         15821 => x"61",
         15822 => x"00",
         15823 => x"7d",
         15824 => x"63",
         15825 => x"96",
         15826 => x"5a",
         15827 => x"08",
         15828 => x"06",
         15829 => x"08",
         15830 => x"08",
         15831 => x"06",
         15832 => x"07",
         15833 => x"52",
         15834 => x"54",
         15835 => x"56",
         15836 => x"60",
         15837 => x"70",
         15838 => x"ba",
         15839 => x"c8",
         15840 => x"ca",
         15841 => x"da",
         15842 => x"f8",
         15843 => x"ea",
         15844 => x"fa",
         15845 => x"80",
         15846 => x"90",
         15847 => x"a0",
         15848 => x"b0",
         15849 => x"b8",
         15850 => x"b2",
         15851 => x"cc",
         15852 => x"c3",
         15853 => x"02",
         15854 => x"02",
         15855 => x"01",
         15856 => x"f3",
         15857 => x"fc",
         15858 => x"01",
         15859 => x"70",
         15860 => x"84",
         15861 => x"83",
         15862 => x"1a",
         15863 => x"2f",
         15864 => x"02",
         15865 => x"06",
         15866 => x"02",
         15867 => x"64",
         15868 => x"26",
         15869 => x"1a",
         15870 => x"00",
         15871 => x"00",
         15872 => x"02",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"04",
         15877 => x"00",
         15878 => x"00",
         15879 => x"00",
         15880 => x"14",
         15881 => x"00",
         15882 => x"00",
         15883 => x"00",
         15884 => x"2b",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"30",
         15889 => x"00",
         15890 => x"00",
         15891 => x"00",
         15892 => x"3c",
         15893 => x"00",
         15894 => x"00",
         15895 => x"00",
         15896 => x"3d",
         15897 => x"00",
         15898 => x"00",
         15899 => x"00",
         15900 => x"3f",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"40",
         15905 => x"00",
         15906 => x"00",
         15907 => x"00",
         15908 => x"41",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"42",
         15913 => x"00",
         15914 => x"00",
         15915 => x"00",
         15916 => x"43",
         15917 => x"00",
         15918 => x"00",
         15919 => x"00",
         15920 => x"50",
         15921 => x"00",
         15922 => x"00",
         15923 => x"00",
         15924 => x"51",
         15925 => x"00",
         15926 => x"00",
         15927 => x"00",
         15928 => x"54",
         15929 => x"00",
         15930 => x"00",
         15931 => x"00",
         15932 => x"55",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"79",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"78",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"82",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"83",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"85",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"87",
         15957 => x"00",
         15958 => x"00",
         15959 => x"00",
         15960 => x"88",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"89",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"8c",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"8d",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"8e",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"8f",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"01",
         15989 => x"00",
         15990 => x"01",
         15991 => x"81",
         15992 => x"00",
         15993 => x"7f",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"f5",
         15999 => x"f5",
         16000 => x"f5",
         16001 => x"00",
         16002 => x"01",
         16003 => x"01",
         16004 => x"01",
         16005 => x"00",
         16006 => x"00",
         16007 => x"00",
         16008 => x"00",
         16009 => x"00",
         16010 => x"00",
         16011 => x"00",
         16012 => x"00",
         16013 => x"00",
         16014 => x"00",
         16015 => x"00",
         16016 => x"00",
         16017 => x"00",
         16018 => x"00",
         16019 => x"00",
         16020 => x"00",
         16021 => x"00",
         16022 => x"00",
         16023 => x"00",
         16024 => x"00",
         16025 => x"00",
         16026 => x"00",
         16027 => x"00",
         16028 => x"00",
         16029 => x"00",
         16030 => x"00",
         16031 => x"00",
         16032 => x"00",
         16033 => x"00",
         16034 => x"00",
         16035 => x"00",
         16036 => x"01",
         16037 => x"fc",
         16038 => x"3b",
         16039 => x"7a",
         16040 => x"f0",
         16041 => x"72",
         16042 => x"76",
         16043 => x"6a",
         16044 => x"6e",
         16045 => x"62",
         16046 => x"66",
         16047 => x"32",
         16048 => x"36",
         16049 => x"f3",
         16050 => x"39",
         16051 => x"7f",
         16052 => x"f2",
         16053 => x"f0",
         16054 => x"f0",
         16055 => x"81",
         16056 => x"f0",
         16057 => x"fc",
         16058 => x"3a",
         16059 => x"5a",
         16060 => x"f0",
         16061 => x"52",
         16062 => x"56",
         16063 => x"4a",
         16064 => x"4e",
         16065 => x"42",
         16066 => x"46",
         16067 => x"32",
         16068 => x"36",
         16069 => x"f3",
         16070 => x"39",
         16071 => x"7f",
         16072 => x"f2",
         16073 => x"f0",
         16074 => x"f0",
         16075 => x"81",
         16076 => x"f0",
         16077 => x"fc",
         16078 => x"2b",
         16079 => x"5a",
         16080 => x"f0",
         16081 => x"52",
         16082 => x"56",
         16083 => x"4a",
         16084 => x"4e",
         16085 => x"42",
         16086 => x"46",
         16087 => x"22",
         16088 => x"26",
         16089 => x"7e",
         16090 => x"29",
         16091 => x"e2",
         16092 => x"f8",
         16093 => x"f0",
         16094 => x"f0",
         16095 => x"86",
         16096 => x"f0",
         16097 => x"fe",
         16098 => x"f0",
         16099 => x"1a",
         16100 => x"f0",
         16101 => x"12",
         16102 => x"16",
         16103 => x"0a",
         16104 => x"0e",
         16105 => x"02",
         16106 => x"06",
         16107 => x"f0",
         16108 => x"f0",
         16109 => x"1e",
         16110 => x"1f",
         16111 => x"f0",
         16112 => x"f0",
         16113 => x"f0",
         16114 => x"f0",
         16115 => x"81",
         16116 => x"f0",
         16117 => x"f0",
         16118 => x"b5",
         16119 => x"77",
         16120 => x"f0",
         16121 => x"70",
         16122 => x"a6",
         16123 => x"5d",
         16124 => x"33",
         16125 => x"6e",
         16126 => x"43",
         16127 => x"36",
         16128 => x"1e",
         16129 => x"9f",
         16130 => x"a3",
         16131 => x"c5",
         16132 => x"c4",
         16133 => x"f0",
         16134 => x"f0",
         16135 => x"81",
         16136 => x"f0",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"01",
         16163 => x"00",
         16164 => x"00",
         16165 => x"00",
         16166 => x"00",
         16167 => x"00",
         16168 => x"00",
         16169 => x"00",
         16170 => x"00",
         16171 => x"00",
         16172 => x"00",
         16173 => x"00",
         16174 => x"00",
         16175 => x"00",
         16176 => x"00",
         16177 => x"00",
         16178 => x"00",
         16179 => x"00",
         16180 => x"00",
         16181 => x"00",
         16182 => x"00",
         16183 => x"00",
         16184 => x"00",
         16185 => x"00",
         16186 => x"00",
         16187 => x"00",
         16188 => x"00",
         16189 => x"00",
         16190 => x"00",
         16191 => x"00",
         16192 => x"00",
         16193 => x"00",
         16194 => x"00",
         16195 => x"00",
         16196 => x"00",
         16197 => x"00",
         16198 => x"00",
         16199 => x"00",
         16200 => x"00",
         16201 => x"00",
         16202 => x"00",
         16203 => x"00",
         16204 => x"00",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"00",
         18207 => x"00",
         18208 => x"e0",
         18209 => x"cf",
         18210 => x"f9",
         18211 => x"fd",
         18212 => x"c1",
         18213 => x"c5",
         18214 => x"e4",
         18215 => x"ee",
         18216 => x"61",
         18217 => x"65",
         18218 => x"69",
         18219 => x"2a",
         18220 => x"21",
         18221 => x"25",
         18222 => x"29",
         18223 => x"2b",
         18224 => x"01",
         18225 => x"05",
         18226 => x"09",
         18227 => x"0d",
         18228 => x"11",
         18229 => x"15",
         18230 => x"19",
         18231 => x"54",
         18232 => x"81",
         18233 => x"85",
         18234 => x"89",
         18235 => x"8d",
         18236 => x"91",
         18237 => x"95",
         18238 => x"99",
         18239 => x"40",
         18240 => x"00",
         18241 => x"00",
         18242 => x"00",
         18243 => x"00",
         18244 => x"00",
         18245 => x"00",
         18246 => x"00",
         18247 => x"00",
         18248 => x"00",
         18249 => x"00",
         18250 => x"00",
         18251 => x"00",
         18252 => x"00",
         18253 => x"00",
         18254 => x"00",
         18255 => x"00",
         18256 => x"00",
         18257 => x"00",
         18258 => x"00",
         18259 => x"00",
         18260 => x"00",
         18261 => x"00",
         18262 => x"00",
         18263 => x"00",
         18264 => x"00",
         18265 => x"00",
         18266 => x"00",
         18267 => x"00",
         18268 => x"00",
         18269 => x"00",
         18270 => x"02",
         18271 => x"04",
         18272 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"cd",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"84",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cc",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"ab",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"96",
           269 => x"0b",
           270 => x"0b",
           271 => x"b6",
           272 => x"0b",
           273 => x"0b",
           274 => x"d6",
           275 => x"0b",
           276 => x"0b",
           277 => x"f6",
           278 => x"0b",
           279 => x"0b",
           280 => x"96",
           281 => x"0b",
           282 => x"0b",
           283 => x"b6",
           284 => x"0b",
           285 => x"0b",
           286 => x"d7",
           287 => x"0b",
           288 => x"0b",
           289 => x"f9",
           290 => x"0b",
           291 => x"0b",
           292 => x"9b",
           293 => x"0b",
           294 => x"0b",
           295 => x"bd",
           296 => x"0b",
           297 => x"0b",
           298 => x"df",
           299 => x"0b",
           300 => x"0b",
           301 => x"81",
           302 => x"0b",
           303 => x"0b",
           304 => x"a3",
           305 => x"0b",
           306 => x"0b",
           307 => x"c5",
           308 => x"0b",
           309 => x"0b",
           310 => x"e7",
           311 => x"0b",
           312 => x"0b",
           313 => x"89",
           314 => x"0b",
           315 => x"0b",
           316 => x"ab",
           317 => x"0b",
           318 => x"0b",
           319 => x"cd",
           320 => x"0b",
           321 => x"0b",
           322 => x"ef",
           323 => x"0b",
           324 => x"0b",
           325 => x"91",
           326 => x"0b",
           327 => x"0b",
           328 => x"b3",
           329 => x"0b",
           330 => x"0b",
           331 => x"d5",
           332 => x"0b",
           333 => x"0b",
           334 => x"f7",
           335 => x"0b",
           336 => x"0b",
           337 => x"99",
           338 => x"0b",
           339 => x"0b",
           340 => x"bb",
           341 => x"0b",
           342 => x"0b",
           343 => x"dc",
           344 => x"0b",
           345 => x"0b",
           346 => x"fe",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"90",
           390 => x"90",
           391 => x"2d",
           392 => x"08",
           393 => x"90",
           394 => x"90",
           395 => x"2d",
           396 => x"08",
           397 => x"90",
           398 => x"90",
           399 => x"2d",
           400 => x"08",
           401 => x"90",
           402 => x"90",
           403 => x"2d",
           404 => x"08",
           405 => x"90",
           406 => x"90",
           407 => x"2d",
           408 => x"08",
           409 => x"90",
           410 => x"90",
           411 => x"2d",
           412 => x"08",
           413 => x"90",
           414 => x"90",
           415 => x"2d",
           416 => x"08",
           417 => x"90",
           418 => x"90",
           419 => x"2d",
           420 => x"08",
           421 => x"90",
           422 => x"90",
           423 => x"2d",
           424 => x"08",
           425 => x"90",
           426 => x"90",
           427 => x"2d",
           428 => x"08",
           429 => x"90",
           430 => x"90",
           431 => x"2d",
           432 => x"08",
           433 => x"90",
           434 => x"90",
           435 => x"fc",
           436 => x"90",
           437 => x"80",
           438 => x"bb",
           439 => x"d5",
           440 => x"bb",
           441 => x"c0",
           442 => x"84",
           443 => x"80",
           444 => x"84",
           445 => x"80",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"90",
           451 => x"90",
           452 => x"f6",
           453 => x"90",
           454 => x"80",
           455 => x"bb",
           456 => x"e3",
           457 => x"bb",
           458 => x"c0",
           459 => x"84",
           460 => x"82",
           461 => x"84",
           462 => x"80",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"90",
           468 => x"90",
           469 => x"a6",
           470 => x"90",
           471 => x"80",
           472 => x"bb",
           473 => x"fa",
           474 => x"bb",
           475 => x"c0",
           476 => x"84",
           477 => x"82",
           478 => x"84",
           479 => x"80",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"90",
           485 => x"90",
           486 => x"e2",
           487 => x"90",
           488 => x"80",
           489 => x"bb",
           490 => x"f4",
           491 => x"bb",
           492 => x"c0",
           493 => x"84",
           494 => x"83",
           495 => x"84",
           496 => x"80",
           497 => x"04",
           498 => x"0c",
           499 => x"2d",
           500 => x"08",
           501 => x"90",
           502 => x"90",
           503 => x"95",
           504 => x"90",
           505 => x"80",
           506 => x"bb",
           507 => x"f6",
           508 => x"bb",
           509 => x"c0",
           510 => x"84",
           511 => x"83",
           512 => x"84",
           513 => x"80",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"90",
           519 => x"90",
           520 => x"d9",
           521 => x"90",
           522 => x"80",
           523 => x"bb",
           524 => x"e3",
           525 => x"bb",
           526 => x"c0",
           527 => x"84",
           528 => x"82",
           529 => x"84",
           530 => x"80",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"90",
           536 => x"90",
           537 => x"a9",
           538 => x"90",
           539 => x"80",
           540 => x"bb",
           541 => x"9b",
           542 => x"bb",
           543 => x"c0",
           544 => x"84",
           545 => x"83",
           546 => x"84",
           547 => x"80",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"90",
           553 => x"90",
           554 => x"a1",
           555 => x"90",
           556 => x"80",
           557 => x"bb",
           558 => x"ba",
           559 => x"bb",
           560 => x"c0",
           561 => x"84",
           562 => x"83",
           563 => x"84",
           564 => x"80",
           565 => x"04",
           566 => x"0c",
           567 => x"2d",
           568 => x"08",
           569 => x"90",
           570 => x"90",
           571 => x"aa",
           572 => x"90",
           573 => x"80",
           574 => x"bb",
           575 => x"f7",
           576 => x"bb",
           577 => x"c0",
           578 => x"84",
           579 => x"80",
           580 => x"84",
           581 => x"80",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"90",
           587 => x"90",
           588 => x"b5",
           589 => x"90",
           590 => x"80",
           591 => x"bb",
           592 => x"9a",
           593 => x"90",
           594 => x"80",
           595 => x"bb",
           596 => x"dc",
           597 => x"bb",
           598 => x"c0",
           599 => x"84",
           600 => x"81",
           601 => x"84",
           602 => x"80",
           603 => x"04",
           604 => x"0c",
           605 => x"2d",
           606 => x"08",
           607 => x"90",
           608 => x"90",
           609 => x"d9",
           610 => x"90",
           611 => x"80",
           612 => x"04",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"53",
           621 => x"00",
           622 => x"06",
           623 => x"09",
           624 => x"05",
           625 => x"2b",
           626 => x"06",
           627 => x"04",
           628 => x"72",
           629 => x"05",
           630 => x"05",
           631 => x"72",
           632 => x"53",
           633 => x"51",
           634 => x"04",
           635 => x"70",
           636 => x"27",
           637 => x"71",
           638 => x"53",
           639 => x"0b",
           640 => x"8c",
           641 => x"ce",
           642 => x"fc",
           643 => x"3d",
           644 => x"05",
           645 => x"53",
           646 => x"e6",
           647 => x"81",
           648 => x"3d",
           649 => x"3d",
           650 => x"7c",
           651 => x"81",
           652 => x"80",
           653 => x"56",
           654 => x"80",
           655 => x"2e",
           656 => x"80",
           657 => x"14",
           658 => x"32",
           659 => x"72",
           660 => x"51",
           661 => x"54",
           662 => x"b7",
           663 => x"2e",
           664 => x"51",
           665 => x"84",
           666 => x"53",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"05",
           671 => x"14",
           672 => x"70",
           673 => x"07",
           674 => x"54",
           675 => x"80",
           676 => x"80",
           677 => x"52",
           678 => x"84",
           679 => x"0d",
           680 => x"84",
           681 => x"88",
           682 => x"f5",
           683 => x"54",
           684 => x"05",
           685 => x"73",
           686 => x"58",
           687 => x"05",
           688 => x"8d",
           689 => x"51",
           690 => x"19",
           691 => x"34",
           692 => x"04",
           693 => x"86",
           694 => x"53",
           695 => x"51",
           696 => x"3d",
           697 => x"3d",
           698 => x"65",
           699 => x"80",
           700 => x"0c",
           701 => x"70",
           702 => x"32",
           703 => x"55",
           704 => x"72",
           705 => x"81",
           706 => x"38",
           707 => x"76",
           708 => x"c5",
           709 => x"7b",
           710 => x"5c",
           711 => x"81",
           712 => x"17",
           713 => x"26",
           714 => x"76",
           715 => x"30",
           716 => x"51",
           717 => x"ae",
           718 => x"2e",
           719 => x"83",
           720 => x"32",
           721 => x"54",
           722 => x"9e",
           723 => x"80",
           724 => x"33",
           725 => x"bd",
           726 => x"08",
           727 => x"bb",
           728 => x"3d",
           729 => x"83",
           730 => x"10",
           731 => x"10",
           732 => x"2b",
           733 => x"19",
           734 => x"0a",
           735 => x"05",
           736 => x"52",
           737 => x"5f",
           738 => x"81",
           739 => x"81",
           740 => x"ff",
           741 => x"7c",
           742 => x"76",
           743 => x"ff",
           744 => x"a5",
           745 => x"06",
           746 => x"73",
           747 => x"5b",
           748 => x"58",
           749 => x"dd",
           750 => x"39",
           751 => x"51",
           752 => x"7b",
           753 => x"fe",
           754 => x"8d",
           755 => x"2a",
           756 => x"54",
           757 => x"38",
           758 => x"06",
           759 => x"95",
           760 => x"53",
           761 => x"26",
           762 => x"10",
           763 => x"94",
           764 => x"08",
           765 => x"18",
           766 => x"d8",
           767 => x"38",
           768 => x"51",
           769 => x"80",
           770 => x"5b",
           771 => x"38",
           772 => x"80",
           773 => x"f6",
           774 => x"7f",
           775 => x"71",
           776 => x"ff",
           777 => x"58",
           778 => x"bb",
           779 => x"52",
           780 => x"9a",
           781 => x"84",
           782 => x"06",
           783 => x"08",
           784 => x"56",
           785 => x"26",
           786 => x"bb",
           787 => x"05",
           788 => x"70",
           789 => x"34",
           790 => x"51",
           791 => x"84",
           792 => x"56",
           793 => x"08",
           794 => x"84",
           795 => x"98",
           796 => x"06",
           797 => x"80",
           798 => x"77",
           799 => x"29",
           800 => x"05",
           801 => x"59",
           802 => x"2a",
           803 => x"55",
           804 => x"2e",
           805 => x"84",
           806 => x"f8",
           807 => x"53",
           808 => x"8b",
           809 => x"80",
           810 => x"80",
           811 => x"72",
           812 => x"7a",
           813 => x"81",
           814 => x"72",
           815 => x"38",
           816 => x"70",
           817 => x"54",
           818 => x"24",
           819 => x"7a",
           820 => x"06",
           821 => x"71",
           822 => x"56",
           823 => x"06",
           824 => x"2e",
           825 => x"77",
           826 => x"2b",
           827 => x"7c",
           828 => x"56",
           829 => x"80",
           830 => x"38",
           831 => x"81",
           832 => x"85",
           833 => x"84",
           834 => x"54",
           835 => x"38",
           836 => x"81",
           837 => x"86",
           838 => x"81",
           839 => x"85",
           840 => x"88",
           841 => x"5f",
           842 => x"b2",
           843 => x"84",
           844 => x"fc",
           845 => x"70",
           846 => x"40",
           847 => x"25",
           848 => x"52",
           849 => x"a9",
           850 => x"84",
           851 => x"fc",
           852 => x"70",
           853 => x"40",
           854 => x"24",
           855 => x"81",
           856 => x"80",
           857 => x"78",
           858 => x"0a",
           859 => x"0a",
           860 => x"2c",
           861 => x"80",
           862 => x"38",
           863 => x"51",
           864 => x"78",
           865 => x"0a",
           866 => x"0a",
           867 => x"2c",
           868 => x"74",
           869 => x"38",
           870 => x"70",
           871 => x"55",
           872 => x"81",
           873 => x"80",
           874 => x"d8",
           875 => x"f3",
           876 => x"38",
           877 => x"2e",
           878 => x"7d",
           879 => x"2e",
           880 => x"52",
           881 => x"33",
           882 => x"a5",
           883 => x"bb",
           884 => x"81",
           885 => x"74",
           886 => x"7a",
           887 => x"a7",
           888 => x"84",
           889 => x"fc",
           890 => x"70",
           891 => x"40",
           892 => x"25",
           893 => x"7c",
           894 => x"86",
           895 => x"39",
           896 => x"5b",
           897 => x"7c",
           898 => x"76",
           899 => x"fa",
           900 => x"80",
           901 => x"80",
           902 => x"60",
           903 => x"71",
           904 => x"ff",
           905 => x"59",
           906 => x"fb",
           907 => x"60",
           908 => x"fe",
           909 => x"83",
           910 => x"98",
           911 => x"7c",
           912 => x"29",
           913 => x"05",
           914 => x"5e",
           915 => x"57",
           916 => x"87",
           917 => x"06",
           918 => x"fe",
           919 => x"78",
           920 => x"29",
           921 => x"05",
           922 => x"5a",
           923 => x"7f",
           924 => x"38",
           925 => x"51",
           926 => x"e2",
           927 => x"70",
           928 => x"06",
           929 => x"83",
           930 => x"fe",
           931 => x"52",
           932 => x"05",
           933 => x"85",
           934 => x"39",
           935 => x"83",
           936 => x"5b",
           937 => x"ff",
           938 => x"ab",
           939 => x"75",
           940 => x"57",
           941 => x"b9",
           942 => x"75",
           943 => x"81",
           944 => x"78",
           945 => x"29",
           946 => x"05",
           947 => x"5a",
           948 => x"e3",
           949 => x"70",
           950 => x"56",
           951 => x"c6",
           952 => x"39",
           953 => x"05",
           954 => x"53",
           955 => x"80",
           956 => x"df",
           957 => x"ff",
           958 => x"84",
           959 => x"fa",
           960 => x"84",
           961 => x"58",
           962 => x"89",
           963 => x"39",
           964 => x"5b",
           965 => x"58",
           966 => x"f9",
           967 => x"39",
           968 => x"05",
           969 => x"81",
           970 => x"41",
           971 => x"8a",
           972 => x"87",
           973 => x"bb",
           974 => x"ff",
           975 => x"71",
           976 => x"54",
           977 => x"2c",
           978 => x"39",
           979 => x"07",
           980 => x"5b",
           981 => x"38",
           982 => x"7f",
           983 => x"71",
           984 => x"06",
           985 => x"54",
           986 => x"38",
           987 => x"bb",
           988 => x"84",
           989 => x"ff",
           990 => x"31",
           991 => x"5a",
           992 => x"81",
           993 => x"33",
           994 => x"f7",
           995 => x"c9",
           996 => x"84",
           997 => x"fc",
           998 => x"70",
           999 => x"54",
          1000 => x"25",
          1001 => x"7c",
          1002 => x"83",
          1003 => x"39",
          1004 => x"51",
          1005 => x"79",
          1006 => x"81",
          1007 => x"38",
          1008 => x"51",
          1009 => x"7a",
          1010 => x"06",
          1011 => x"2e",
          1012 => x"fa",
          1013 => x"98",
          1014 => x"31",
          1015 => x"90",
          1016 => x"80",
          1017 => x"51",
          1018 => x"90",
          1019 => x"39",
          1020 => x"51",
          1021 => x"7e",
          1022 => x"73",
          1023 => x"a2",
          1024 => x"39",
          1025 => x"98",
          1026 => x"e5",
          1027 => x"06",
          1028 => x"2e",
          1029 => x"fb",
          1030 => x"74",
          1031 => x"70",
          1032 => x"53",
          1033 => x"7c",
          1034 => x"82",
          1035 => x"39",
          1036 => x"51",
          1037 => x"ff",
          1038 => x"52",
          1039 => x"8b",
          1040 => x"84",
          1041 => x"ff",
          1042 => x"31",
          1043 => x"5a",
          1044 => x"7a",
          1045 => x"30",
          1046 => x"bf",
          1047 => x"5b",
          1048 => x"fe",
          1049 => x"e6",
          1050 => x"75",
          1051 => x"f3",
          1052 => x"3d",
          1053 => x"3d",
          1054 => x"80",
          1055 => x"e8",
          1056 => x"33",
          1057 => x"81",
          1058 => x"06",
          1059 => x"55",
          1060 => x"72",
          1061 => x"81",
          1062 => x"38",
          1063 => x"05",
          1064 => x"72",
          1065 => x"38",
          1066 => x"08",
          1067 => x"90",
          1068 => x"72",
          1069 => x"84",
          1070 => x"83",
          1071 => x"74",
          1072 => x"56",
          1073 => x"80",
          1074 => x"84",
          1075 => x"54",
          1076 => x"e6",
          1077 => x"84",
          1078 => x"52",
          1079 => x"14",
          1080 => x"2d",
          1081 => x"08",
          1082 => x"38",
          1083 => x"56",
          1084 => x"84",
          1085 => x"0d",
          1086 => x"0d",
          1087 => x"54",
          1088 => x"16",
          1089 => x"2a",
          1090 => x"81",
          1091 => x"57",
          1092 => x"72",
          1093 => x"81",
          1094 => x"73",
          1095 => x"55",
          1096 => x"77",
          1097 => x"06",
          1098 => x"56",
          1099 => x"84",
          1100 => x"0d",
          1101 => x"81",
          1102 => x"53",
          1103 => x"ea",
          1104 => x"72",
          1105 => x"08",
          1106 => x"84",
          1107 => x"80",
          1108 => x"ff",
          1109 => x"05",
          1110 => x"57",
          1111 => x"ca",
          1112 => x"0d",
          1113 => x"08",
          1114 => x"85",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"11",
          1118 => x"2a",
          1119 => x"06",
          1120 => x"57",
          1121 => x"ae",
          1122 => x"2a",
          1123 => x"73",
          1124 => x"38",
          1125 => x"53",
          1126 => x"08",
          1127 => x"74",
          1128 => x"76",
          1129 => x"81",
          1130 => x"8c",
          1131 => x"81",
          1132 => x"0c",
          1133 => x"84",
          1134 => x"88",
          1135 => x"74",
          1136 => x"ff",
          1137 => x"15",
          1138 => x"2d",
          1139 => x"bb",
          1140 => x"38",
          1141 => x"81",
          1142 => x"0c",
          1143 => x"39",
          1144 => x"77",
          1145 => x"70",
          1146 => x"70",
          1147 => x"06",
          1148 => x"56",
          1149 => x"b3",
          1150 => x"2a",
          1151 => x"71",
          1152 => x"82",
          1153 => x"52",
          1154 => x"80",
          1155 => x"08",
          1156 => x"53",
          1157 => x"80",
          1158 => x"13",
          1159 => x"16",
          1160 => x"8c",
          1161 => x"81",
          1162 => x"73",
          1163 => x"0c",
          1164 => x"04",
          1165 => x"06",
          1166 => x"17",
          1167 => x"08",
          1168 => x"17",
          1169 => x"33",
          1170 => x"0c",
          1171 => x"04",
          1172 => x"16",
          1173 => x"2d",
          1174 => x"08",
          1175 => x"84",
          1176 => x"ff",
          1177 => x"16",
          1178 => x"07",
          1179 => x"bb",
          1180 => x"2e",
          1181 => x"a0",
          1182 => x"85",
          1183 => x"54",
          1184 => x"84",
          1185 => x"0d",
          1186 => x"07",
          1187 => x"17",
          1188 => x"ec",
          1189 => x"0d",
          1190 => x"54",
          1191 => x"70",
          1192 => x"33",
          1193 => x"38",
          1194 => x"72",
          1195 => x"54",
          1196 => x"72",
          1197 => x"54",
          1198 => x"38",
          1199 => x"84",
          1200 => x"0d",
          1201 => x"0d",
          1202 => x"7a",
          1203 => x"54",
          1204 => x"9d",
          1205 => x"27",
          1206 => x"80",
          1207 => x"71",
          1208 => x"53",
          1209 => x"81",
          1210 => x"ff",
          1211 => x"ef",
          1212 => x"bb",
          1213 => x"3d",
          1214 => x"12",
          1215 => x"27",
          1216 => x"14",
          1217 => x"ff",
          1218 => x"53",
          1219 => x"73",
          1220 => x"51",
          1221 => x"d9",
          1222 => x"ff",
          1223 => x"71",
          1224 => x"ff",
          1225 => x"df",
          1226 => x"fe",
          1227 => x"70",
          1228 => x"70",
          1229 => x"33",
          1230 => x"38",
          1231 => x"74",
          1232 => x"84",
          1233 => x"3d",
          1234 => x"3d",
          1235 => x"71",
          1236 => x"72",
          1237 => x"54",
          1238 => x"72",
          1239 => x"54",
          1240 => x"38",
          1241 => x"84",
          1242 => x"0d",
          1243 => x"0d",
          1244 => x"79",
          1245 => x"54",
          1246 => x"93",
          1247 => x"81",
          1248 => x"73",
          1249 => x"55",
          1250 => x"51",
          1251 => x"73",
          1252 => x"0c",
          1253 => x"04",
          1254 => x"76",
          1255 => x"56",
          1256 => x"2e",
          1257 => x"33",
          1258 => x"05",
          1259 => x"52",
          1260 => x"09",
          1261 => x"38",
          1262 => x"71",
          1263 => x"38",
          1264 => x"72",
          1265 => x"51",
          1266 => x"84",
          1267 => x"0d",
          1268 => x"2e",
          1269 => x"33",
          1270 => x"72",
          1271 => x"38",
          1272 => x"52",
          1273 => x"80",
          1274 => x"72",
          1275 => x"bb",
          1276 => x"3d",
          1277 => x"84",
          1278 => x"86",
          1279 => x"fb",
          1280 => x"79",
          1281 => x"56",
          1282 => x"84",
          1283 => x"84",
          1284 => x"81",
          1285 => x"81",
          1286 => x"84",
          1287 => x"54",
          1288 => x"08",
          1289 => x"38",
          1290 => x"08",
          1291 => x"74",
          1292 => x"75",
          1293 => x"84",
          1294 => x"b1",
          1295 => x"84",
          1296 => x"84",
          1297 => x"87",
          1298 => x"fd",
          1299 => x"77",
          1300 => x"55",
          1301 => x"80",
          1302 => x"72",
          1303 => x"54",
          1304 => x"80",
          1305 => x"ff",
          1306 => x"ff",
          1307 => x"06",
          1308 => x"13",
          1309 => x"52",
          1310 => x"bb",
          1311 => x"3d",
          1312 => x"3d",
          1313 => x"79",
          1314 => x"54",
          1315 => x"2e",
          1316 => x"72",
          1317 => x"54",
          1318 => x"51",
          1319 => x"73",
          1320 => x"0c",
          1321 => x"04",
          1322 => x"78",
          1323 => x"a0",
          1324 => x"2e",
          1325 => x"51",
          1326 => x"84",
          1327 => x"52",
          1328 => x"73",
          1329 => x"38",
          1330 => x"e3",
          1331 => x"bb",
          1332 => x"53",
          1333 => x"9f",
          1334 => x"38",
          1335 => x"9f",
          1336 => x"38",
          1337 => x"71",
          1338 => x"31",
          1339 => x"57",
          1340 => x"80",
          1341 => x"2e",
          1342 => x"10",
          1343 => x"07",
          1344 => x"07",
          1345 => x"ff",
          1346 => x"70",
          1347 => x"72",
          1348 => x"31",
          1349 => x"56",
          1350 => x"58",
          1351 => x"da",
          1352 => x"76",
          1353 => x"84",
          1354 => x"88",
          1355 => x"fc",
          1356 => x"70",
          1357 => x"06",
          1358 => x"72",
          1359 => x"70",
          1360 => x"71",
          1361 => x"2a",
          1362 => x"80",
          1363 => x"70",
          1364 => x"2b",
          1365 => x"74",
          1366 => x"81",
          1367 => x"30",
          1368 => x"82",
          1369 => x"31",
          1370 => x"55",
          1371 => x"05",
          1372 => x"70",
          1373 => x"25",
          1374 => x"31",
          1375 => x"70",
          1376 => x"32",
          1377 => x"70",
          1378 => x"31",
          1379 => x"05",
          1380 => x"0c",
          1381 => x"55",
          1382 => x"5a",
          1383 => x"55",
          1384 => x"56",
          1385 => x"56",
          1386 => x"3d",
          1387 => x"3d",
          1388 => x"70",
          1389 => x"54",
          1390 => x"3f",
          1391 => x"08",
          1392 => x"71",
          1393 => x"84",
          1394 => x"3d",
          1395 => x"3d",
          1396 => x"58",
          1397 => x"76",
          1398 => x"38",
          1399 => x"cf",
          1400 => x"84",
          1401 => x"13",
          1402 => x"2e",
          1403 => x"51",
          1404 => x"72",
          1405 => x"08",
          1406 => x"53",
          1407 => x"80",
          1408 => x"53",
          1409 => x"be",
          1410 => x"74",
          1411 => x"72",
          1412 => x"2b",
          1413 => x"55",
          1414 => x"76",
          1415 => x"72",
          1416 => x"2a",
          1417 => x"77",
          1418 => x"31",
          1419 => x"2c",
          1420 => x"7b",
          1421 => x"71",
          1422 => x"5c",
          1423 => x"55",
          1424 => x"74",
          1425 => x"84",
          1426 => x"88",
          1427 => x"fa",
          1428 => x"9f",
          1429 => x"2c",
          1430 => x"7b",
          1431 => x"2c",
          1432 => x"73",
          1433 => x"31",
          1434 => x"31",
          1435 => x"59",
          1436 => x"b4",
          1437 => x"84",
          1438 => x"75",
          1439 => x"84",
          1440 => x"0d",
          1441 => x"0d",
          1442 => x"57",
          1443 => x"0c",
          1444 => x"33",
          1445 => x"73",
          1446 => x"81",
          1447 => x"81",
          1448 => x"0c",
          1449 => x"55",
          1450 => x"f3",
          1451 => x"2e",
          1452 => x"73",
          1453 => x"83",
          1454 => x"58",
          1455 => x"89",
          1456 => x"38",
          1457 => x"56",
          1458 => x"80",
          1459 => x"e0",
          1460 => x"38",
          1461 => x"81",
          1462 => x"53",
          1463 => x"81",
          1464 => x"53",
          1465 => x"8f",
          1466 => x"70",
          1467 => x"54",
          1468 => x"27",
          1469 => x"72",
          1470 => x"83",
          1471 => x"29",
          1472 => x"70",
          1473 => x"33",
          1474 => x"73",
          1475 => x"be",
          1476 => x"2e",
          1477 => x"30",
          1478 => x"0c",
          1479 => x"84",
          1480 => x"8b",
          1481 => x"81",
          1482 => x"79",
          1483 => x"56",
          1484 => x"b0",
          1485 => x"06",
          1486 => x"81",
          1487 => x"0c",
          1488 => x"55",
          1489 => x"2e",
          1490 => x"58",
          1491 => x"2e",
          1492 => x"56",
          1493 => x"c6",
          1494 => x"53",
          1495 => x"58",
          1496 => x"fe",
          1497 => x"84",
          1498 => x"8b",
          1499 => x"82",
          1500 => x"70",
          1501 => x"33",
          1502 => x"56",
          1503 => x"80",
          1504 => x"84",
          1505 => x"0d",
          1506 => x"0d",
          1507 => x"57",
          1508 => x"0c",
          1509 => x"33",
          1510 => x"73",
          1511 => x"81",
          1512 => x"81",
          1513 => x"0c",
          1514 => x"55",
          1515 => x"f3",
          1516 => x"2e",
          1517 => x"73",
          1518 => x"83",
          1519 => x"58",
          1520 => x"89",
          1521 => x"38",
          1522 => x"56",
          1523 => x"80",
          1524 => x"e0",
          1525 => x"38",
          1526 => x"81",
          1527 => x"53",
          1528 => x"81",
          1529 => x"53",
          1530 => x"8f",
          1531 => x"70",
          1532 => x"54",
          1533 => x"27",
          1534 => x"72",
          1535 => x"83",
          1536 => x"29",
          1537 => x"70",
          1538 => x"33",
          1539 => x"73",
          1540 => x"be",
          1541 => x"2e",
          1542 => x"30",
          1543 => x"0c",
          1544 => x"84",
          1545 => x"8b",
          1546 => x"81",
          1547 => x"79",
          1548 => x"56",
          1549 => x"b0",
          1550 => x"06",
          1551 => x"81",
          1552 => x"0c",
          1553 => x"55",
          1554 => x"2e",
          1555 => x"58",
          1556 => x"2e",
          1557 => x"56",
          1558 => x"c6",
          1559 => x"53",
          1560 => x"58",
          1561 => x"fe",
          1562 => x"84",
          1563 => x"8b",
          1564 => x"82",
          1565 => x"70",
          1566 => x"33",
          1567 => x"56",
          1568 => x"80",
          1569 => x"84",
          1570 => x"0d",
          1571 => x"aa",
          1572 => x"84",
          1573 => x"06",
          1574 => x"0c",
          1575 => x"0d",
          1576 => x"93",
          1577 => x"71",
          1578 => x"bf",
          1579 => x"71",
          1580 => x"cf",
          1581 => x"be",
          1582 => x"0d",
          1583 => x"bc",
          1584 => x"3f",
          1585 => x"04",
          1586 => x"51",
          1587 => x"83",
          1588 => x"83",
          1589 => x"ef",
          1590 => x"3d",
          1591 => x"d0",
          1592 => x"92",
          1593 => x"0d",
          1594 => x"94",
          1595 => x"3f",
          1596 => x"04",
          1597 => x"51",
          1598 => x"83",
          1599 => x"83",
          1600 => x"ee",
          1601 => x"3d",
          1602 => x"d0",
          1603 => x"e6",
          1604 => x"0d",
          1605 => x"80",
          1606 => x"3f",
          1607 => x"04",
          1608 => x"51",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ee",
          1612 => x"3d",
          1613 => x"d1",
          1614 => x"ba",
          1615 => x"0d",
          1616 => x"e4",
          1617 => x"3f",
          1618 => x"04",
          1619 => x"51",
          1620 => x"83",
          1621 => x"83",
          1622 => x"ee",
          1623 => x"3d",
          1624 => x"d2",
          1625 => x"8e",
          1626 => x"0d",
          1627 => x"a8",
          1628 => x"3f",
          1629 => x"04",
          1630 => x"51",
          1631 => x"83",
          1632 => x"83",
          1633 => x"ed",
          1634 => x"3d",
          1635 => x"d2",
          1636 => x"e2",
          1637 => x"0d",
          1638 => x"3d",
          1639 => x"3d",
          1640 => x"05",
          1641 => x"33",
          1642 => x"0b",
          1643 => x"08",
          1644 => x"7b",
          1645 => x"51",
          1646 => x"78",
          1647 => x"ff",
          1648 => x"81",
          1649 => x"07",
          1650 => x"06",
          1651 => x"57",
          1652 => x"38",
          1653 => x"52",
          1654 => x"52",
          1655 => x"99",
          1656 => x"84",
          1657 => x"bb",
          1658 => x"2e",
          1659 => x"77",
          1660 => x"98",
          1661 => x"70",
          1662 => x"25",
          1663 => x"9f",
          1664 => x"53",
          1665 => x"77",
          1666 => x"38",
          1667 => x"88",
          1668 => x"87",
          1669 => x"e3",
          1670 => x"78",
          1671 => x"51",
          1672 => x"84",
          1673 => x"54",
          1674 => x"53",
          1675 => x"d2",
          1676 => x"d7",
          1677 => x"bb",
          1678 => x"96",
          1679 => x"84",
          1680 => x"87",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"3d",
          1684 => x"54",
          1685 => x"75",
          1686 => x"82",
          1687 => x"84",
          1688 => x"57",
          1689 => x"08",
          1690 => x"7a",
          1691 => x"2e",
          1692 => x"74",
          1693 => x"57",
          1694 => x"87",
          1695 => x"51",
          1696 => x"84",
          1697 => x"52",
          1698 => x"9c",
          1699 => x"84",
          1700 => x"d3",
          1701 => x"52",
          1702 => x"51",
          1703 => x"ff",
          1704 => x"3d",
          1705 => x"84",
          1706 => x"33",
          1707 => x"58",
          1708 => x"52",
          1709 => x"e1",
          1710 => x"84",
          1711 => x"76",
          1712 => x"38",
          1713 => x"8a",
          1714 => x"bb",
          1715 => x"3d",
          1716 => x"04",
          1717 => x"56",
          1718 => x"54",
          1719 => x"53",
          1720 => x"51",
          1721 => x"bb",
          1722 => x"bb",
          1723 => x"3d",
          1724 => x"3d",
          1725 => x"63",
          1726 => x"80",
          1727 => x"73",
          1728 => x"41",
          1729 => x"5f",
          1730 => x"80",
          1731 => x"38",
          1732 => x"d3",
          1733 => x"f3",
          1734 => x"94",
          1735 => x"3f",
          1736 => x"79",
          1737 => x"7c",
          1738 => x"ed",
          1739 => x"2e",
          1740 => x"73",
          1741 => x"7a",
          1742 => x"38",
          1743 => x"83",
          1744 => x"dd",
          1745 => x"14",
          1746 => x"08",
          1747 => x"51",
          1748 => x"78",
          1749 => x"38",
          1750 => x"51",
          1751 => x"80",
          1752 => x"27",
          1753 => x"75",
          1754 => x"55",
          1755 => x"72",
          1756 => x"38",
          1757 => x"53",
          1758 => x"83",
          1759 => x"74",
          1760 => x"81",
          1761 => x"57",
          1762 => x"88",
          1763 => x"74",
          1764 => x"38",
          1765 => x"08",
          1766 => x"eb",
          1767 => x"16",
          1768 => x"26",
          1769 => x"d3",
          1770 => x"ca",
          1771 => x"79",
          1772 => x"80",
          1773 => x"3f",
          1774 => x"08",
          1775 => x"98",
          1776 => x"76",
          1777 => x"ee",
          1778 => x"2e",
          1779 => x"7b",
          1780 => x"78",
          1781 => x"38",
          1782 => x"bb",
          1783 => x"3d",
          1784 => x"d3",
          1785 => x"a3",
          1786 => x"84",
          1787 => x"53",
          1788 => x"ea",
          1789 => x"74",
          1790 => x"38",
          1791 => x"83",
          1792 => x"dc",
          1793 => x"14",
          1794 => x"08",
          1795 => x"51",
          1796 => x"73",
          1797 => x"c0",
          1798 => x"53",
          1799 => x"df",
          1800 => x"52",
          1801 => x"51",
          1802 => x"82",
          1803 => x"e8",
          1804 => x"a0",
          1805 => x"3f",
          1806 => x"dd",
          1807 => x"39",
          1808 => x"51",
          1809 => x"84",
          1810 => x"e8",
          1811 => x"a0",
          1812 => x"3f",
          1813 => x"fd",
          1814 => x"18",
          1815 => x"27",
          1816 => x"08",
          1817 => x"8c",
          1818 => x"3f",
          1819 => x"e6",
          1820 => x"54",
          1821 => x"f9",
          1822 => x"26",
          1823 => x"d8",
          1824 => x"e8",
          1825 => x"51",
          1826 => x"81",
          1827 => x"91",
          1828 => x"a6",
          1829 => x"84",
          1830 => x"06",
          1831 => x"72",
          1832 => x"ec",
          1833 => x"72",
          1834 => x"09",
          1835 => x"e0",
          1836 => x"fc",
          1837 => x"51",
          1838 => x"84",
          1839 => x"98",
          1840 => x"2c",
          1841 => x"70",
          1842 => x"32",
          1843 => x"72",
          1844 => x"07",
          1845 => x"58",
          1846 => x"53",
          1847 => x"fd",
          1848 => x"51",
          1849 => x"84",
          1850 => x"98",
          1851 => x"2c",
          1852 => x"70",
          1853 => x"32",
          1854 => x"72",
          1855 => x"07",
          1856 => x"58",
          1857 => x"53",
          1858 => x"ff",
          1859 => x"b9",
          1860 => x"84",
          1861 => x"8f",
          1862 => x"fe",
          1863 => x"c0",
          1864 => x"53",
          1865 => x"81",
          1866 => x"3f",
          1867 => x"51",
          1868 => x"80",
          1869 => x"3f",
          1870 => x"70",
          1871 => x"52",
          1872 => x"38",
          1873 => x"70",
          1874 => x"52",
          1875 => x"38",
          1876 => x"70",
          1877 => x"52",
          1878 => x"38",
          1879 => x"70",
          1880 => x"52",
          1881 => x"38",
          1882 => x"70",
          1883 => x"52",
          1884 => x"38",
          1885 => x"70",
          1886 => x"52",
          1887 => x"38",
          1888 => x"70",
          1889 => x"52",
          1890 => x"72",
          1891 => x"06",
          1892 => x"38",
          1893 => x"84",
          1894 => x"81",
          1895 => x"3f",
          1896 => x"51",
          1897 => x"80",
          1898 => x"3f",
          1899 => x"84",
          1900 => x"81",
          1901 => x"3f",
          1902 => x"51",
          1903 => x"80",
          1904 => x"3f",
          1905 => x"81",
          1906 => x"80",
          1907 => x"cb",
          1908 => x"9b",
          1909 => x"d5",
          1910 => x"f4",
          1911 => x"9b",
          1912 => x"87",
          1913 => x"06",
          1914 => x"80",
          1915 => x"38",
          1916 => x"51",
          1917 => x"83",
          1918 => x"9b",
          1919 => x"51",
          1920 => x"72",
          1921 => x"81",
          1922 => x"71",
          1923 => x"f0",
          1924 => x"39",
          1925 => x"a0",
          1926 => x"b8",
          1927 => x"3f",
          1928 => x"94",
          1929 => x"2a",
          1930 => x"51",
          1931 => x"2e",
          1932 => x"ff",
          1933 => x"51",
          1934 => x"83",
          1935 => x"9b",
          1936 => x"51",
          1937 => x"72",
          1938 => x"81",
          1939 => x"71",
          1940 => x"94",
          1941 => x"39",
          1942 => x"dc",
          1943 => x"e0",
          1944 => x"3f",
          1945 => x"d0",
          1946 => x"2a",
          1947 => x"51",
          1948 => x"2e",
          1949 => x"ff",
          1950 => x"51",
          1951 => x"83",
          1952 => x"9a",
          1953 => x"51",
          1954 => x"72",
          1955 => x"81",
          1956 => x"71",
          1957 => x"b8",
          1958 => x"39",
          1959 => x"80",
          1960 => x"ff",
          1961 => x"90",
          1962 => x"52",
          1963 => x"b7",
          1964 => x"bb",
          1965 => x"ff",
          1966 => x"40",
          1967 => x"2e",
          1968 => x"83",
          1969 => x"e3",
          1970 => x"3d",
          1971 => x"fc",
          1972 => x"3f",
          1973 => x"f8",
          1974 => x"7e",
          1975 => x"3f",
          1976 => x"ef",
          1977 => x"81",
          1978 => x"59",
          1979 => x"82",
          1980 => x"81",
          1981 => x"38",
          1982 => x"06",
          1983 => x"2e",
          1984 => x"67",
          1985 => x"79",
          1986 => x"e0",
          1987 => x"5c",
          1988 => x"09",
          1989 => x"38",
          1990 => x"33",
          1991 => x"a0",
          1992 => x"80",
          1993 => x"26",
          1994 => x"90",
          1995 => x"fc",
          1996 => x"52",
          1997 => x"3f",
          1998 => x"08",
          1999 => x"08",
          2000 => x"7b",
          2001 => x"e8",
          2002 => x"bb",
          2003 => x"38",
          2004 => x"5e",
          2005 => x"83",
          2006 => x"1c",
          2007 => x"06",
          2008 => x"7c",
          2009 => x"9a",
          2010 => x"7b",
          2011 => x"dd",
          2012 => x"52",
          2013 => x"87",
          2014 => x"84",
          2015 => x"bb",
          2016 => x"2e",
          2017 => x"84",
          2018 => x"48",
          2019 => x"80",
          2020 => x"a9",
          2021 => x"84",
          2022 => x"06",
          2023 => x"80",
          2024 => x"38",
          2025 => x"08",
          2026 => x"3f",
          2027 => x"08",
          2028 => x"f3",
          2029 => x"a5",
          2030 => x"7a",
          2031 => x"8a",
          2032 => x"24",
          2033 => x"7a",
          2034 => x"e8",
          2035 => x"80",
          2036 => x"80",
          2037 => x"d5",
          2038 => x"f3",
          2039 => x"bb",
          2040 => x"56",
          2041 => x"54",
          2042 => x"53",
          2043 => x"52",
          2044 => x"ae",
          2045 => x"84",
          2046 => x"84",
          2047 => x"30",
          2048 => x"80",
          2049 => x"5b",
          2050 => x"7a",
          2051 => x"38",
          2052 => x"7a",
          2053 => x"80",
          2054 => x"81",
          2055 => x"ff",
          2056 => x"7a",
          2057 => x"7f",
          2058 => x"81",
          2059 => x"7c",
          2060 => x"61",
          2061 => x"ec",
          2062 => x"81",
          2063 => x"83",
          2064 => x"d3",
          2065 => x"48",
          2066 => x"80",
          2067 => x"e8",
          2068 => x"0b",
          2069 => x"33",
          2070 => x"06",
          2071 => x"fd",
          2072 => x"53",
          2073 => x"52",
          2074 => x"51",
          2075 => x"3f",
          2076 => x"08",
          2077 => x"81",
          2078 => x"83",
          2079 => x"84",
          2080 => x"80",
          2081 => x"51",
          2082 => x"3f",
          2083 => x"08",
          2084 => x"38",
          2085 => x"08",
          2086 => x"3f",
          2087 => x"ef",
          2088 => x"81",
          2089 => x"59",
          2090 => x"09",
          2091 => x"d3",
          2092 => x"84",
          2093 => x"82",
          2094 => x"82",
          2095 => x"83",
          2096 => x"80",
          2097 => x"b8",
          2098 => x"80",
          2099 => x"51",
          2100 => x"67",
          2101 => x"79",
          2102 => x"90",
          2103 => x"63",
          2104 => x"33",
          2105 => x"89",
          2106 => x"38",
          2107 => x"83",
          2108 => x"5a",
          2109 => x"83",
          2110 => x"88",
          2111 => x"e4",
          2112 => x"53",
          2113 => x"c8",
          2114 => x"86",
          2115 => x"bb",
          2116 => x"2e",
          2117 => x"fb",
          2118 => x"70",
          2119 => x"41",
          2120 => x"39",
          2121 => x"51",
          2122 => x"7d",
          2123 => x"ac",
          2124 => x"39",
          2125 => x"56",
          2126 => x"d7",
          2127 => x"53",
          2128 => x"52",
          2129 => x"e3",
          2130 => x"39",
          2131 => x"3f",
          2132 => x"9a",
          2133 => x"f5",
          2134 => x"83",
          2135 => x"dc",
          2136 => x"39",
          2137 => x"3f",
          2138 => x"83",
          2139 => x"de",
          2140 => x"59",
          2141 => x"d7",
          2142 => x"fa",
          2143 => x"3f",
          2144 => x"b8",
          2145 => x"11",
          2146 => x"05",
          2147 => x"3f",
          2148 => x"08",
          2149 => x"b5",
          2150 => x"83",
          2151 => x"d0",
          2152 => x"5a",
          2153 => x"bb",
          2154 => x"2e",
          2155 => x"84",
          2156 => x"52",
          2157 => x"51",
          2158 => x"fa",
          2159 => x"3d",
          2160 => x"53",
          2161 => x"51",
          2162 => x"84",
          2163 => x"80",
          2164 => x"38",
          2165 => x"d8",
          2166 => x"af",
          2167 => x"78",
          2168 => x"fe",
          2169 => x"ff",
          2170 => x"e9",
          2171 => x"bb",
          2172 => x"2e",
          2173 => x"b8",
          2174 => x"11",
          2175 => x"05",
          2176 => x"3f",
          2177 => x"08",
          2178 => x"64",
          2179 => x"53",
          2180 => x"d8",
          2181 => x"f3",
          2182 => x"e4",
          2183 => x"f8",
          2184 => x"d0",
          2185 => x"48",
          2186 => x"78",
          2187 => x"9d",
          2188 => x"26",
          2189 => x"64",
          2190 => x"46",
          2191 => x"b8",
          2192 => x"11",
          2193 => x"05",
          2194 => x"3f",
          2195 => x"08",
          2196 => x"f9",
          2197 => x"fe",
          2198 => x"ff",
          2199 => x"e8",
          2200 => x"bb",
          2201 => x"b0",
          2202 => x"78",
          2203 => x"52",
          2204 => x"51",
          2205 => x"84",
          2206 => x"53",
          2207 => x"7e",
          2208 => x"3f",
          2209 => x"33",
          2210 => x"2e",
          2211 => x"78",
          2212 => x"ca",
          2213 => x"05",
          2214 => x"cf",
          2215 => x"ff",
          2216 => x"ff",
          2217 => x"e9",
          2218 => x"bb",
          2219 => x"2e",
          2220 => x"b8",
          2221 => x"11",
          2222 => x"05",
          2223 => x"3f",
          2224 => x"08",
          2225 => x"85",
          2226 => x"fe",
          2227 => x"ff",
          2228 => x"e9",
          2229 => x"bb",
          2230 => x"2e",
          2231 => x"83",
          2232 => x"ce",
          2233 => x"67",
          2234 => x"7c",
          2235 => x"38",
          2236 => x"7a",
          2237 => x"5a",
          2238 => x"95",
          2239 => x"79",
          2240 => x"53",
          2241 => x"d8",
          2242 => x"ff",
          2243 => x"5b",
          2244 => x"81",
          2245 => x"d2",
          2246 => x"ff",
          2247 => x"ff",
          2248 => x"e8",
          2249 => x"bb",
          2250 => x"2e",
          2251 => x"b8",
          2252 => x"11",
          2253 => x"05",
          2254 => x"3f",
          2255 => x"08",
          2256 => x"89",
          2257 => x"fe",
          2258 => x"ff",
          2259 => x"e8",
          2260 => x"bb",
          2261 => x"2e",
          2262 => x"83",
          2263 => x"cd",
          2264 => x"5a",
          2265 => x"82",
          2266 => x"5c",
          2267 => x"05",
          2268 => x"34",
          2269 => x"46",
          2270 => x"3d",
          2271 => x"53",
          2272 => x"51",
          2273 => x"84",
          2274 => x"80",
          2275 => x"38",
          2276 => x"fc",
          2277 => x"80",
          2278 => x"ed",
          2279 => x"84",
          2280 => x"68",
          2281 => x"52",
          2282 => x"51",
          2283 => x"84",
          2284 => x"53",
          2285 => x"7e",
          2286 => x"3f",
          2287 => x"33",
          2288 => x"2e",
          2289 => x"78",
          2290 => x"97",
          2291 => x"05",
          2292 => x"68",
          2293 => x"db",
          2294 => x"34",
          2295 => x"49",
          2296 => x"fc",
          2297 => x"80",
          2298 => x"9d",
          2299 => x"84",
          2300 => x"f5",
          2301 => x"59",
          2302 => x"05",
          2303 => x"68",
          2304 => x"b8",
          2305 => x"11",
          2306 => x"05",
          2307 => x"3f",
          2308 => x"08",
          2309 => x"f5",
          2310 => x"3d",
          2311 => x"53",
          2312 => x"51",
          2313 => x"84",
          2314 => x"80",
          2315 => x"38",
          2316 => x"fc",
          2317 => x"80",
          2318 => x"cd",
          2319 => x"84",
          2320 => x"f5",
          2321 => x"3d",
          2322 => x"53",
          2323 => x"51",
          2324 => x"84",
          2325 => x"86",
          2326 => x"84",
          2327 => x"d9",
          2328 => x"a7",
          2329 => x"5b",
          2330 => x"27",
          2331 => x"5b",
          2332 => x"84",
          2333 => x"79",
          2334 => x"38",
          2335 => x"e1",
          2336 => x"39",
          2337 => x"80",
          2338 => x"b1",
          2339 => x"84",
          2340 => x"ff",
          2341 => x"59",
          2342 => x"81",
          2343 => x"84",
          2344 => x"51",
          2345 => x"84",
          2346 => x"80",
          2347 => x"38",
          2348 => x"08",
          2349 => x"3f",
          2350 => x"b8",
          2351 => x"11",
          2352 => x"05",
          2353 => x"3f",
          2354 => x"08",
          2355 => x"f4",
          2356 => x"79",
          2357 => x"c0",
          2358 => x"c0",
          2359 => x"3d",
          2360 => x"53",
          2361 => x"51",
          2362 => x"84",
          2363 => x"91",
          2364 => x"88",
          2365 => x"80",
          2366 => x"38",
          2367 => x"08",
          2368 => x"fe",
          2369 => x"ff",
          2370 => x"e4",
          2371 => x"bb",
          2372 => x"2e",
          2373 => x"66",
          2374 => x"88",
          2375 => x"81",
          2376 => x"32",
          2377 => x"72",
          2378 => x"7e",
          2379 => x"5d",
          2380 => x"88",
          2381 => x"2e",
          2382 => x"46",
          2383 => x"51",
          2384 => x"80",
          2385 => x"65",
          2386 => x"68",
          2387 => x"3f",
          2388 => x"51",
          2389 => x"f2",
          2390 => x"64",
          2391 => x"64",
          2392 => x"b8",
          2393 => x"11",
          2394 => x"05",
          2395 => x"3f",
          2396 => x"08",
          2397 => x"d5",
          2398 => x"71",
          2399 => x"84",
          2400 => x"3d",
          2401 => x"53",
          2402 => x"51",
          2403 => x"84",
          2404 => x"c6",
          2405 => x"39",
          2406 => x"80",
          2407 => x"7e",
          2408 => x"40",
          2409 => x"b8",
          2410 => x"11",
          2411 => x"05",
          2412 => x"3f",
          2413 => x"08",
          2414 => x"91",
          2415 => x"02",
          2416 => x"22",
          2417 => x"05",
          2418 => x"45",
          2419 => x"f0",
          2420 => x"80",
          2421 => x"ad",
          2422 => x"84",
          2423 => x"38",
          2424 => x"b8",
          2425 => x"11",
          2426 => x"05",
          2427 => x"3f",
          2428 => x"08",
          2429 => x"dc",
          2430 => x"02",
          2431 => x"33",
          2432 => x"81",
          2433 => x"9b",
          2434 => x"fe",
          2435 => x"ff",
          2436 => x"e0",
          2437 => x"bb",
          2438 => x"2e",
          2439 => x"64",
          2440 => x"5d",
          2441 => x"70",
          2442 => x"e1",
          2443 => x"2e",
          2444 => x"f3",
          2445 => x"55",
          2446 => x"54",
          2447 => x"d9",
          2448 => x"51",
          2449 => x"f3",
          2450 => x"52",
          2451 => x"fa",
          2452 => x"39",
          2453 => x"51",
          2454 => x"f0",
          2455 => x"3d",
          2456 => x"53",
          2457 => x"51",
          2458 => x"84",
          2459 => x"80",
          2460 => x"64",
          2461 => x"ce",
          2462 => x"70",
          2463 => x"23",
          2464 => x"e7",
          2465 => x"89",
          2466 => x"80",
          2467 => x"38",
          2468 => x"08",
          2469 => x"39",
          2470 => x"33",
          2471 => x"2e",
          2472 => x"f3",
          2473 => x"fc",
          2474 => x"d9",
          2475 => x"c6",
          2476 => x"f7",
          2477 => x"d9",
          2478 => x"ba",
          2479 => x"f6",
          2480 => x"f4",
          2481 => x"78",
          2482 => x"38",
          2483 => x"08",
          2484 => x"39",
          2485 => x"51",
          2486 => x"f9",
          2487 => x"f4",
          2488 => x"78",
          2489 => x"38",
          2490 => x"08",
          2491 => x"39",
          2492 => x"33",
          2493 => x"2e",
          2494 => x"f3",
          2495 => x"fb",
          2496 => x"f4",
          2497 => x"7d",
          2498 => x"38",
          2499 => x"08",
          2500 => x"39",
          2501 => x"33",
          2502 => x"2e",
          2503 => x"f3",
          2504 => x"fb",
          2505 => x"f4",
          2506 => x"7c",
          2507 => x"38",
          2508 => x"08",
          2509 => x"39",
          2510 => x"08",
          2511 => x"49",
          2512 => x"83",
          2513 => x"88",
          2514 => x"b5",
          2515 => x"0d",
          2516 => x"bb",
          2517 => x"c0",
          2518 => x"08",
          2519 => x"84",
          2520 => x"51",
          2521 => x"84",
          2522 => x"90",
          2523 => x"57",
          2524 => x"80",
          2525 => x"da",
          2526 => x"84",
          2527 => x"07",
          2528 => x"c0",
          2529 => x"08",
          2530 => x"84",
          2531 => x"51",
          2532 => x"84",
          2533 => x"90",
          2534 => x"57",
          2535 => x"80",
          2536 => x"da",
          2537 => x"84",
          2538 => x"07",
          2539 => x"80",
          2540 => x"c0",
          2541 => x"8c",
          2542 => x"87",
          2543 => x"0c",
          2544 => x"5c",
          2545 => x"5d",
          2546 => x"05",
          2547 => x"80",
          2548 => x"e4",
          2549 => x"70",
          2550 => x"70",
          2551 => x"e6",
          2552 => x"b8",
          2553 => x"9e",
          2554 => x"3f",
          2555 => x"95",
          2556 => x"d3",
          2557 => x"d3",
          2558 => x"8f",
          2559 => x"f4",
          2560 => x"55",
          2561 => x"83",
          2562 => x"83",
          2563 => x"81",
          2564 => x"83",
          2565 => x"c3",
          2566 => x"b2",
          2567 => x"fc",
          2568 => x"3f",
          2569 => x"d4",
          2570 => x"df",
          2571 => x"0a",
          2572 => x"a8",
          2573 => x"3f",
          2574 => x"80",
          2575 => x"0d",
          2576 => x"56",
          2577 => x"52",
          2578 => x"2e",
          2579 => x"74",
          2580 => x"ff",
          2581 => x"70",
          2582 => x"81",
          2583 => x"81",
          2584 => x"70",
          2585 => x"53",
          2586 => x"a0",
          2587 => x"71",
          2588 => x"54",
          2589 => x"81",
          2590 => x"52",
          2591 => x"80",
          2592 => x"72",
          2593 => x"ff",
          2594 => x"54",
          2595 => x"83",
          2596 => x"70",
          2597 => x"38",
          2598 => x"86",
          2599 => x"52",
          2600 => x"73",
          2601 => x"52",
          2602 => x"2e",
          2603 => x"83",
          2604 => x"70",
          2605 => x"30",
          2606 => x"76",
          2607 => x"53",
          2608 => x"88",
          2609 => x"70",
          2610 => x"34",
          2611 => x"74",
          2612 => x"bb",
          2613 => x"3d",
          2614 => x"80",
          2615 => x"73",
          2616 => x"be",
          2617 => x"52",
          2618 => x"70",
          2619 => x"53",
          2620 => x"a2",
          2621 => x"81",
          2622 => x"81",
          2623 => x"75",
          2624 => x"81",
          2625 => x"06",
          2626 => x"dc",
          2627 => x"0d",
          2628 => x"08",
          2629 => x"0b",
          2630 => x"0c",
          2631 => x"04",
          2632 => x"05",
          2633 => x"da",
          2634 => x"bb",
          2635 => x"2e",
          2636 => x"84",
          2637 => x"86",
          2638 => x"fc",
          2639 => x"82",
          2640 => x"05",
          2641 => x"52",
          2642 => x"81",
          2643 => x"13",
          2644 => x"54",
          2645 => x"9e",
          2646 => x"38",
          2647 => x"51",
          2648 => x"97",
          2649 => x"38",
          2650 => x"54",
          2651 => x"bb",
          2652 => x"38",
          2653 => x"55",
          2654 => x"bb",
          2655 => x"38",
          2656 => x"55",
          2657 => x"87",
          2658 => x"d9",
          2659 => x"22",
          2660 => x"73",
          2661 => x"80",
          2662 => x"0b",
          2663 => x"9c",
          2664 => x"87",
          2665 => x"0c",
          2666 => x"87",
          2667 => x"0c",
          2668 => x"87",
          2669 => x"0c",
          2670 => x"87",
          2671 => x"0c",
          2672 => x"87",
          2673 => x"0c",
          2674 => x"87",
          2675 => x"0c",
          2676 => x"98",
          2677 => x"87",
          2678 => x"0c",
          2679 => x"c0",
          2680 => x"80",
          2681 => x"bb",
          2682 => x"3d",
          2683 => x"3d",
          2684 => x"87",
          2685 => x"5d",
          2686 => x"87",
          2687 => x"08",
          2688 => x"23",
          2689 => x"b8",
          2690 => x"82",
          2691 => x"c0",
          2692 => x"5a",
          2693 => x"34",
          2694 => x"b0",
          2695 => x"84",
          2696 => x"c0",
          2697 => x"5a",
          2698 => x"34",
          2699 => x"a8",
          2700 => x"86",
          2701 => x"c0",
          2702 => x"5c",
          2703 => x"23",
          2704 => x"a0",
          2705 => x"8a",
          2706 => x"7d",
          2707 => x"ff",
          2708 => x"7b",
          2709 => x"06",
          2710 => x"33",
          2711 => x"33",
          2712 => x"33",
          2713 => x"33",
          2714 => x"33",
          2715 => x"ff",
          2716 => x"83",
          2717 => x"ff",
          2718 => x"8f",
          2719 => x"fe",
          2720 => x"93",
          2721 => x"72",
          2722 => x"38",
          2723 => x"e9",
          2724 => x"bb",
          2725 => x"2b",
          2726 => x"51",
          2727 => x"2e",
          2728 => x"86",
          2729 => x"2e",
          2730 => x"84",
          2731 => x"84",
          2732 => x"72",
          2733 => x"b7",
          2734 => x"84",
          2735 => x"70",
          2736 => x"52",
          2737 => x"09",
          2738 => x"38",
          2739 => x"e9",
          2740 => x"bb",
          2741 => x"2b",
          2742 => x"51",
          2743 => x"2e",
          2744 => x"39",
          2745 => x"80",
          2746 => x"71",
          2747 => x"81",
          2748 => x"fb",
          2749 => x"84",
          2750 => x"70",
          2751 => x"52",
          2752 => x"eb",
          2753 => x"07",
          2754 => x"52",
          2755 => x"db",
          2756 => x"bb",
          2757 => x"3d",
          2758 => x"3d",
          2759 => x"05",
          2760 => x"bc",
          2761 => x"ff",
          2762 => x"55",
          2763 => x"80",
          2764 => x"c0",
          2765 => x"70",
          2766 => x"81",
          2767 => x"52",
          2768 => x"8c",
          2769 => x"2a",
          2770 => x"51",
          2771 => x"38",
          2772 => x"81",
          2773 => x"80",
          2774 => x"71",
          2775 => x"06",
          2776 => x"38",
          2777 => x"06",
          2778 => x"94",
          2779 => x"80",
          2780 => x"87",
          2781 => x"52",
          2782 => x"74",
          2783 => x"0c",
          2784 => x"04",
          2785 => x"70",
          2786 => x"51",
          2787 => x"72",
          2788 => x"06",
          2789 => x"2e",
          2790 => x"93",
          2791 => x"52",
          2792 => x"c0",
          2793 => x"94",
          2794 => x"96",
          2795 => x"06",
          2796 => x"70",
          2797 => x"39",
          2798 => x"02",
          2799 => x"70",
          2800 => x"2a",
          2801 => x"70",
          2802 => x"34",
          2803 => x"04",
          2804 => x"78",
          2805 => x"33",
          2806 => x"57",
          2807 => x"80",
          2808 => x"15",
          2809 => x"33",
          2810 => x"06",
          2811 => x"71",
          2812 => x"ff",
          2813 => x"94",
          2814 => x"96",
          2815 => x"06",
          2816 => x"70",
          2817 => x"38",
          2818 => x"70",
          2819 => x"51",
          2820 => x"72",
          2821 => x"06",
          2822 => x"2e",
          2823 => x"93",
          2824 => x"52",
          2825 => x"75",
          2826 => x"51",
          2827 => x"80",
          2828 => x"2e",
          2829 => x"c0",
          2830 => x"73",
          2831 => x"17",
          2832 => x"57",
          2833 => x"38",
          2834 => x"84",
          2835 => x"0d",
          2836 => x"2a",
          2837 => x"51",
          2838 => x"38",
          2839 => x"81",
          2840 => x"80",
          2841 => x"71",
          2842 => x"06",
          2843 => x"2e",
          2844 => x"87",
          2845 => x"08",
          2846 => x"70",
          2847 => x"54",
          2848 => x"38",
          2849 => x"3d",
          2850 => x"9e",
          2851 => x"9c",
          2852 => x"52",
          2853 => x"2e",
          2854 => x"87",
          2855 => x"08",
          2856 => x"0c",
          2857 => x"a8",
          2858 => x"c4",
          2859 => x"9e",
          2860 => x"f3",
          2861 => x"c0",
          2862 => x"83",
          2863 => x"87",
          2864 => x"08",
          2865 => x"0c",
          2866 => x"a0",
          2867 => x"d4",
          2868 => x"9e",
          2869 => x"f3",
          2870 => x"c0",
          2871 => x"83",
          2872 => x"87",
          2873 => x"08",
          2874 => x"0c",
          2875 => x"b8",
          2876 => x"e4",
          2877 => x"9e",
          2878 => x"f3",
          2879 => x"c0",
          2880 => x"83",
          2881 => x"87",
          2882 => x"08",
          2883 => x"0c",
          2884 => x"80",
          2885 => x"83",
          2886 => x"87",
          2887 => x"08",
          2888 => x"0c",
          2889 => x"88",
          2890 => x"fc",
          2891 => x"9e",
          2892 => x"f4",
          2893 => x"0b",
          2894 => x"34",
          2895 => x"c0",
          2896 => x"70",
          2897 => x"06",
          2898 => x"70",
          2899 => x"71",
          2900 => x"34",
          2901 => x"c0",
          2902 => x"70",
          2903 => x"06",
          2904 => x"70",
          2905 => x"38",
          2906 => x"83",
          2907 => x"80",
          2908 => x"9e",
          2909 => x"90",
          2910 => x"51",
          2911 => x"80",
          2912 => x"81",
          2913 => x"f4",
          2914 => x"0b",
          2915 => x"90",
          2916 => x"80",
          2917 => x"52",
          2918 => x"2e",
          2919 => x"52",
          2920 => x"88",
          2921 => x"87",
          2922 => x"08",
          2923 => x"80",
          2924 => x"52",
          2925 => x"83",
          2926 => x"71",
          2927 => x"34",
          2928 => x"c0",
          2929 => x"70",
          2930 => x"06",
          2931 => x"70",
          2932 => x"38",
          2933 => x"83",
          2934 => x"80",
          2935 => x"9e",
          2936 => x"84",
          2937 => x"51",
          2938 => x"80",
          2939 => x"81",
          2940 => x"f4",
          2941 => x"0b",
          2942 => x"90",
          2943 => x"80",
          2944 => x"52",
          2945 => x"2e",
          2946 => x"52",
          2947 => x"8c",
          2948 => x"87",
          2949 => x"08",
          2950 => x"80",
          2951 => x"52",
          2952 => x"83",
          2953 => x"71",
          2954 => x"34",
          2955 => x"c0",
          2956 => x"70",
          2957 => x"06",
          2958 => x"70",
          2959 => x"38",
          2960 => x"83",
          2961 => x"80",
          2962 => x"9e",
          2963 => x"a0",
          2964 => x"52",
          2965 => x"2e",
          2966 => x"52",
          2967 => x"8f",
          2968 => x"9e",
          2969 => x"80",
          2970 => x"2a",
          2971 => x"83",
          2972 => x"80",
          2973 => x"9e",
          2974 => x"84",
          2975 => x"52",
          2976 => x"2e",
          2977 => x"52",
          2978 => x"91",
          2979 => x"9e",
          2980 => x"f0",
          2981 => x"2a",
          2982 => x"83",
          2983 => x"80",
          2984 => x"9e",
          2985 => x"88",
          2986 => x"52",
          2987 => x"83",
          2988 => x"71",
          2989 => x"34",
          2990 => x"90",
          2991 => x"51",
          2992 => x"94",
          2993 => x"0d",
          2994 => x"fd",
          2995 => x"3d",
          2996 => x"94",
          2997 => x"b3",
          2998 => x"84",
          2999 => x"86",
          3000 => x"da",
          3001 => x"8e",
          3002 => x"86",
          3003 => x"85",
          3004 => x"f4",
          3005 => x"73",
          3006 => x"83",
          3007 => x"56",
          3008 => x"38",
          3009 => x"33",
          3010 => x"f5",
          3011 => x"8a",
          3012 => x"84",
          3013 => x"f4",
          3014 => x"75",
          3015 => x"83",
          3016 => x"54",
          3017 => x"38",
          3018 => x"33",
          3019 => x"e3",
          3020 => x"85",
          3021 => x"83",
          3022 => x"f4",
          3023 => x"73",
          3024 => x"83",
          3025 => x"55",
          3026 => x"38",
          3027 => x"33",
          3028 => x"ea",
          3029 => x"8e",
          3030 => x"81",
          3031 => x"da",
          3032 => x"92",
          3033 => x"e8",
          3034 => x"da",
          3035 => x"b5",
          3036 => x"f3",
          3037 => x"83",
          3038 => x"ff",
          3039 => x"83",
          3040 => x"52",
          3041 => x"51",
          3042 => x"3f",
          3043 => x"51",
          3044 => x"83",
          3045 => x"52",
          3046 => x"51",
          3047 => x"3f",
          3048 => x"08",
          3049 => x"c0",
          3050 => x"c9",
          3051 => x"bb",
          3052 => x"84",
          3053 => x"71",
          3054 => x"84",
          3055 => x"52",
          3056 => x"51",
          3057 => x"3f",
          3058 => x"33",
          3059 => x"38",
          3060 => x"33",
          3061 => x"38",
          3062 => x"04",
          3063 => x"08",
          3064 => x"c0",
          3065 => x"c9",
          3066 => x"bb",
          3067 => x"84",
          3068 => x"71",
          3069 => x"84",
          3070 => x"52",
          3071 => x"51",
          3072 => x"3f",
          3073 => x"04",
          3074 => x"08",
          3075 => x"c0",
          3076 => x"c9",
          3077 => x"bb",
          3078 => x"84",
          3079 => x"71",
          3080 => x"84",
          3081 => x"52",
          3082 => x"51",
          3083 => x"3f",
          3084 => x"33",
          3085 => x"2e",
          3086 => x"ff",
          3087 => x"dc",
          3088 => x"b2",
          3089 => x"c0",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"cc",
          3093 => x"b3",
          3094 => x"ec",
          3095 => x"da",
          3096 => x"b3",
          3097 => x"f3",
          3098 => x"83",
          3099 => x"ff",
          3100 => x"83",
          3101 => x"ff",
          3102 => x"83",
          3103 => x"52",
          3104 => x"51",
          3105 => x"3f",
          3106 => x"08",
          3107 => x"c0",
          3108 => x"c8",
          3109 => x"bb",
          3110 => x"84",
          3111 => x"71",
          3112 => x"84",
          3113 => x"52",
          3114 => x"51",
          3115 => x"3f",
          3116 => x"33",
          3117 => x"2e",
          3118 => x"fe",
          3119 => x"dd",
          3120 => x"bf",
          3121 => x"f4",
          3122 => x"73",
          3123 => x"8e",
          3124 => x"39",
          3125 => x"51",
          3126 => x"3f",
          3127 => x"33",
          3128 => x"2e",
          3129 => x"d6",
          3130 => x"94",
          3131 => x"86",
          3132 => x"8c",
          3133 => x"80",
          3134 => x"38",
          3135 => x"dd",
          3136 => x"be",
          3137 => x"f4",
          3138 => x"73",
          3139 => x"b3",
          3140 => x"83",
          3141 => x"52",
          3142 => x"51",
          3143 => x"3f",
          3144 => x"33",
          3145 => x"2e",
          3146 => x"d2",
          3147 => x"94",
          3148 => x"dd",
          3149 => x"b1",
          3150 => x"f4",
          3151 => x"74",
          3152 => x"ed",
          3153 => x"83",
          3154 => x"52",
          3155 => x"51",
          3156 => x"3f",
          3157 => x"33",
          3158 => x"2e",
          3159 => x"cd",
          3160 => x"d0",
          3161 => x"d4",
          3162 => x"52",
          3163 => x"51",
          3164 => x"3f",
          3165 => x"33",
          3166 => x"2e",
          3167 => x"c7",
          3168 => x"c8",
          3169 => x"cc",
          3170 => x"52",
          3171 => x"51",
          3172 => x"3f",
          3173 => x"33",
          3174 => x"2e",
          3175 => x"c1",
          3176 => x"c0",
          3177 => x"c4",
          3178 => x"52",
          3179 => x"51",
          3180 => x"3f",
          3181 => x"33",
          3182 => x"2e",
          3183 => x"c1",
          3184 => x"d8",
          3185 => x"dc",
          3186 => x"52",
          3187 => x"51",
          3188 => x"3f",
          3189 => x"33",
          3190 => x"2e",
          3191 => x"c1",
          3192 => x"e0",
          3193 => x"e4",
          3194 => x"52",
          3195 => x"51",
          3196 => x"3f",
          3197 => x"33",
          3198 => x"2e",
          3199 => x"c1",
          3200 => x"a0",
          3201 => x"83",
          3202 => x"a8",
          3203 => x"e6",
          3204 => x"86",
          3205 => x"80",
          3206 => x"38",
          3207 => x"3d",
          3208 => x"05",
          3209 => x"85",
          3210 => x"71",
          3211 => x"c4",
          3212 => x"71",
          3213 => x"df",
          3214 => x"af",
          3215 => x"3d",
          3216 => x"df",
          3217 => x"af",
          3218 => x"3d",
          3219 => x"df",
          3220 => x"af",
          3221 => x"3d",
          3222 => x"df",
          3223 => x"af",
          3224 => x"3d",
          3225 => x"df",
          3226 => x"af",
          3227 => x"3d",
          3228 => x"df",
          3229 => x"af",
          3230 => x"3d",
          3231 => x"88",
          3232 => x"80",
          3233 => x"96",
          3234 => x"83",
          3235 => x"87",
          3236 => x"0c",
          3237 => x"0d",
          3238 => x"ad",
          3239 => x"5a",
          3240 => x"58",
          3241 => x"f4",
          3242 => x"82",
          3243 => x"84",
          3244 => x"80",
          3245 => x"3d",
          3246 => x"83",
          3247 => x"54",
          3248 => x"52",
          3249 => x"d3",
          3250 => x"bb",
          3251 => x"2e",
          3252 => x"51",
          3253 => x"84",
          3254 => x"81",
          3255 => x"80",
          3256 => x"84",
          3257 => x"38",
          3258 => x"08",
          3259 => x"18",
          3260 => x"74",
          3261 => x"70",
          3262 => x"07",
          3263 => x"55",
          3264 => x"2e",
          3265 => x"ff",
          3266 => x"f4",
          3267 => x"11",
          3268 => x"82",
          3269 => x"84",
          3270 => x"8f",
          3271 => x"2e",
          3272 => x"84",
          3273 => x"a9",
          3274 => x"83",
          3275 => x"ff",
          3276 => x"78",
          3277 => x"81",
          3278 => x"76",
          3279 => x"c0",
          3280 => x"51",
          3281 => x"3f",
          3282 => x"56",
          3283 => x"08",
          3284 => x"52",
          3285 => x"51",
          3286 => x"3f",
          3287 => x"bb",
          3288 => x"3d",
          3289 => x"3d",
          3290 => x"08",
          3291 => x"71",
          3292 => x"33",
          3293 => x"57",
          3294 => x"81",
          3295 => x"0b",
          3296 => x"56",
          3297 => x"10",
          3298 => x"05",
          3299 => x"54",
          3300 => x"3f",
          3301 => x"08",
          3302 => x"73",
          3303 => x"bf",
          3304 => x"bb",
          3305 => x"38",
          3306 => x"54",
          3307 => x"81",
          3308 => x"82",
          3309 => x"81",
          3310 => x"ff",
          3311 => x"82",
          3312 => x"38",
          3313 => x"84",
          3314 => x"aa",
          3315 => x"81",
          3316 => x"3d",
          3317 => x"53",
          3318 => x"51",
          3319 => x"84",
          3320 => x"80",
          3321 => x"ff",
          3322 => x"52",
          3323 => x"a5",
          3324 => x"84",
          3325 => x"06",
          3326 => x"2e",
          3327 => x"16",
          3328 => x"06",
          3329 => x"76",
          3330 => x"38",
          3331 => x"78",
          3332 => x"56",
          3333 => x"fe",
          3334 => x"15",
          3335 => x"33",
          3336 => x"a0",
          3337 => x"06",
          3338 => x"75",
          3339 => x"38",
          3340 => x"3d",
          3341 => x"cc",
          3342 => x"bb",
          3343 => x"83",
          3344 => x"52",
          3345 => x"e1",
          3346 => x"84",
          3347 => x"38",
          3348 => x"08",
          3349 => x"52",
          3350 => x"cf",
          3351 => x"bb",
          3352 => x"2e",
          3353 => x"51",
          3354 => x"3f",
          3355 => x"08",
          3356 => x"84",
          3357 => x"25",
          3358 => x"bb",
          3359 => x"05",
          3360 => x"55",
          3361 => x"77",
          3362 => x"81",
          3363 => x"ac",
          3364 => x"aa",
          3365 => x"ff",
          3366 => x"06",
          3367 => x"81",
          3368 => x"84",
          3369 => x"0d",
          3370 => x"0d",
          3371 => x"b8",
          3372 => x"3d",
          3373 => x"08",
          3374 => x"42",
          3375 => x"5c",
          3376 => x"3d",
          3377 => x"f4",
          3378 => x"83",
          3379 => x"83",
          3380 => x"55",
          3381 => x"74",
          3382 => x"06",
          3383 => x"80",
          3384 => x"38",
          3385 => x"91",
          3386 => x"70",
          3387 => x"56",
          3388 => x"38",
          3389 => x"90",
          3390 => x"3d",
          3391 => x"40",
          3392 => x"fb",
          3393 => x"84",
          3394 => x"70",
          3395 => x"57",
          3396 => x"81",
          3397 => x"81",
          3398 => x"e2",
          3399 => x"98",
          3400 => x"2c",
          3401 => x"33",
          3402 => x"70",
          3403 => x"98",
          3404 => x"10",
          3405 => x"e0",
          3406 => x"15",
          3407 => x"53",
          3408 => x"52",
          3409 => x"59",
          3410 => x"79",
          3411 => x"38",
          3412 => x"81",
          3413 => x"81",
          3414 => x"81",
          3415 => x"70",
          3416 => x"42",
          3417 => x"81",
          3418 => x"10",
          3419 => x"2b",
          3420 => x"0b",
          3421 => x"16",
          3422 => x"77",
          3423 => x"38",
          3424 => x"15",
          3425 => x"33",
          3426 => x"75",
          3427 => x"38",
          3428 => x"c2",
          3429 => x"e2",
          3430 => x"57",
          3431 => x"81",
          3432 => x"1b",
          3433 => x"70",
          3434 => x"e2",
          3435 => x"98",
          3436 => x"2c",
          3437 => x"05",
          3438 => x"83",
          3439 => x"33",
          3440 => x"5e",
          3441 => x"57",
          3442 => x"81",
          3443 => x"84",
          3444 => x"80",
          3445 => x"3f",
          3446 => x"08",
          3447 => x"98",
          3448 => x"79",
          3449 => x"81",
          3450 => x"38",
          3451 => x"fe",
          3452 => x"2d",
          3453 => x"81",
          3454 => x"99",
          3455 => x"80",
          3456 => x"80",
          3457 => x"98",
          3458 => x"ff",
          3459 => x"42",
          3460 => x"80",
          3461 => x"10",
          3462 => x"2b",
          3463 => x"0b",
          3464 => x"16",
          3465 => x"77",
          3466 => x"38",
          3467 => x"15",
          3468 => x"33",
          3469 => x"62",
          3470 => x"38",
          3471 => x"ff",
          3472 => x"d1",
          3473 => x"76",
          3474 => x"8a",
          3475 => x"39",
          3476 => x"90",
          3477 => x"76",
          3478 => x"76",
          3479 => x"34",
          3480 => x"bc",
          3481 => x"34",
          3482 => x"63",
          3483 => x"26",
          3484 => x"74",
          3485 => x"c4",
          3486 => x"76",
          3487 => x"df",
          3488 => x"60",
          3489 => x"84",
          3490 => x"80",
          3491 => x"bc",
          3492 => x"84",
          3493 => x"56",
          3494 => x"fc",
          3495 => x"e6",
          3496 => x"88",
          3497 => x"c9",
          3498 => x"c8",
          3499 => x"5b",
          3500 => x"c8",
          3501 => x"39",
          3502 => x"33",
          3503 => x"06",
          3504 => x"33",
          3505 => x"75",
          3506 => x"b4",
          3507 => x"e8",
          3508 => x"15",
          3509 => x"e2",
          3510 => x"16",
          3511 => x"55",
          3512 => x"3f",
          3513 => x"7c",
          3514 => x"bd",
          3515 => x"26",
          3516 => x"10",
          3517 => x"a0",
          3518 => x"57",
          3519 => x"a5",
          3520 => x"84",
          3521 => x"80",
          3522 => x"e2",
          3523 => x"e2",
          3524 => x"56",
          3525 => x"b6",
          3526 => x"e8",
          3527 => x"51",
          3528 => x"3f",
          3529 => x"08",
          3530 => x"ff",
          3531 => x"84",
          3532 => x"52",
          3533 => x"b4",
          3534 => x"e2",
          3535 => x"05",
          3536 => x"e2",
          3537 => x"81",
          3538 => x"74",
          3539 => x"51",
          3540 => x"3f",
          3541 => x"c8",
          3542 => x"39",
          3543 => x"83",
          3544 => x"56",
          3545 => x"38",
          3546 => x"81",
          3547 => x"58",
          3548 => x"90",
          3549 => x"10",
          3550 => x"05",
          3551 => x"55",
          3552 => x"38",
          3553 => x"fa",
          3554 => x"10",
          3555 => x"9c",
          3556 => x"57",
          3557 => x"2e",
          3558 => x"75",
          3559 => x"8b",
          3560 => x"84",
          3561 => x"c4",
          3562 => x"84",
          3563 => x"06",
          3564 => x"75",
          3565 => x"ff",
          3566 => x"84",
          3567 => x"84",
          3568 => x"56",
          3569 => x"2e",
          3570 => x"84",
          3571 => x"52",
          3572 => x"b3",
          3573 => x"e6",
          3574 => x"a0",
          3575 => x"91",
          3576 => x"e8",
          3577 => x"51",
          3578 => x"3f",
          3579 => x"33",
          3580 => x"74",
          3581 => x"34",
          3582 => x"06",
          3583 => x"84",
          3584 => x"70",
          3585 => x"84",
          3586 => x"5c",
          3587 => x"7a",
          3588 => x"38",
          3589 => x"08",
          3590 => x"57",
          3591 => x"c8",
          3592 => x"70",
          3593 => x"ff",
          3594 => x"84",
          3595 => x"70",
          3596 => x"84",
          3597 => x"5a",
          3598 => x"78",
          3599 => x"38",
          3600 => x"08",
          3601 => x"57",
          3602 => x"c8",
          3603 => x"70",
          3604 => x"ff",
          3605 => x"84",
          3606 => x"70",
          3607 => x"84",
          3608 => x"5a",
          3609 => x"76",
          3610 => x"38",
          3611 => x"84",
          3612 => x"84",
          3613 => x"56",
          3614 => x"2e",
          3615 => x"ff",
          3616 => x"84",
          3617 => x"75",
          3618 => x"98",
          3619 => x"ff",
          3620 => x"59",
          3621 => x"80",
          3622 => x"e6",
          3623 => x"a0",
          3624 => x"cd",
          3625 => x"c8",
          3626 => x"2b",
          3627 => x"84",
          3628 => x"5a",
          3629 => x"74",
          3630 => x"c4",
          3631 => x"e8",
          3632 => x"51",
          3633 => x"3f",
          3634 => x"0a",
          3635 => x"0a",
          3636 => x"2c",
          3637 => x"33",
          3638 => x"74",
          3639 => x"a0",
          3640 => x"e8",
          3641 => x"51",
          3642 => x"3f",
          3643 => x"0a",
          3644 => x"0a",
          3645 => x"2c",
          3646 => x"33",
          3647 => x"7a",
          3648 => x"b9",
          3649 => x"39",
          3650 => x"81",
          3651 => x"34",
          3652 => x"08",
          3653 => x"51",
          3654 => x"3f",
          3655 => x"0a",
          3656 => x"0a",
          3657 => x"2c",
          3658 => x"33",
          3659 => x"75",
          3660 => x"e6",
          3661 => x"58",
          3662 => x"78",
          3663 => x"e8",
          3664 => x"33",
          3665 => x"a9",
          3666 => x"80",
          3667 => x"80",
          3668 => x"98",
          3669 => x"c4",
          3670 => x"55",
          3671 => x"ff",
          3672 => x"b6",
          3673 => x"c8",
          3674 => x"80",
          3675 => x"38",
          3676 => x"08",
          3677 => x"ff",
          3678 => x"84",
          3679 => x"ff",
          3680 => x"84",
          3681 => x"76",
          3682 => x"55",
          3683 => x"e2",
          3684 => x"05",
          3685 => x"34",
          3686 => x"08",
          3687 => x"ff",
          3688 => x"84",
          3689 => x"7b",
          3690 => x"3f",
          3691 => x"08",
          3692 => x"58",
          3693 => x"38",
          3694 => x"33",
          3695 => x"2e",
          3696 => x"83",
          3697 => x"70",
          3698 => x"f4",
          3699 => x"08",
          3700 => x"74",
          3701 => x"75",
          3702 => x"fc",
          3703 => x"9c",
          3704 => x"70",
          3705 => x"80",
          3706 => x"84",
          3707 => x"79",
          3708 => x"f4",
          3709 => x"10",
          3710 => x"05",
          3711 => x"43",
          3712 => x"52",
          3713 => x"83",
          3714 => x"f4",
          3715 => x"10",
          3716 => x"05",
          3717 => x"5e",
          3718 => x"cf",
          3719 => x"ec",
          3720 => x"80",
          3721 => x"83",
          3722 => x"58",
          3723 => x"8b",
          3724 => x"0b",
          3725 => x"34",
          3726 => x"e2",
          3727 => x"84",
          3728 => x"b5",
          3729 => x"84",
          3730 => x"55",
          3731 => x"b6",
          3732 => x"e8",
          3733 => x"51",
          3734 => x"3f",
          3735 => x"08",
          3736 => x"ff",
          3737 => x"84",
          3738 => x"52",
          3739 => x"ae",
          3740 => x"e2",
          3741 => x"05",
          3742 => x"e2",
          3743 => x"81",
          3744 => x"74",
          3745 => x"d3",
          3746 => x"9e",
          3747 => x"0b",
          3748 => x"34",
          3749 => x"e2",
          3750 => x"e4",
          3751 => x"c8",
          3752 => x"ff",
          3753 => x"7a",
          3754 => x"d4",
          3755 => x"c4",
          3756 => x"5a",
          3757 => x"c4",
          3758 => x"58",
          3759 => x"c8",
          3760 => x"e8",
          3761 => x"51",
          3762 => x"3f",
          3763 => x"33",
          3764 => x"70",
          3765 => x"e2",
          3766 => x"52",
          3767 => x"76",
          3768 => x"38",
          3769 => x"08",
          3770 => x"ff",
          3771 => x"84",
          3772 => x"70",
          3773 => x"98",
          3774 => x"c4",
          3775 => x"59",
          3776 => x"24",
          3777 => x"84",
          3778 => x"52",
          3779 => x"ac",
          3780 => x"81",
          3781 => x"81",
          3782 => x"70",
          3783 => x"e2",
          3784 => x"51",
          3785 => x"24",
          3786 => x"84",
          3787 => x"52",
          3788 => x"ac",
          3789 => x"81",
          3790 => x"81",
          3791 => x"70",
          3792 => x"e2",
          3793 => x"51",
          3794 => x"25",
          3795 => x"f3",
          3796 => x"16",
          3797 => x"33",
          3798 => x"e6",
          3799 => x"76",
          3800 => x"ac",
          3801 => x"81",
          3802 => x"81",
          3803 => x"70",
          3804 => x"e2",
          3805 => x"57",
          3806 => x"25",
          3807 => x"7b",
          3808 => x"17",
          3809 => x"84",
          3810 => x"52",
          3811 => x"ff",
          3812 => x"75",
          3813 => x"29",
          3814 => x"05",
          3815 => x"84",
          3816 => x"44",
          3817 => x"76",
          3818 => x"38",
          3819 => x"83",
          3820 => x"0b",
          3821 => x"84",
          3822 => x"55",
          3823 => x"b6",
          3824 => x"e8",
          3825 => x"51",
          3826 => x"3f",
          3827 => x"08",
          3828 => x"ff",
          3829 => x"84",
          3830 => x"52",
          3831 => x"ab",
          3832 => x"e2",
          3833 => x"05",
          3834 => x"e2",
          3835 => x"81",
          3836 => x"74",
          3837 => x"d3",
          3838 => x"9c",
          3839 => x"0b",
          3840 => x"34",
          3841 => x"e2",
          3842 => x"84",
          3843 => x"b5",
          3844 => x"84",
          3845 => x"70",
          3846 => x"58",
          3847 => x"2e",
          3848 => x"84",
          3849 => x"55",
          3850 => x"ae",
          3851 => x"2b",
          3852 => x"57",
          3853 => x"24",
          3854 => x"16",
          3855 => x"81",
          3856 => x"81",
          3857 => x"81",
          3858 => x"70",
          3859 => x"e2",
          3860 => x"57",
          3861 => x"25",
          3862 => x"18",
          3863 => x"e2",
          3864 => x"81",
          3865 => x"05",
          3866 => x"33",
          3867 => x"e2",
          3868 => x"76",
          3869 => x"38",
          3870 => x"75",
          3871 => x"34",
          3872 => x"e2",
          3873 => x"81",
          3874 => x"81",
          3875 => x"70",
          3876 => x"81",
          3877 => x"58",
          3878 => x"76",
          3879 => x"38",
          3880 => x"70",
          3881 => x"81",
          3882 => x"57",
          3883 => x"25",
          3884 => x"84",
          3885 => x"52",
          3886 => x"a9",
          3887 => x"81",
          3888 => x"81",
          3889 => x"70",
          3890 => x"e2",
          3891 => x"57",
          3892 => x"25",
          3893 => x"84",
          3894 => x"52",
          3895 => x"a9",
          3896 => x"81",
          3897 => x"81",
          3898 => x"70",
          3899 => x"e2",
          3900 => x"57",
          3901 => x"24",
          3902 => x"f0",
          3903 => x"a8",
          3904 => x"c8",
          3905 => x"84",
          3906 => x"ec",
          3907 => x"84",
          3908 => x"e2",
          3909 => x"99",
          3910 => x"f4",
          3911 => x"74",
          3912 => x"75",
          3913 => x"34",
          3914 => x"38",
          3915 => x"84",
          3916 => x"52",
          3917 => x"33",
          3918 => x"a8",
          3919 => x"81",
          3920 => x"81",
          3921 => x"70",
          3922 => x"e2",
          3923 => x"57",
          3924 => x"24",
          3925 => x"e2",
          3926 => x"98",
          3927 => x"2c",
          3928 => x"06",
          3929 => x"58",
          3930 => x"ef",
          3931 => x"c3",
          3932 => x"ec",
          3933 => x"ef",
          3934 => x"f4",
          3935 => x"56",
          3936 => x"74",
          3937 => x"16",
          3938 => x"56",
          3939 => x"f0",
          3940 => x"83",
          3941 => x"83",
          3942 => x"55",
          3943 => x"ee",
          3944 => x"51",
          3945 => x"3f",
          3946 => x"08",
          3947 => x"ac",
          3948 => x"83",
          3949 => x"94",
          3950 => x"40",
          3951 => x"39",
          3952 => x"db",
          3953 => x"77",
          3954 => x"84",
          3955 => x"75",
          3956 => x"ac",
          3957 => x"39",
          3958 => x"aa",
          3959 => x"bb",
          3960 => x"e2",
          3961 => x"bb",
          3962 => x"ff",
          3963 => x"53",
          3964 => x"51",
          3965 => x"3f",
          3966 => x"e2",
          3967 => x"e2",
          3968 => x"57",
          3969 => x"2e",
          3970 => x"84",
          3971 => x"52",
          3972 => x"a6",
          3973 => x"e6",
          3974 => x"a0",
          3975 => x"d1",
          3976 => x"e8",
          3977 => x"51",
          3978 => x"3f",
          3979 => x"33",
          3980 => x"78",
          3981 => x"34",
          3982 => x"06",
          3983 => x"75",
          3984 => x"e7",
          3985 => x"84",
          3986 => x"c4",
          3987 => x"84",
          3988 => x"06",
          3989 => x"75",
          3990 => x"ff",
          3991 => x"76",
          3992 => x"33",
          3993 => x"33",
          3994 => x"74",
          3995 => x"de",
          3996 => x"e8",
          3997 => x"51",
          3998 => x"3f",
          3999 => x"08",
          4000 => x"ff",
          4001 => x"84",
          4002 => x"52",
          4003 => x"a5",
          4004 => x"e2",
          4005 => x"05",
          4006 => x"e2",
          4007 => x"81",
          4008 => x"c7",
          4009 => x"ff",
          4010 => x"84",
          4011 => x"84",
          4012 => x"84",
          4013 => x"81",
          4014 => x"05",
          4015 => x"7b",
          4016 => x"a9",
          4017 => x"70",
          4018 => x"84",
          4019 => x"84",
          4020 => x"58",
          4021 => x"74",
          4022 => x"f2",
          4023 => x"e8",
          4024 => x"51",
          4025 => x"3f",
          4026 => x"08",
          4027 => x"ff",
          4028 => x"84",
          4029 => x"52",
          4030 => x"a4",
          4031 => x"e2",
          4032 => x"05",
          4033 => x"e2",
          4034 => x"81",
          4035 => x"c7",
          4036 => x"34",
          4037 => x"e2",
          4038 => x"0b",
          4039 => x"34",
          4040 => x"84",
          4041 => x"0d",
          4042 => x"9c",
          4043 => x"80",
          4044 => x"38",
          4045 => x"a7",
          4046 => x"bb",
          4047 => x"e2",
          4048 => x"bb",
          4049 => x"ff",
          4050 => x"53",
          4051 => x"51",
          4052 => x"3f",
          4053 => x"33",
          4054 => x"33",
          4055 => x"80",
          4056 => x"38",
          4057 => x"08",
          4058 => x"ff",
          4059 => x"84",
          4060 => x"52",
          4061 => x"a3",
          4062 => x"e6",
          4063 => x"88",
          4064 => x"ed",
          4065 => x"c8",
          4066 => x"59",
          4067 => x"c8",
          4068 => x"ff",
          4069 => x"39",
          4070 => x"d7",
          4071 => x"f4",
          4072 => x"82",
          4073 => x"06",
          4074 => x"05",
          4075 => x"54",
          4076 => x"80",
          4077 => x"84",
          4078 => x"79",
          4079 => x"f4",
          4080 => x"10",
          4081 => x"05",
          4082 => x"43",
          4083 => x"52",
          4084 => x"b7",
          4085 => x"f4",
          4086 => x"10",
          4087 => x"05",
          4088 => x"5e",
          4089 => x"2e",
          4090 => x"75",
          4091 => x"74",
          4092 => x"f9",
          4093 => x"f4",
          4094 => x"70",
          4095 => x"56",
          4096 => x"27",
          4097 => x"77",
          4098 => x"34",
          4099 => x"b5",
          4100 => x"05",
          4101 => x"7b",
          4102 => x"81",
          4103 => x"83",
          4104 => x"52",
          4105 => x"b9",
          4106 => x"f4",
          4107 => x"81",
          4108 => x"80",
          4109 => x"c8",
          4110 => x"84",
          4111 => x"7b",
          4112 => x"0c",
          4113 => x"04",
          4114 => x"52",
          4115 => x"ca",
          4116 => x"bb",
          4117 => x"d5",
          4118 => x"84",
          4119 => x"5c",
          4120 => x"ec",
          4121 => x"f8",
          4122 => x"82",
          4123 => x"84",
          4124 => x"5a",
          4125 => x"08",
          4126 => x"81",
          4127 => x"38",
          4128 => x"08",
          4129 => x"a3",
          4130 => x"84",
          4131 => x"0b",
          4132 => x"08",
          4133 => x"38",
          4134 => x"08",
          4135 => x"1b",
          4136 => x"76",
          4137 => x"ff",
          4138 => x"f4",
          4139 => x"10",
          4140 => x"05",
          4141 => x"41",
          4142 => x"81",
          4143 => x"82",
          4144 => x"06",
          4145 => x"05",
          4146 => x"53",
          4147 => x"da",
          4148 => x"bb",
          4149 => x"0c",
          4150 => x"33",
          4151 => x"83",
          4152 => x"70",
          4153 => x"83",
          4154 => x"59",
          4155 => x"3f",
          4156 => x"33",
          4157 => x"83",
          4158 => x"70",
          4159 => x"42",
          4160 => x"81",
          4161 => x"ff",
          4162 => x"93",
          4163 => x"38",
          4164 => x"ff",
          4165 => x"06",
          4166 => x"77",
          4167 => x"f8",
          4168 => x"53",
          4169 => x"51",
          4170 => x"3f",
          4171 => x"33",
          4172 => x"81",
          4173 => x"56",
          4174 => x"80",
          4175 => x"0b",
          4176 => x"34",
          4177 => x"74",
          4178 => x"90",
          4179 => x"f4",
          4180 => x"2b",
          4181 => x"83",
          4182 => x"81",
          4183 => x"52",
          4184 => x"d9",
          4185 => x"bb",
          4186 => x"0c",
          4187 => x"33",
          4188 => x"83",
          4189 => x"70",
          4190 => x"83",
          4191 => x"59",
          4192 => x"3f",
          4193 => x"33",
          4194 => x"83",
          4195 => x"70",
          4196 => x"42",
          4197 => x"fe",
          4198 => x"86",
          4199 => x"f4",
          4200 => x"df",
          4201 => x"f4",
          4202 => x"f1",
          4203 => x"d4",
          4204 => x"c2",
          4205 => x"c2",
          4206 => x"39",
          4207 => x"02",
          4208 => x"33",
          4209 => x"80",
          4210 => x"5b",
          4211 => x"26",
          4212 => x"72",
          4213 => x"8b",
          4214 => x"25",
          4215 => x"72",
          4216 => x"a8",
          4217 => x"a0",
          4218 => x"c7",
          4219 => x"5e",
          4220 => x"9f",
          4221 => x"76",
          4222 => x"75",
          4223 => x"34",
          4224 => x"b5",
          4225 => x"fa",
          4226 => x"fa",
          4227 => x"98",
          4228 => x"2b",
          4229 => x"2b",
          4230 => x"7a",
          4231 => x"56",
          4232 => x"27",
          4233 => x"74",
          4234 => x"56",
          4235 => x"70",
          4236 => x"0c",
          4237 => x"ee",
          4238 => x"27",
          4239 => x"fa",
          4240 => x"99",
          4241 => x"78",
          4242 => x"55",
          4243 => x"e0",
          4244 => x"74",
          4245 => x"56",
          4246 => x"53",
          4247 => x"90",
          4248 => x"86",
          4249 => x"0b",
          4250 => x"33",
          4251 => x"11",
          4252 => x"33",
          4253 => x"11",
          4254 => x"41",
          4255 => x"86",
          4256 => x"0b",
          4257 => x"33",
          4258 => x"06",
          4259 => x"33",
          4260 => x"06",
          4261 => x"22",
          4262 => x"ff",
          4263 => x"29",
          4264 => x"58",
          4265 => x"5d",
          4266 => x"87",
          4267 => x"31",
          4268 => x"79",
          4269 => x"7e",
          4270 => x"7c",
          4271 => x"7a",
          4272 => x"06",
          4273 => x"06",
          4274 => x"14",
          4275 => x"57",
          4276 => x"74",
          4277 => x"83",
          4278 => x"74",
          4279 => x"70",
          4280 => x"59",
          4281 => x"06",
          4282 => x"2e",
          4283 => x"78",
          4284 => x"72",
          4285 => x"c1",
          4286 => x"70",
          4287 => x"34",
          4288 => x"33",
          4289 => x"05",
          4290 => x"39",
          4291 => x"80",
          4292 => x"b0",
          4293 => x"b8",
          4294 => x"81",
          4295 => x"b8",
          4296 => x"81",
          4297 => x"fa",
          4298 => x"74",
          4299 => x"5d",
          4300 => x"5e",
          4301 => x"27",
          4302 => x"73",
          4303 => x"73",
          4304 => x"71",
          4305 => x"5a",
          4306 => x"80",
          4307 => x"38",
          4308 => x"fa",
          4309 => x"0b",
          4310 => x"34",
          4311 => x"33",
          4312 => x"71",
          4313 => x"71",
          4314 => x"71",
          4315 => x"56",
          4316 => x"76",
          4317 => x"ae",
          4318 => x"39",
          4319 => x"38",
          4320 => x"33",
          4321 => x"06",
          4322 => x"11",
          4323 => x"33",
          4324 => x"11",
          4325 => x"80",
          4326 => x"5b",
          4327 => x"86",
          4328 => x"70",
          4329 => x"f8",
          4330 => x"ff",
          4331 => x"f7",
          4332 => x"ff",
          4333 => x"b2",
          4334 => x"ff",
          4335 => x"75",
          4336 => x"5e",
          4337 => x"58",
          4338 => x"57",
          4339 => x"8b",
          4340 => x"31",
          4341 => x"29",
          4342 => x"7d",
          4343 => x"74",
          4344 => x"71",
          4345 => x"83",
          4346 => x"62",
          4347 => x"70",
          4348 => x"5f",
          4349 => x"55",
          4350 => x"85",
          4351 => x"29",
          4352 => x"31",
          4353 => x"06",
          4354 => x"fd",
          4355 => x"83",
          4356 => x"fd",
          4357 => x"f2",
          4358 => x"31",
          4359 => x"fe",
          4360 => x"3d",
          4361 => x"80",
          4362 => x"8a",
          4363 => x"73",
          4364 => x"34",
          4365 => x"87",
          4366 => x"55",
          4367 => x"34",
          4368 => x"34",
          4369 => x"98",
          4370 => x"34",
          4371 => x"87",
          4372 => x"54",
          4373 => x"80",
          4374 => x"80",
          4375 => x"52",
          4376 => x"d8",
          4377 => x"87",
          4378 => x"54",
          4379 => x"56",
          4380 => x"f8",
          4381 => x"84",
          4382 => x"72",
          4383 => x"08",
          4384 => x"06",
          4385 => x"51",
          4386 => x"34",
          4387 => x"cc",
          4388 => x"06",
          4389 => x"53",
          4390 => x"81",
          4391 => x"08",
          4392 => x"88",
          4393 => x"75",
          4394 => x"0b",
          4395 => x"34",
          4396 => x"bb",
          4397 => x"3d",
          4398 => x"b8",
          4399 => x"bb",
          4400 => x"f7",
          4401 => x"af",
          4402 => x"84",
          4403 => x"33",
          4404 => x"33",
          4405 => x"81",
          4406 => x"26",
          4407 => x"84",
          4408 => x"83",
          4409 => x"83",
          4410 => x"72",
          4411 => x"86",
          4412 => x"11",
          4413 => x"22",
          4414 => x"59",
          4415 => x"05",
          4416 => x"ff",
          4417 => x"8a",
          4418 => x"58",
          4419 => x"2e",
          4420 => x"83",
          4421 => x"76",
          4422 => x"83",
          4423 => x"83",
          4424 => x"76",
          4425 => x"ff",
          4426 => x"ff",
          4427 => x"55",
          4428 => x"82",
          4429 => x"19",
          4430 => x"fa",
          4431 => x"fa",
          4432 => x"83",
          4433 => x"84",
          4434 => x"5c",
          4435 => x"74",
          4436 => x"38",
          4437 => x"33",
          4438 => x"54",
          4439 => x"72",
          4440 => x"ac",
          4441 => x"d6",
          4442 => x"55",
          4443 => x"33",
          4444 => x"34",
          4445 => x"05",
          4446 => x"70",
          4447 => x"34",
          4448 => x"84",
          4449 => x"27",
          4450 => x"9f",
          4451 => x"38",
          4452 => x"33",
          4453 => x"15",
          4454 => x"0b",
          4455 => x"34",
          4456 => x"81",
          4457 => x"81",
          4458 => x"9f",
          4459 => x"38",
          4460 => x"33",
          4461 => x"75",
          4462 => x"23",
          4463 => x"81",
          4464 => x"83",
          4465 => x"54",
          4466 => x"26",
          4467 => x"72",
          4468 => x"05",
          4469 => x"33",
          4470 => x"58",
          4471 => x"55",
          4472 => x"80",
          4473 => x"b0",
          4474 => x"ff",
          4475 => x"ff",
          4476 => x"29",
          4477 => x"54",
          4478 => x"27",
          4479 => x"99",
          4480 => x"e0",
          4481 => x"53",
          4482 => x"13",
          4483 => x"81",
          4484 => x"73",
          4485 => x"55",
          4486 => x"81",
          4487 => x"81",
          4488 => x"f8",
          4489 => x"f7",
          4490 => x"29",
          4491 => x"5a",
          4492 => x"26",
          4493 => x"53",
          4494 => x"84",
          4495 => x"0d",
          4496 => x"fa",
          4497 => x"fa",
          4498 => x"83",
          4499 => x"84",
          4500 => x"5c",
          4501 => x"7a",
          4502 => x"38",
          4503 => x"fe",
          4504 => x"81",
          4505 => x"05",
          4506 => x"33",
          4507 => x"75",
          4508 => x"06",
          4509 => x"73",
          4510 => x"05",
          4511 => x"33",
          4512 => x"78",
          4513 => x"56",
          4514 => x"73",
          4515 => x"ae",
          4516 => x"b0",
          4517 => x"d6",
          4518 => x"31",
          4519 => x"a0",
          4520 => x"16",
          4521 => x"70",
          4522 => x"34",
          4523 => x"72",
          4524 => x"8a",
          4525 => x"e0",
          4526 => x"75",
          4527 => x"05",
          4528 => x"13",
          4529 => x"38",
          4530 => x"80",
          4531 => x"f8",
          4532 => x"fe",
          4533 => x"fa",
          4534 => x"59",
          4535 => x"19",
          4536 => x"84",
          4537 => x"59",
          4538 => x"fc",
          4539 => x"02",
          4540 => x"05",
          4541 => x"70",
          4542 => x"38",
          4543 => x"83",
          4544 => x"51",
          4545 => x"84",
          4546 => x"51",
          4547 => x"86",
          4548 => x"fa",
          4549 => x"0b",
          4550 => x"0c",
          4551 => x"04",
          4552 => x"fa",
          4553 => x"fa",
          4554 => x"81",
          4555 => x"52",
          4556 => x"e2",
          4557 => x"51",
          4558 => x"b4",
          4559 => x"84",
          4560 => x"86",
          4561 => x"83",
          4562 => x"70",
          4563 => x"09",
          4564 => x"72",
          4565 => x"53",
          4566 => x"fa",
          4567 => x"39",
          4568 => x"33",
          4569 => x"b8",
          4570 => x"11",
          4571 => x"70",
          4572 => x"38",
          4573 => x"83",
          4574 => x"80",
          4575 => x"84",
          4576 => x"0d",
          4577 => x"b5",
          4578 => x"31",
          4579 => x"9f",
          4580 => x"54",
          4581 => x"70",
          4582 => x"34",
          4583 => x"bb",
          4584 => x"3d",
          4585 => x"fa",
          4586 => x"05",
          4587 => x"33",
          4588 => x"55",
          4589 => x"25",
          4590 => x"53",
          4591 => x"b5",
          4592 => x"84",
          4593 => x"86",
          4594 => x"80",
          4595 => x"b5",
          4596 => x"b4",
          4597 => x"f7",
          4598 => x"56",
          4599 => x"25",
          4600 => x"81",
          4601 => x"83",
          4602 => x"fe",
          4603 => x"3d",
          4604 => x"05",
          4605 => x"b1",
          4606 => x"70",
          4607 => x"c5",
          4608 => x"70",
          4609 => x"fa",
          4610 => x"80",
          4611 => x"84",
          4612 => x"06",
          4613 => x"2a",
          4614 => x"53",
          4615 => x"f0",
          4616 => x"06",
          4617 => x"f2",
          4618 => x"b0",
          4619 => x"84",
          4620 => x"83",
          4621 => x"83",
          4622 => x"81",
          4623 => x"07",
          4624 => x"fa",
          4625 => x"0b",
          4626 => x"0c",
          4627 => x"04",
          4628 => x"33",
          4629 => x"51",
          4630 => x"b0",
          4631 => x"83",
          4632 => x"81",
          4633 => x"07",
          4634 => x"fa",
          4635 => x"39",
          4636 => x"83",
          4637 => x"80",
          4638 => x"84",
          4639 => x"0d",
          4640 => x"b0",
          4641 => x"06",
          4642 => x"70",
          4643 => x"34",
          4644 => x"83",
          4645 => x"87",
          4646 => x"83",
          4647 => x"ff",
          4648 => x"fa",
          4649 => x"fd",
          4650 => x"51",
          4651 => x"b0",
          4652 => x"39",
          4653 => x"33",
          4654 => x"83",
          4655 => x"83",
          4656 => x"ff",
          4657 => x"fa",
          4658 => x"f9",
          4659 => x"51",
          4660 => x"b0",
          4661 => x"39",
          4662 => x"33",
          4663 => x"51",
          4664 => x"b0",
          4665 => x"39",
          4666 => x"33",
          4667 => x"80",
          4668 => x"70",
          4669 => x"34",
          4670 => x"83",
          4671 => x"81",
          4672 => x"07",
          4673 => x"fa",
          4674 => x"ba",
          4675 => x"b0",
          4676 => x"06",
          4677 => x"51",
          4678 => x"b0",
          4679 => x"39",
          4680 => x"33",
          4681 => x"80",
          4682 => x"70",
          4683 => x"34",
          4684 => x"83",
          4685 => x"81",
          4686 => x"07",
          4687 => x"fa",
          4688 => x"82",
          4689 => x"b0",
          4690 => x"06",
          4691 => x"fa",
          4692 => x"f2",
          4693 => x"b0",
          4694 => x"06",
          4695 => x"70",
          4696 => x"34",
          4697 => x"f3",
          4698 => x"bf",
          4699 => x"84",
          4700 => x"05",
          4701 => x"b4",
          4702 => x"b3",
          4703 => x"b5",
          4704 => x"fa",
          4705 => x"5f",
          4706 => x"78",
          4707 => x"a1",
          4708 => x"24",
          4709 => x"81",
          4710 => x"38",
          4711 => x"fa",
          4712 => x"84",
          4713 => x"7a",
          4714 => x"34",
          4715 => x"b2",
          4716 => x"fa",
          4717 => x"3d",
          4718 => x"83",
          4719 => x"06",
          4720 => x"0b",
          4721 => x"34",
          4722 => x"b8",
          4723 => x"0b",
          4724 => x"34",
          4725 => x"fa",
          4726 => x"0b",
          4727 => x"23",
          4728 => x"b8",
          4729 => x"84",
          4730 => x"56",
          4731 => x"33",
          4732 => x"7c",
          4733 => x"83",
          4734 => x"ff",
          4735 => x"7d",
          4736 => x"34",
          4737 => x"b8",
          4738 => x"83",
          4739 => x"7b",
          4740 => x"23",
          4741 => x"b5",
          4742 => x"0d",
          4743 => x"84",
          4744 => x"81",
          4745 => x"fc",
          4746 => x"83",
          4747 => x"a8",
          4748 => x"b5",
          4749 => x"83",
          4750 => x"84",
          4751 => x"58",
          4752 => x"33",
          4753 => x"85",
          4754 => x"55",
          4755 => x"53",
          4756 => x"e5",
          4757 => x"ff",
          4758 => x"0b",
          4759 => x"33",
          4760 => x"79",
          4761 => x"79",
          4762 => x"d8",
          4763 => x"53",
          4764 => x"ac",
          4765 => x"93",
          4766 => x"70",
          4767 => x"84",
          4768 => x"52",
          4769 => x"7a",
          4770 => x"83",
          4771 => x"fe",
          4772 => x"7d",
          4773 => x"34",
          4774 => x"b8",
          4775 => x"83",
          4776 => x"7b",
          4777 => x"23",
          4778 => x"b5",
          4779 => x"0d",
          4780 => x"84",
          4781 => x"81",
          4782 => x"fc",
          4783 => x"83",
          4784 => x"a8",
          4785 => x"b5",
          4786 => x"83",
          4787 => x"83",
          4788 => x"ff",
          4789 => x"84",
          4790 => x"52",
          4791 => x"51",
          4792 => x"3f",
          4793 => x"f8",
          4794 => x"90",
          4795 => x"84",
          4796 => x"27",
          4797 => x"83",
          4798 => x"33",
          4799 => x"b8",
          4800 => x"87",
          4801 => x"70",
          4802 => x"5a",
          4803 => x"f9",
          4804 => x"02",
          4805 => x"05",
          4806 => x"f8",
          4807 => x"b5",
          4808 => x"b4",
          4809 => x"29",
          4810 => x"a0",
          4811 => x"fa",
          4812 => x"51",
          4813 => x"7c",
          4814 => x"83",
          4815 => x"83",
          4816 => x"52",
          4817 => x"57",
          4818 => x"2e",
          4819 => x"75",
          4820 => x"f9",
          4821 => x"24",
          4822 => x"75",
          4823 => x"85",
          4824 => x"2e",
          4825 => x"84",
          4826 => x"83",
          4827 => x"83",
          4828 => x"72",
          4829 => x"55",
          4830 => x"b9",
          4831 => x"86",
          4832 => x"14",
          4833 => x"f8",
          4834 => x"b5",
          4835 => x"b2",
          4836 => x"29",
          4837 => x"56",
          4838 => x"fa",
          4839 => x"83",
          4840 => x"73",
          4841 => x"58",
          4842 => x"b0",
          4843 => x"b0",
          4844 => x"84",
          4845 => x"70",
          4846 => x"83",
          4847 => x"83",
          4848 => x"72",
          4849 => x"57",
          4850 => x"57",
          4851 => x"33",
          4852 => x"14",
          4853 => x"70",
          4854 => x"59",
          4855 => x"26",
          4856 => x"84",
          4857 => x"58",
          4858 => x"38",
          4859 => x"72",
          4860 => x"34",
          4861 => x"33",
          4862 => x"2e",
          4863 => x"b8",
          4864 => x"76",
          4865 => x"fb",
          4866 => x"84",
          4867 => x"89",
          4868 => x"75",
          4869 => x"38",
          4870 => x"80",
          4871 => x"8a",
          4872 => x"06",
          4873 => x"81",
          4874 => x"f1",
          4875 => x"0b",
          4876 => x"34",
          4877 => x"83",
          4878 => x"33",
          4879 => x"80",
          4880 => x"34",
          4881 => x"09",
          4882 => x"89",
          4883 => x"76",
          4884 => x"fd",
          4885 => x"13",
          4886 => x"06",
          4887 => x"83",
          4888 => x"38",
          4889 => x"51",
          4890 => x"81",
          4891 => x"ff",
          4892 => x"83",
          4893 => x"38",
          4894 => x"74",
          4895 => x"34",
          4896 => x"75",
          4897 => x"f9",
          4898 => x"0b",
          4899 => x"0c",
          4900 => x"04",
          4901 => x"2e",
          4902 => x"fd",
          4903 => x"fa",
          4904 => x"81",
          4905 => x"ff",
          4906 => x"83",
          4907 => x"72",
          4908 => x"34",
          4909 => x"51",
          4910 => x"83",
          4911 => x"70",
          4912 => x"55",
          4913 => x"73",
          4914 => x"73",
          4915 => x"fa",
          4916 => x"a0",
          4917 => x"83",
          4918 => x"81",
          4919 => x"ef",
          4920 => x"90",
          4921 => x"75",
          4922 => x"3f",
          4923 => x"e6",
          4924 => x"80",
          4925 => x"84",
          4926 => x"57",
          4927 => x"2e",
          4928 => x"75",
          4929 => x"82",
          4930 => x"2e",
          4931 => x"78",
          4932 => x"d1",
          4933 => x"2e",
          4934 => x"78",
          4935 => x"8f",
          4936 => x"f8",
          4937 => x"b4",
          4938 => x"b5",
          4939 => x"29",
          4940 => x"5c",
          4941 => x"19",
          4942 => x"a0",
          4943 => x"84",
          4944 => x"83",
          4945 => x"83",
          4946 => x"72",
          4947 => x"5a",
          4948 => x"78",
          4949 => x"18",
          4950 => x"b4",
          4951 => x"29",
          4952 => x"5a",
          4953 => x"33",
          4954 => x"b0",
          4955 => x"84",
          4956 => x"70",
          4957 => x"83",
          4958 => x"83",
          4959 => x"72",
          4960 => x"42",
          4961 => x"59",
          4962 => x"33",
          4963 => x"1f",
          4964 => x"70",
          4965 => x"42",
          4966 => x"26",
          4967 => x"84",
          4968 => x"5a",
          4969 => x"38",
          4970 => x"75",
          4971 => x"34",
          4972 => x"bb",
          4973 => x"3d",
          4974 => x"b7",
          4975 => x"38",
          4976 => x"81",
          4977 => x"b8",
          4978 => x"38",
          4979 => x"2e",
          4980 => x"80",
          4981 => x"80",
          4982 => x"f8",
          4983 => x"b4",
          4984 => x"b5",
          4985 => x"29",
          4986 => x"40",
          4987 => x"19",
          4988 => x"a0",
          4989 => x"84",
          4990 => x"83",
          4991 => x"83",
          4992 => x"72",
          4993 => x"41",
          4994 => x"78",
          4995 => x"1f",
          4996 => x"b4",
          4997 => x"29",
          4998 => x"83",
          4999 => x"86",
          5000 => x"1b",
          5001 => x"f8",
          5002 => x"ff",
          5003 => x"b2",
          5004 => x"b5",
          5005 => x"29",
          5006 => x"43",
          5007 => x"fa",
          5008 => x"84",
          5009 => x"34",
          5010 => x"77",
          5011 => x"41",
          5012 => x"fe",
          5013 => x"83",
          5014 => x"80",
          5015 => x"84",
          5016 => x"0d",
          5017 => x"2e",
          5018 => x"78",
          5019 => x"81",
          5020 => x"2e",
          5021 => x"fd",
          5022 => x"0b",
          5023 => x"34",
          5024 => x"bb",
          5025 => x"3d",
          5026 => x"9b",
          5027 => x"38",
          5028 => x"75",
          5029 => x"d0",
          5030 => x"84",
          5031 => x"59",
          5032 => x"ba",
          5033 => x"84",
          5034 => x"34",
          5035 => x"06",
          5036 => x"84",
          5037 => x"34",
          5038 => x"bb",
          5039 => x"3d",
          5040 => x"9b",
          5041 => x"38",
          5042 => x"ba",
          5043 => x"b8",
          5044 => x"fa",
          5045 => x"fa",
          5046 => x"72",
          5047 => x"40",
          5048 => x"80",
          5049 => x"c7",
          5050 => x"34",
          5051 => x"33",
          5052 => x"33",
          5053 => x"22",
          5054 => x"12",
          5055 => x"56",
          5056 => x"b6",
          5057 => x"fa",
          5058 => x"71",
          5059 => x"57",
          5060 => x"33",
          5061 => x"80",
          5062 => x"b8",
          5063 => x"81",
          5064 => x"fa",
          5065 => x"fa",
          5066 => x"72",
          5067 => x"42",
          5068 => x"83",
          5069 => x"60",
          5070 => x"05",
          5071 => x"58",
          5072 => x"81",
          5073 => x"ea",
          5074 => x"0b",
          5075 => x"34",
          5076 => x"84",
          5077 => x"83",
          5078 => x"70",
          5079 => x"83",
          5080 => x"73",
          5081 => x"86",
          5082 => x"05",
          5083 => x"22",
          5084 => x"72",
          5085 => x"70",
          5086 => x"06",
          5087 => x"33",
          5088 => x"5a",
          5089 => x"2e",
          5090 => x"78",
          5091 => x"ff",
          5092 => x"76",
          5093 => x"76",
          5094 => x"fa",
          5095 => x"90",
          5096 => x"84",
          5097 => x"80",
          5098 => x"85",
          5099 => x"84",
          5100 => x"80",
          5101 => x"87",
          5102 => x"84",
          5103 => x"80",
          5104 => x"84",
          5105 => x"0d",
          5106 => x"b4",
          5107 => x"ec",
          5108 => x"b5",
          5109 => x"ed",
          5110 => x"b3",
          5111 => x"ee",
          5112 => x"84",
          5113 => x"80",
          5114 => x"84",
          5115 => x"0d",
          5116 => x"ff",
          5117 => x"06",
          5118 => x"83",
          5119 => x"84",
          5120 => x"70",
          5121 => x"83",
          5122 => x"70",
          5123 => x"72",
          5124 => x"86",
          5125 => x"05",
          5126 => x"22",
          5127 => x"7b",
          5128 => x"83",
          5129 => x"83",
          5130 => x"44",
          5131 => x"42",
          5132 => x"81",
          5133 => x"38",
          5134 => x"06",
          5135 => x"56",
          5136 => x"75",
          5137 => x"fa",
          5138 => x"81",
          5139 => x"81",
          5140 => x"81",
          5141 => x"72",
          5142 => x"40",
          5143 => x"a0",
          5144 => x"a0",
          5145 => x"84",
          5146 => x"83",
          5147 => x"83",
          5148 => x"72",
          5149 => x"5a",
          5150 => x"a0",
          5151 => x"b6",
          5152 => x"fa",
          5153 => x"71",
          5154 => x"5a",
          5155 => x"b0",
          5156 => x"b0",
          5157 => x"84",
          5158 => x"70",
          5159 => x"83",
          5160 => x"83",
          5161 => x"72",
          5162 => x"43",
          5163 => x"59",
          5164 => x"33",
          5165 => x"d6",
          5166 => x"1a",
          5167 => x"06",
          5168 => x"7b",
          5169 => x"38",
          5170 => x"33",
          5171 => x"d0",
          5172 => x"58",
          5173 => x"b5",
          5174 => x"b5",
          5175 => x"ff",
          5176 => x"05",
          5177 => x"39",
          5178 => x"95",
          5179 => x"bd",
          5180 => x"38",
          5181 => x"95",
          5182 => x"ba",
          5183 => x"7e",
          5184 => x"ff",
          5185 => x"75",
          5186 => x"c8",
          5187 => x"10",
          5188 => x"05",
          5189 => x"04",
          5190 => x"fa",
          5191 => x"52",
          5192 => x"9f",
          5193 => x"84",
          5194 => x"9c",
          5195 => x"83",
          5196 => x"84",
          5197 => x"70",
          5198 => x"83",
          5199 => x"70",
          5200 => x"72",
          5201 => x"86",
          5202 => x"05",
          5203 => x"22",
          5204 => x"7b",
          5205 => x"83",
          5206 => x"83",
          5207 => x"46",
          5208 => x"59",
          5209 => x"81",
          5210 => x"38",
          5211 => x"81",
          5212 => x"81",
          5213 => x"81",
          5214 => x"72",
          5215 => x"58",
          5216 => x"a0",
          5217 => x"a0",
          5218 => x"84",
          5219 => x"83",
          5220 => x"83",
          5221 => x"72",
          5222 => x"5e",
          5223 => x"a0",
          5224 => x"b6",
          5225 => x"fa",
          5226 => x"71",
          5227 => x"5e",
          5228 => x"33",
          5229 => x"80",
          5230 => x"b8",
          5231 => x"81",
          5232 => x"fa",
          5233 => x"fa",
          5234 => x"72",
          5235 => x"44",
          5236 => x"83",
          5237 => x"84",
          5238 => x"34",
          5239 => x"70",
          5240 => x"5b",
          5241 => x"26",
          5242 => x"84",
          5243 => x"58",
          5244 => x"38",
          5245 => x"75",
          5246 => x"34",
          5247 => x"81",
          5248 => x"59",
          5249 => x"f7",
          5250 => x"fa",
          5251 => x"b8",
          5252 => x"fa",
          5253 => x"81",
          5254 => x"81",
          5255 => x"81",
          5256 => x"72",
          5257 => x"5b",
          5258 => x"5b",
          5259 => x"33",
          5260 => x"80",
          5261 => x"b8",
          5262 => x"fa",
          5263 => x"fa",
          5264 => x"71",
          5265 => x"41",
          5266 => x"0b",
          5267 => x"1c",
          5268 => x"b4",
          5269 => x"29",
          5270 => x"83",
          5271 => x"86",
          5272 => x"1a",
          5273 => x"f8",
          5274 => x"ff",
          5275 => x"b2",
          5276 => x"b5",
          5277 => x"29",
          5278 => x"5a",
          5279 => x"fa",
          5280 => x"99",
          5281 => x"60",
          5282 => x"81",
          5283 => x"58",
          5284 => x"fe",
          5285 => x"83",
          5286 => x"fe",
          5287 => x"0b",
          5288 => x"0c",
          5289 => x"bb",
          5290 => x"3d",
          5291 => x"fa",
          5292 => x"59",
          5293 => x"19",
          5294 => x"83",
          5295 => x"70",
          5296 => x"58",
          5297 => x"f9",
          5298 => x"0b",
          5299 => x"34",
          5300 => x"bb",
          5301 => x"3d",
          5302 => x"fa",
          5303 => x"5b",
          5304 => x"1b",
          5305 => x"83",
          5306 => x"84",
          5307 => x"83",
          5308 => x"5b",
          5309 => x"5c",
          5310 => x"84",
          5311 => x"9c",
          5312 => x"53",
          5313 => x"ff",
          5314 => x"84",
          5315 => x"80",
          5316 => x"38",
          5317 => x"33",
          5318 => x"5a",
          5319 => x"85",
          5320 => x"83",
          5321 => x"02",
          5322 => x"22",
          5323 => x"d8",
          5324 => x"cf",
          5325 => x"b6",
          5326 => x"84",
          5327 => x"33",
          5328 => x"fa",
          5329 => x"b8",
          5330 => x"fa",
          5331 => x"5b",
          5332 => x"39",
          5333 => x"33",
          5334 => x"33",
          5335 => x"33",
          5336 => x"05",
          5337 => x"84",
          5338 => x"33",
          5339 => x"a0",
          5340 => x"84",
          5341 => x"83",
          5342 => x"83",
          5343 => x"72",
          5344 => x"5a",
          5345 => x"78",
          5346 => x"18",
          5347 => x"b4",
          5348 => x"29",
          5349 => x"83",
          5350 => x"60",
          5351 => x"80",
          5352 => x"b8",
          5353 => x"81",
          5354 => x"fa",
          5355 => x"fa",
          5356 => x"72",
          5357 => x"5f",
          5358 => x"83",
          5359 => x"84",
          5360 => x"34",
          5361 => x"81",
          5362 => x"58",
          5363 => x"90",
          5364 => x"b8",
          5365 => x"77",
          5366 => x"ff",
          5367 => x"83",
          5368 => x"80",
          5369 => x"80",
          5370 => x"fb",
          5371 => x"80",
          5372 => x"38",
          5373 => x"33",
          5374 => x"b4",
          5375 => x"81",
          5376 => x"3f",
          5377 => x"bb",
          5378 => x"3d",
          5379 => x"ba",
          5380 => x"fa",
          5381 => x"ba",
          5382 => x"fa",
          5383 => x"ba",
          5384 => x"76",
          5385 => x"23",
          5386 => x"83",
          5387 => x"84",
          5388 => x"83",
          5389 => x"84",
          5390 => x"83",
          5391 => x"84",
          5392 => x"ff",
          5393 => x"ba",
          5394 => x"7a",
          5395 => x"93",
          5396 => x"d8",
          5397 => x"86",
          5398 => x"06",
          5399 => x"83",
          5400 => x"81",
          5401 => x"fa",
          5402 => x"05",
          5403 => x"83",
          5404 => x"94",
          5405 => x"57",
          5406 => x"3f",
          5407 => x"fd",
          5408 => x"bb",
          5409 => x"ff",
          5410 => x"88",
          5411 => x"05",
          5412 => x"24",
          5413 => x"76",
          5414 => x"e8",
          5415 => x"f5",
          5416 => x"39",
          5417 => x"ba",
          5418 => x"58",
          5419 => x"06",
          5420 => x"27",
          5421 => x"77",
          5422 => x"d8",
          5423 => x"33",
          5424 => x"b1",
          5425 => x"38",
          5426 => x"83",
          5427 => x"5f",
          5428 => x"84",
          5429 => x"5e",
          5430 => x"8f",
          5431 => x"fa",
          5432 => x"ba",
          5433 => x"71",
          5434 => x"70",
          5435 => x"06",
          5436 => x"5e",
          5437 => x"fa",
          5438 => x"e7",
          5439 => x"85",
          5440 => x"80",
          5441 => x"38",
          5442 => x"33",
          5443 => x"81",
          5444 => x"b8",
          5445 => x"57",
          5446 => x"27",
          5447 => x"75",
          5448 => x"34",
          5449 => x"80",
          5450 => x"b5",
          5451 => x"b4",
          5452 => x"ff",
          5453 => x"7b",
          5454 => x"a7",
          5455 => x"56",
          5456 => x"b4",
          5457 => x"39",
          5458 => x"fa",
          5459 => x"fa",
          5460 => x"b8",
          5461 => x"05",
          5462 => x"76",
          5463 => x"38",
          5464 => x"75",
          5465 => x"34",
          5466 => x"84",
          5467 => x"40",
          5468 => x"8d",
          5469 => x"fa",
          5470 => x"ba",
          5471 => x"71",
          5472 => x"70",
          5473 => x"06",
          5474 => x"42",
          5475 => x"fa",
          5476 => x"cf",
          5477 => x"85",
          5478 => x"80",
          5479 => x"38",
          5480 => x"22",
          5481 => x"2e",
          5482 => x"fc",
          5483 => x"b8",
          5484 => x"fa",
          5485 => x"fa",
          5486 => x"71",
          5487 => x"c7",
          5488 => x"83",
          5489 => x"43",
          5490 => x"71",
          5491 => x"70",
          5492 => x"06",
          5493 => x"08",
          5494 => x"80",
          5495 => x"5d",
          5496 => x"82",
          5497 => x"bf",
          5498 => x"83",
          5499 => x"fb",
          5500 => x"ba",
          5501 => x"79",
          5502 => x"e7",
          5503 => x"d8",
          5504 => x"99",
          5505 => x"06",
          5506 => x"81",
          5507 => x"89",
          5508 => x"39",
          5509 => x"33",
          5510 => x"2e",
          5511 => x"84",
          5512 => x"83",
          5513 => x"5d",
          5514 => x"b8",
          5515 => x"11",
          5516 => x"75",
          5517 => x"38",
          5518 => x"83",
          5519 => x"fb",
          5520 => x"ba",
          5521 => x"76",
          5522 => x"c8",
          5523 => x"d9",
          5524 => x"b4",
          5525 => x"05",
          5526 => x"33",
          5527 => x"41",
          5528 => x"25",
          5529 => x"57",
          5530 => x"b4",
          5531 => x"39",
          5532 => x"51",
          5533 => x"3f",
          5534 => x"ba",
          5535 => x"57",
          5536 => x"8b",
          5537 => x"10",
          5538 => x"05",
          5539 => x"5a",
          5540 => x"51",
          5541 => x"3f",
          5542 => x"81",
          5543 => x"ba",
          5544 => x"58",
          5545 => x"82",
          5546 => x"85",
          5547 => x"7d",
          5548 => x"38",
          5549 => x"22",
          5550 => x"26",
          5551 => x"57",
          5552 => x"81",
          5553 => x"d5",
          5554 => x"97",
          5555 => x"85",
          5556 => x"77",
          5557 => x"38",
          5558 => x"33",
          5559 => x"81",
          5560 => x"ba",
          5561 => x"05",
          5562 => x"06",
          5563 => x"33",
          5564 => x"06",
          5565 => x"43",
          5566 => x"5c",
          5567 => x"27",
          5568 => x"5a",
          5569 => x"b2",
          5570 => x"ff",
          5571 => x"58",
          5572 => x"27",
          5573 => x"57",
          5574 => x"b4",
          5575 => x"f8",
          5576 => x"57",
          5577 => x"27",
          5578 => x"7a",
          5579 => x"fa",
          5580 => x"af",
          5581 => x"85",
          5582 => x"80",
          5583 => x"38",
          5584 => x"33",
          5585 => x"33",
          5586 => x"7f",
          5587 => x"38",
          5588 => x"33",
          5589 => x"33",
          5590 => x"06",
          5591 => x"33",
          5592 => x"11",
          5593 => x"80",
          5594 => x"b2",
          5595 => x"71",
          5596 => x"70",
          5597 => x"06",
          5598 => x"33",
          5599 => x"59",
          5600 => x"81",
          5601 => x"38",
          5602 => x"ff",
          5603 => x"31",
          5604 => x"7c",
          5605 => x"38",
          5606 => x"33",
          5607 => x"27",
          5608 => x"ff",
          5609 => x"83",
          5610 => x"7c",
          5611 => x"70",
          5612 => x"57",
          5613 => x"8e",
          5614 => x"b8",
          5615 => x"76",
          5616 => x"ee",
          5617 => x"56",
          5618 => x"b4",
          5619 => x"ff",
          5620 => x"b2",
          5621 => x"80",
          5622 => x"26",
          5623 => x"77",
          5624 => x"7e",
          5625 => x"71",
          5626 => x"5e",
          5627 => x"86",
          5628 => x"5b",
          5629 => x"80",
          5630 => x"06",
          5631 => x"06",
          5632 => x"1d",
          5633 => x"5c",
          5634 => x"f7",
          5635 => x"99",
          5636 => x"e0",
          5637 => x"5f",
          5638 => x"1f",
          5639 => x"81",
          5640 => x"76",
          5641 => x"58",
          5642 => x"81",
          5643 => x"81",
          5644 => x"f8",
          5645 => x"f7",
          5646 => x"29",
          5647 => x"5e",
          5648 => x"27",
          5649 => x"e0",
          5650 => x"5f",
          5651 => x"1f",
          5652 => x"81",
          5653 => x"76",
          5654 => x"58",
          5655 => x"81",
          5656 => x"81",
          5657 => x"f8",
          5658 => x"f7",
          5659 => x"29",
          5660 => x"5e",
          5661 => x"26",
          5662 => x"f6",
          5663 => x"ba",
          5664 => x"75",
          5665 => x"e0",
          5666 => x"84",
          5667 => x"51",
          5668 => x"f6",
          5669 => x"0b",
          5670 => x"33",
          5671 => x"ba",
          5672 => x"59",
          5673 => x"78",
          5674 => x"84",
          5675 => x"56",
          5676 => x"09",
          5677 => x"be",
          5678 => x"b5",
          5679 => x"81",
          5680 => x"fa",
          5681 => x"43",
          5682 => x"ff",
          5683 => x"38",
          5684 => x"33",
          5685 => x"26",
          5686 => x"7e",
          5687 => x"56",
          5688 => x"f5",
          5689 => x"76",
          5690 => x"27",
          5691 => x"f5",
          5692 => x"10",
          5693 => x"90",
          5694 => x"86",
          5695 => x"11",
          5696 => x"5a",
          5697 => x"80",
          5698 => x"06",
          5699 => x"75",
          5700 => x"79",
          5701 => x"76",
          5702 => x"83",
          5703 => x"70",
          5704 => x"90",
          5705 => x"88",
          5706 => x"07",
          5707 => x"52",
          5708 => x"7a",
          5709 => x"80",
          5710 => x"05",
          5711 => x"76",
          5712 => x"58",
          5713 => x"26",
          5714 => x"b8",
          5715 => x"b8",
          5716 => x"5f",
          5717 => x"06",
          5718 => x"06",
          5719 => x"22",
          5720 => x"64",
          5721 => x"59",
          5722 => x"26",
          5723 => x"78",
          5724 => x"7b",
          5725 => x"57",
          5726 => x"1d",
          5727 => x"76",
          5728 => x"38",
          5729 => x"33",
          5730 => x"18",
          5731 => x"0b",
          5732 => x"34",
          5733 => x"81",
          5734 => x"81",
          5735 => x"76",
          5736 => x"38",
          5737 => x"e0",
          5738 => x"78",
          5739 => x"5a",
          5740 => x"57",
          5741 => x"d6",
          5742 => x"39",
          5743 => x"81",
          5744 => x"58",
          5745 => x"83",
          5746 => x"70",
          5747 => x"71",
          5748 => x"f0",
          5749 => x"2a",
          5750 => x"57",
          5751 => x"2e",
          5752 => x"be",
          5753 => x"0b",
          5754 => x"34",
          5755 => x"81",
          5756 => x"56",
          5757 => x"83",
          5758 => x"33",
          5759 => x"80",
          5760 => x"34",
          5761 => x"33",
          5762 => x"33",
          5763 => x"22",
          5764 => x"33",
          5765 => x"5d",
          5766 => x"83",
          5767 => x"87",
          5768 => x"83",
          5769 => x"81",
          5770 => x"ff",
          5771 => x"f4",
          5772 => x"fa",
          5773 => x"fd",
          5774 => x"56",
          5775 => x"b0",
          5776 => x"83",
          5777 => x"81",
          5778 => x"07",
          5779 => x"fa",
          5780 => x"39",
          5781 => x"33",
          5782 => x"81",
          5783 => x"83",
          5784 => x"c3",
          5785 => x"b0",
          5786 => x"06",
          5787 => x"75",
          5788 => x"34",
          5789 => x"80",
          5790 => x"fa",
          5791 => x"18",
          5792 => x"06",
          5793 => x"a4",
          5794 => x"b0",
          5795 => x"06",
          5796 => x"fa",
          5797 => x"8f",
          5798 => x"b0",
          5799 => x"06",
          5800 => x"75",
          5801 => x"34",
          5802 => x"83",
          5803 => x"81",
          5804 => x"e0",
          5805 => x"83",
          5806 => x"fe",
          5807 => x"fa",
          5808 => x"cf",
          5809 => x"07",
          5810 => x"fa",
          5811 => x"d7",
          5812 => x"b0",
          5813 => x"06",
          5814 => x"75",
          5815 => x"34",
          5816 => x"83",
          5817 => x"81",
          5818 => x"07",
          5819 => x"fa",
          5820 => x"b3",
          5821 => x"b0",
          5822 => x"06",
          5823 => x"75",
          5824 => x"34",
          5825 => x"83",
          5826 => x"81",
          5827 => x"07",
          5828 => x"fa",
          5829 => x"8f",
          5830 => x"b0",
          5831 => x"06",
          5832 => x"fa",
          5833 => x"ff",
          5834 => x"b0",
          5835 => x"07",
          5836 => x"fa",
          5837 => x"ef",
          5838 => x"b0",
          5839 => x"07",
          5840 => x"fa",
          5841 => x"df",
          5842 => x"b0",
          5843 => x"06",
          5844 => x"56",
          5845 => x"b0",
          5846 => x"39",
          5847 => x"33",
          5848 => x"b0",
          5849 => x"83",
          5850 => x"fd",
          5851 => x"0b",
          5852 => x"34",
          5853 => x"51",
          5854 => x"ec",
          5855 => x"ba",
          5856 => x"fa",
          5857 => x"ba",
          5858 => x"fa",
          5859 => x"ba",
          5860 => x"78",
          5861 => x"23",
          5862 => x"ba",
          5863 => x"c7",
          5864 => x"84",
          5865 => x"80",
          5866 => x"84",
          5867 => x"0d",
          5868 => x"fa",
          5869 => x"fa",
          5870 => x"81",
          5871 => x"ff",
          5872 => x"cf",
          5873 => x"88",
          5874 => x"dc",
          5875 => x"05",
          5876 => x"b5",
          5877 => x"84",
          5878 => x"84",
          5879 => x"84",
          5880 => x"80",
          5881 => x"84",
          5882 => x"84",
          5883 => x"9c",
          5884 => x"77",
          5885 => x"34",
          5886 => x"84",
          5887 => x"81",
          5888 => x"7a",
          5889 => x"34",
          5890 => x"fe",
          5891 => x"80",
          5892 => x"84",
          5893 => x"23",
          5894 => x"ba",
          5895 => x"39",
          5896 => x"fa",
          5897 => x"52",
          5898 => x"97",
          5899 => x"b5",
          5900 => x"ff",
          5901 => x"05",
          5902 => x"39",
          5903 => x"fa",
          5904 => x"52",
          5905 => x"fb",
          5906 => x"39",
          5907 => x"ea",
          5908 => x"8f",
          5909 => x"b5",
          5910 => x"70",
          5911 => x"2c",
          5912 => x"5f",
          5913 => x"39",
          5914 => x"51",
          5915 => x"b8",
          5916 => x"75",
          5917 => x"eb",
          5918 => x"fa",
          5919 => x"e3",
          5920 => x"b4",
          5921 => x"70",
          5922 => x"2c",
          5923 => x"40",
          5924 => x"39",
          5925 => x"33",
          5926 => x"b8",
          5927 => x"11",
          5928 => x"75",
          5929 => x"c0",
          5930 => x"f3",
          5931 => x"b8",
          5932 => x"81",
          5933 => x"5c",
          5934 => x"ee",
          5935 => x"fa",
          5936 => x"b8",
          5937 => x"81",
          5938 => x"fa",
          5939 => x"74",
          5940 => x"c7",
          5941 => x"83",
          5942 => x"5f",
          5943 => x"29",
          5944 => x"ff",
          5945 => x"f9",
          5946 => x"5b",
          5947 => x"5d",
          5948 => x"81",
          5949 => x"83",
          5950 => x"ff",
          5951 => x"80",
          5952 => x"89",
          5953 => x"f7",
          5954 => x"76",
          5955 => x"38",
          5956 => x"75",
          5957 => x"23",
          5958 => x"06",
          5959 => x"57",
          5960 => x"83",
          5961 => x"b8",
          5962 => x"76",
          5963 => x"ec",
          5964 => x"56",
          5965 => x"b4",
          5966 => x"ff",
          5967 => x"b2",
          5968 => x"80",
          5969 => x"26",
          5970 => x"77",
          5971 => x"7e",
          5972 => x"71",
          5973 => x"5e",
          5974 => x"86",
          5975 => x"5b",
          5976 => x"80",
          5977 => x"06",
          5978 => x"06",
          5979 => x"1d",
          5980 => x"5d",
          5981 => x"ec",
          5982 => x"99",
          5983 => x"e0",
          5984 => x"5e",
          5985 => x"1e",
          5986 => x"81",
          5987 => x"76",
          5988 => x"58",
          5989 => x"81",
          5990 => x"81",
          5991 => x"f8",
          5992 => x"f7",
          5993 => x"29",
          5994 => x"5d",
          5995 => x"27",
          5996 => x"e0",
          5997 => x"5e",
          5998 => x"1e",
          5999 => x"81",
          6000 => x"76",
          6001 => x"58",
          6002 => x"81",
          6003 => x"81",
          6004 => x"f8",
          6005 => x"f7",
          6006 => x"29",
          6007 => x"5d",
          6008 => x"26",
          6009 => x"eb",
          6010 => x"fa",
          6011 => x"5c",
          6012 => x"1c",
          6013 => x"83",
          6014 => x"84",
          6015 => x"83",
          6016 => x"84",
          6017 => x"5f",
          6018 => x"fd",
          6019 => x"eb",
          6020 => x"b8",
          6021 => x"81",
          6022 => x"11",
          6023 => x"76",
          6024 => x"38",
          6025 => x"83",
          6026 => x"77",
          6027 => x"ff",
          6028 => x"80",
          6029 => x"38",
          6030 => x"83",
          6031 => x"84",
          6032 => x"70",
          6033 => x"ff",
          6034 => x"56",
          6035 => x"eb",
          6036 => x"56",
          6037 => x"b5",
          6038 => x"39",
          6039 => x"33",
          6040 => x"b8",
          6041 => x"11",
          6042 => x"75",
          6043 => x"ca",
          6044 => x"ef",
          6045 => x"81",
          6046 => x"06",
          6047 => x"83",
          6048 => x"70",
          6049 => x"83",
          6050 => x"7a",
          6051 => x"57",
          6052 => x"09",
          6053 => x"b8",
          6054 => x"39",
          6055 => x"75",
          6056 => x"34",
          6057 => x"ff",
          6058 => x"83",
          6059 => x"fc",
          6060 => x"7b",
          6061 => x"83",
          6062 => x"f2",
          6063 => x"7d",
          6064 => x"7a",
          6065 => x"38",
          6066 => x"81",
          6067 => x"83",
          6068 => x"77",
          6069 => x"59",
          6070 => x"26",
          6071 => x"80",
          6072 => x"05",
          6073 => x"fa",
          6074 => x"70",
          6075 => x"34",
          6076 => x"d4",
          6077 => x"39",
          6078 => x"56",
          6079 => x"b2",
          6080 => x"39",
          6081 => x"fa",
          6082 => x"ad",
          6083 => x"fa",
          6084 => x"84",
          6085 => x"83",
          6086 => x"f1",
          6087 => x"0b",
          6088 => x"34",
          6089 => x"83",
          6090 => x"33",
          6091 => x"80",
          6092 => x"34",
          6093 => x"f9",
          6094 => x"a7",
          6095 => x"0d",
          6096 => x"33",
          6097 => x"33",
          6098 => x"80",
          6099 => x"73",
          6100 => x"3f",
          6101 => x"bb",
          6102 => x"3d",
          6103 => x"52",
          6104 => x"ab",
          6105 => x"84",
          6106 => x"85",
          6107 => x"f3",
          6108 => x"bf",
          6109 => x"ff",
          6110 => x"88",
          6111 => x"ff",
          6112 => x"e8",
          6113 => x"55",
          6114 => x"80",
          6115 => x"38",
          6116 => x"75",
          6117 => x"34",
          6118 => x"84",
          6119 => x"8f",
          6120 => x"83",
          6121 => x"54",
          6122 => x"80",
          6123 => x"73",
          6124 => x"30",
          6125 => x"09",
          6126 => x"56",
          6127 => x"72",
          6128 => x"0c",
          6129 => x"54",
          6130 => x"09",
          6131 => x"38",
          6132 => x"83",
          6133 => x"70",
          6134 => x"07",
          6135 => x"79",
          6136 => x"c4",
          6137 => x"f8",
          6138 => x"b5",
          6139 => x"b4",
          6140 => x"29",
          6141 => x"a0",
          6142 => x"fa",
          6143 => x"59",
          6144 => x"29",
          6145 => x"ff",
          6146 => x"f9",
          6147 => x"59",
          6148 => x"81",
          6149 => x"38",
          6150 => x"73",
          6151 => x"80",
          6152 => x"87",
          6153 => x"0c",
          6154 => x"88",
          6155 => x"80",
          6156 => x"87",
          6157 => x"08",
          6158 => x"f6",
          6159 => x"81",
          6160 => x"ff",
          6161 => x"81",
          6162 => x"cf",
          6163 => x"83",
          6164 => x"33",
          6165 => x"06",
          6166 => x"16",
          6167 => x"55",
          6168 => x"85",
          6169 => x"81",
          6170 => x"b4",
          6171 => x"f8",
          6172 => x"75",
          6173 => x"5a",
          6174 => x"2e",
          6175 => x"75",
          6176 => x"15",
          6177 => x"a4",
          6178 => x"f8",
          6179 => x"81",
          6180 => x"ff",
          6181 => x"89",
          6182 => x"b3",
          6183 => x"ac",
          6184 => x"2b",
          6185 => x"58",
          6186 => x"83",
          6187 => x"73",
          6188 => x"70",
          6189 => x"32",
          6190 => x"51",
          6191 => x"80",
          6192 => x"38",
          6193 => x"f8",
          6194 => x"09",
          6195 => x"72",
          6196 => x"e4",
          6197 => x"83",
          6198 => x"80",
          6199 => x"dd",
          6200 => x"e4",
          6201 => x"de",
          6202 => x"f8",
          6203 => x"f8",
          6204 => x"5d",
          6205 => x"5e",
          6206 => x"b8",
          6207 => x"74",
          6208 => x"8d",
          6209 => x"cc",
          6210 => x"73",
          6211 => x"82",
          6212 => x"c2",
          6213 => x"72",
          6214 => x"8b",
          6215 => x"cc",
          6216 => x"73",
          6217 => x"74",
          6218 => x"54",
          6219 => x"2e",
          6220 => x"f8",
          6221 => x"53",
          6222 => x"81",
          6223 => x"81",
          6224 => x"72",
          6225 => x"84",
          6226 => x"f8",
          6227 => x"54",
          6228 => x"84",
          6229 => x"f8",
          6230 => x"e8",
          6231 => x"98",
          6232 => x"54",
          6233 => x"83",
          6234 => x"0b",
          6235 => x"9c",
          6236 => x"d8",
          6237 => x"16",
          6238 => x"06",
          6239 => x"76",
          6240 => x"38",
          6241 => x"df",
          6242 => x"f8",
          6243 => x"9e",
          6244 => x"9c",
          6245 => x"38",
          6246 => x"83",
          6247 => x"5a",
          6248 => x"83",
          6249 => x"54",
          6250 => x"91",
          6251 => x"14",
          6252 => x"9c",
          6253 => x"7d",
          6254 => x"dc",
          6255 => x"83",
          6256 => x"54",
          6257 => x"2e",
          6258 => x"54",
          6259 => x"8a",
          6260 => x"98",
          6261 => x"f9",
          6262 => x"81",
          6263 => x"77",
          6264 => x"38",
          6265 => x"17",
          6266 => x"b9",
          6267 => x"76",
          6268 => x"54",
          6269 => x"83",
          6270 => x"53",
          6271 => x"82",
          6272 => x"81",
          6273 => x"38",
          6274 => x"34",
          6275 => x"fc",
          6276 => x"58",
          6277 => x"80",
          6278 => x"83",
          6279 => x"2e",
          6280 => x"77",
          6281 => x"06",
          6282 => x"7d",
          6283 => x"ed",
          6284 => x"2e",
          6285 => x"79",
          6286 => x"59",
          6287 => x"75",
          6288 => x"54",
          6289 => x"a1",
          6290 => x"2e",
          6291 => x"17",
          6292 => x"06",
          6293 => x"fe",
          6294 => x"27",
          6295 => x"57",
          6296 => x"54",
          6297 => x"e1",
          6298 => x"10",
          6299 => x"05",
          6300 => x"2b",
          6301 => x"f5",
          6302 => x"33",
          6303 => x"78",
          6304 => x"9c",
          6305 => x"d8",
          6306 => x"ea",
          6307 => x"7d",
          6308 => x"a8",
          6309 => x"ff",
          6310 => x"a0",
          6311 => x"ff",
          6312 => x"ff",
          6313 => x"38",
          6314 => x"b8",
          6315 => x"54",
          6316 => x"83",
          6317 => x"82",
          6318 => x"70",
          6319 => x"07",
          6320 => x"7d",
          6321 => x"83",
          6322 => x"06",
          6323 => x"78",
          6324 => x"c6",
          6325 => x"72",
          6326 => x"83",
          6327 => x"70",
          6328 => x"78",
          6329 => x"ba",
          6330 => x"70",
          6331 => x"54",
          6332 => x"27",
          6333 => x"b8",
          6334 => x"72",
          6335 => x"9a",
          6336 => x"fc",
          6337 => x"f9",
          6338 => x"81",
          6339 => x"82",
          6340 => x"3f",
          6341 => x"84",
          6342 => x"0d",
          6343 => x"34",
          6344 => x"f9",
          6345 => x"81",
          6346 => x"38",
          6347 => x"14",
          6348 => x"5b",
          6349 => x"cc",
          6350 => x"c9",
          6351 => x"83",
          6352 => x"34",
          6353 => x"f8",
          6354 => x"ff",
          6355 => x"c2",
          6356 => x"b1",
          6357 => x"ff",
          6358 => x"81",
          6359 => x"96",
          6360 => x"cc",
          6361 => x"81",
          6362 => x"8a",
          6363 => x"ff",
          6364 => x"81",
          6365 => x"06",
          6366 => x"83",
          6367 => x"81",
          6368 => x"c0",
          6369 => x"54",
          6370 => x"27",
          6371 => x"87",
          6372 => x"08",
          6373 => x"0c",
          6374 => x"06",
          6375 => x"39",
          6376 => x"f8",
          6377 => x"f9",
          6378 => x"83",
          6379 => x"73",
          6380 => x"53",
          6381 => x"38",
          6382 => x"de",
          6383 => x"83",
          6384 => x"83",
          6385 => x"83",
          6386 => x"70",
          6387 => x"33",
          6388 => x"33",
          6389 => x"5e",
          6390 => x"fa",
          6391 => x"82",
          6392 => x"06",
          6393 => x"7a",
          6394 => x"2e",
          6395 => x"79",
          6396 => x"81",
          6397 => x"38",
          6398 => x"ef",
          6399 => x"f0",
          6400 => x"39",
          6401 => x"b8",
          6402 => x"54",
          6403 => x"81",
          6404 => x"b8",
          6405 => x"59",
          6406 => x"80",
          6407 => x"fa",
          6408 => x"76",
          6409 => x"54",
          6410 => x"fa",
          6411 => x"f7",
          6412 => x"53",
          6413 => x"08",
          6414 => x"83",
          6415 => x"83",
          6416 => x"f6",
          6417 => x"b8",
          6418 => x"81",
          6419 => x"11",
          6420 => x"80",
          6421 => x"38",
          6422 => x"83",
          6423 => x"73",
          6424 => x"ff",
          6425 => x"80",
          6426 => x"38",
          6427 => x"83",
          6428 => x"84",
          6429 => x"70",
          6430 => x"56",
          6431 => x"80",
          6432 => x"38",
          6433 => x"83",
          6434 => x"ff",
          6435 => x"39",
          6436 => x"51",
          6437 => x"3f",
          6438 => x"aa",
          6439 => x"fc",
          6440 => x"14",
          6441 => x"f8",
          6442 => x"dd",
          6443 => x"0b",
          6444 => x"34",
          6445 => x"33",
          6446 => x"39",
          6447 => x"81",
          6448 => x"3f",
          6449 => x"04",
          6450 => x"80",
          6451 => x"90",
          6452 => x"02",
          6453 => x"82",
          6454 => x"f5",
          6455 => x"80",
          6456 => x"85",
          6457 => x"90",
          6458 => x"fe",
          6459 => x"34",
          6460 => x"90",
          6461 => x"87",
          6462 => x"08",
          6463 => x"08",
          6464 => x"90",
          6465 => x"c0",
          6466 => x"52",
          6467 => x"9c",
          6468 => x"72",
          6469 => x"81",
          6470 => x"c0",
          6471 => x"56",
          6472 => x"27",
          6473 => x"81",
          6474 => x"38",
          6475 => x"a4",
          6476 => x"55",
          6477 => x"80",
          6478 => x"55",
          6479 => x"80",
          6480 => x"c0",
          6481 => x"80",
          6482 => x"53",
          6483 => x"9c",
          6484 => x"c0",
          6485 => x"55",
          6486 => x"f6",
          6487 => x"33",
          6488 => x"9c",
          6489 => x"70",
          6490 => x"38",
          6491 => x"2e",
          6492 => x"c0",
          6493 => x"55",
          6494 => x"83",
          6495 => x"71",
          6496 => x"70",
          6497 => x"57",
          6498 => x"2e",
          6499 => x"81",
          6500 => x"71",
          6501 => x"74",
          6502 => x"38",
          6503 => x"84",
          6504 => x"0d",
          6505 => x"84",
          6506 => x"88",
          6507 => x"fa",
          6508 => x"02",
          6509 => x"05",
          6510 => x"80",
          6511 => x"90",
          6512 => x"2b",
          6513 => x"80",
          6514 => x"98",
          6515 => x"55",
          6516 => x"83",
          6517 => x"90",
          6518 => x"84",
          6519 => x"90",
          6520 => x"85",
          6521 => x"86",
          6522 => x"f5",
          6523 => x"74",
          6524 => x"83",
          6525 => x"51",
          6526 => x"34",
          6527 => x"f5",
          6528 => x"56",
          6529 => x"15",
          6530 => x"87",
          6531 => x"34",
          6532 => x"9c",
          6533 => x"90",
          6534 => x"ce",
          6535 => x"87",
          6536 => x"08",
          6537 => x"98",
          6538 => x"70",
          6539 => x"38",
          6540 => x"87",
          6541 => x"08",
          6542 => x"73",
          6543 => x"71",
          6544 => x"db",
          6545 => x"98",
          6546 => x"ff",
          6547 => x"27",
          6548 => x"71",
          6549 => x"2e",
          6550 => x"87",
          6551 => x"08",
          6552 => x"05",
          6553 => x"98",
          6554 => x"87",
          6555 => x"08",
          6556 => x"2e",
          6557 => x"14",
          6558 => x"98",
          6559 => x"52",
          6560 => x"87",
          6561 => x"ff",
          6562 => x"87",
          6563 => x"08",
          6564 => x"26",
          6565 => x"52",
          6566 => x"16",
          6567 => x"06",
          6568 => x"80",
          6569 => x"38",
          6570 => x"06",
          6571 => x"d4",
          6572 => x"70",
          6573 => x"56",
          6574 => x"80",
          6575 => x"84",
          6576 => x"52",
          6577 => x"27",
          6578 => x"70",
          6579 => x"33",
          6580 => x"05",
          6581 => x"71",
          6582 => x"76",
          6583 => x"0c",
          6584 => x"04",
          6585 => x"bb",
          6586 => x"3d",
          6587 => x"51",
          6588 => x"3d",
          6589 => x"84",
          6590 => x"33",
          6591 => x"0b",
          6592 => x"08",
          6593 => x"87",
          6594 => x"06",
          6595 => x"2a",
          6596 => x"55",
          6597 => x"15",
          6598 => x"2a",
          6599 => x"15",
          6600 => x"2a",
          6601 => x"15",
          6602 => x"15",
          6603 => x"f5",
          6604 => x"c6",
          6605 => x"13",
          6606 => x"51",
          6607 => x"97",
          6608 => x"81",
          6609 => x"72",
          6610 => x"54",
          6611 => x"26",
          6612 => x"f5",
          6613 => x"74",
          6614 => x"83",
          6615 => x"55",
          6616 => x"34",
          6617 => x"f5",
          6618 => x"56",
          6619 => x"15",
          6620 => x"87",
          6621 => x"34",
          6622 => x"9c",
          6623 => x"90",
          6624 => x"ce",
          6625 => x"87",
          6626 => x"08",
          6627 => x"98",
          6628 => x"70",
          6629 => x"38",
          6630 => x"87",
          6631 => x"08",
          6632 => x"73",
          6633 => x"71",
          6634 => x"db",
          6635 => x"98",
          6636 => x"ff",
          6637 => x"27",
          6638 => x"71",
          6639 => x"2e",
          6640 => x"87",
          6641 => x"08",
          6642 => x"05",
          6643 => x"98",
          6644 => x"87",
          6645 => x"08",
          6646 => x"2e",
          6647 => x"14",
          6648 => x"98",
          6649 => x"52",
          6650 => x"87",
          6651 => x"ff",
          6652 => x"87",
          6653 => x"08",
          6654 => x"26",
          6655 => x"52",
          6656 => x"16",
          6657 => x"06",
          6658 => x"80",
          6659 => x"74",
          6660 => x"52",
          6661 => x"38",
          6662 => x"81",
          6663 => x"73",
          6664 => x"38",
          6665 => x"84",
          6666 => x"88",
          6667 => x"ff",
          6668 => x"fb",
          6669 => x"f5",
          6670 => x"80",
          6671 => x"85",
          6672 => x"90",
          6673 => x"fe",
          6674 => x"34",
          6675 => x"90",
          6676 => x"87",
          6677 => x"08",
          6678 => x"08",
          6679 => x"90",
          6680 => x"c0",
          6681 => x"52",
          6682 => x"9c",
          6683 => x"72",
          6684 => x"81",
          6685 => x"c0",
          6686 => x"52",
          6687 => x"27",
          6688 => x"81",
          6689 => x"38",
          6690 => x"a4",
          6691 => x"53",
          6692 => x"80",
          6693 => x"53",
          6694 => x"80",
          6695 => x"c0",
          6696 => x"80",
          6697 => x"53",
          6698 => x"9c",
          6699 => x"c0",
          6700 => x"51",
          6701 => x"f6",
          6702 => x"33",
          6703 => x"9c",
          6704 => x"73",
          6705 => x"38",
          6706 => x"2e",
          6707 => x"c0",
          6708 => x"51",
          6709 => x"83",
          6710 => x"71",
          6711 => x"70",
          6712 => x"57",
          6713 => x"2e",
          6714 => x"81",
          6715 => x"73",
          6716 => x"ff",
          6717 => x"0d",
          6718 => x"51",
          6719 => x"3f",
          6720 => x"04",
          6721 => x"84",
          6722 => x"7a",
          6723 => x"2a",
          6724 => x"ff",
          6725 => x"2b",
          6726 => x"33",
          6727 => x"71",
          6728 => x"83",
          6729 => x"11",
          6730 => x"12",
          6731 => x"2b",
          6732 => x"07",
          6733 => x"53",
          6734 => x"59",
          6735 => x"53",
          6736 => x"81",
          6737 => x"16",
          6738 => x"83",
          6739 => x"8b",
          6740 => x"2b",
          6741 => x"70",
          6742 => x"33",
          6743 => x"71",
          6744 => x"57",
          6745 => x"59",
          6746 => x"71",
          6747 => x"38",
          6748 => x"85",
          6749 => x"8b",
          6750 => x"2b",
          6751 => x"76",
          6752 => x"54",
          6753 => x"86",
          6754 => x"81",
          6755 => x"73",
          6756 => x"84",
          6757 => x"70",
          6758 => x"33",
          6759 => x"71",
          6760 => x"70",
          6761 => x"55",
          6762 => x"77",
          6763 => x"71",
          6764 => x"84",
          6765 => x"16",
          6766 => x"86",
          6767 => x"0b",
          6768 => x"84",
          6769 => x"53",
          6770 => x"34",
          6771 => x"34",
          6772 => x"08",
          6773 => x"81",
          6774 => x"88",
          6775 => x"80",
          6776 => x"88",
          6777 => x"52",
          6778 => x"34",
          6779 => x"34",
          6780 => x"04",
          6781 => x"87",
          6782 => x"8b",
          6783 => x"2b",
          6784 => x"84",
          6785 => x"17",
          6786 => x"2b",
          6787 => x"2a",
          6788 => x"51",
          6789 => x"71",
          6790 => x"72",
          6791 => x"84",
          6792 => x"70",
          6793 => x"33",
          6794 => x"71",
          6795 => x"83",
          6796 => x"5a",
          6797 => x"05",
          6798 => x"87",
          6799 => x"88",
          6800 => x"88",
          6801 => x"59",
          6802 => x"13",
          6803 => x"13",
          6804 => x"f4",
          6805 => x"33",
          6806 => x"71",
          6807 => x"81",
          6808 => x"70",
          6809 => x"5a",
          6810 => x"72",
          6811 => x"13",
          6812 => x"f4",
          6813 => x"70",
          6814 => x"33",
          6815 => x"71",
          6816 => x"74",
          6817 => x"81",
          6818 => x"88",
          6819 => x"83",
          6820 => x"f8",
          6821 => x"7b",
          6822 => x"52",
          6823 => x"5a",
          6824 => x"77",
          6825 => x"73",
          6826 => x"84",
          6827 => x"70",
          6828 => x"81",
          6829 => x"8b",
          6830 => x"2b",
          6831 => x"70",
          6832 => x"33",
          6833 => x"07",
          6834 => x"06",
          6835 => x"5f",
          6836 => x"5a",
          6837 => x"77",
          6838 => x"81",
          6839 => x"ba",
          6840 => x"17",
          6841 => x"83",
          6842 => x"8b",
          6843 => x"2b",
          6844 => x"70",
          6845 => x"33",
          6846 => x"71",
          6847 => x"58",
          6848 => x"5a",
          6849 => x"70",
          6850 => x"e4",
          6851 => x"81",
          6852 => x"88",
          6853 => x"80",
          6854 => x"88",
          6855 => x"54",
          6856 => x"77",
          6857 => x"84",
          6858 => x"70",
          6859 => x"81",
          6860 => x"8b",
          6861 => x"2b",
          6862 => x"82",
          6863 => x"15",
          6864 => x"2b",
          6865 => x"2a",
          6866 => x"52",
          6867 => x"53",
          6868 => x"34",
          6869 => x"34",
          6870 => x"04",
          6871 => x"79",
          6872 => x"08",
          6873 => x"80",
          6874 => x"77",
          6875 => x"38",
          6876 => x"90",
          6877 => x"0d",
          6878 => x"f4",
          6879 => x"f4",
          6880 => x"0b",
          6881 => x"23",
          6882 => x"53",
          6883 => x"ff",
          6884 => x"d1",
          6885 => x"ba",
          6886 => x"76",
          6887 => x"0b",
          6888 => x"84",
          6889 => x"54",
          6890 => x"34",
          6891 => x"15",
          6892 => x"f4",
          6893 => x"86",
          6894 => x"0b",
          6895 => x"84",
          6896 => x"84",
          6897 => x"ff",
          6898 => x"80",
          6899 => x"ff",
          6900 => x"88",
          6901 => x"55",
          6902 => x"17",
          6903 => x"17",
          6904 => x"f0",
          6905 => x"10",
          6906 => x"f4",
          6907 => x"05",
          6908 => x"82",
          6909 => x"0b",
          6910 => x"fe",
          6911 => x"3d",
          6912 => x"80",
          6913 => x"84",
          6914 => x"38",
          6915 => x"2a",
          6916 => x"83",
          6917 => x"51",
          6918 => x"ff",
          6919 => x"ba",
          6920 => x"11",
          6921 => x"33",
          6922 => x"07",
          6923 => x"5a",
          6924 => x"ff",
          6925 => x"80",
          6926 => x"38",
          6927 => x"10",
          6928 => x"81",
          6929 => x"88",
          6930 => x"81",
          6931 => x"79",
          6932 => x"ff",
          6933 => x"7a",
          6934 => x"5c",
          6935 => x"72",
          6936 => x"38",
          6937 => x"85",
          6938 => x"55",
          6939 => x"33",
          6940 => x"71",
          6941 => x"57",
          6942 => x"38",
          6943 => x"ff",
          6944 => x"77",
          6945 => x"80",
          6946 => x"78",
          6947 => x"81",
          6948 => x"88",
          6949 => x"81",
          6950 => x"56",
          6951 => x"59",
          6952 => x"2e",
          6953 => x"59",
          6954 => x"73",
          6955 => x"38",
          6956 => x"80",
          6957 => x"38",
          6958 => x"82",
          6959 => x"16",
          6960 => x"78",
          6961 => x"80",
          6962 => x"88",
          6963 => x"56",
          6964 => x"74",
          6965 => x"15",
          6966 => x"f4",
          6967 => x"88",
          6968 => x"71",
          6969 => x"75",
          6970 => x"84",
          6971 => x"70",
          6972 => x"81",
          6973 => x"88",
          6974 => x"83",
          6975 => x"f8",
          6976 => x"7e",
          6977 => x"06",
          6978 => x"5c",
          6979 => x"59",
          6980 => x"82",
          6981 => x"81",
          6982 => x"72",
          6983 => x"84",
          6984 => x"18",
          6985 => x"34",
          6986 => x"34",
          6987 => x"08",
          6988 => x"11",
          6989 => x"33",
          6990 => x"71",
          6991 => x"74",
          6992 => x"5c",
          6993 => x"84",
          6994 => x"85",
          6995 => x"ba",
          6996 => x"16",
          6997 => x"86",
          6998 => x"12",
          6999 => x"2b",
          7000 => x"2a",
          7001 => x"59",
          7002 => x"34",
          7003 => x"34",
          7004 => x"08",
          7005 => x"11",
          7006 => x"33",
          7007 => x"71",
          7008 => x"74",
          7009 => x"5c",
          7010 => x"86",
          7011 => x"87",
          7012 => x"ba",
          7013 => x"16",
          7014 => x"84",
          7015 => x"12",
          7016 => x"2b",
          7017 => x"2a",
          7018 => x"59",
          7019 => x"34",
          7020 => x"34",
          7021 => x"08",
          7022 => x"51",
          7023 => x"84",
          7024 => x"0d",
          7025 => x"33",
          7026 => x"71",
          7027 => x"83",
          7028 => x"05",
          7029 => x"85",
          7030 => x"88",
          7031 => x"88",
          7032 => x"59",
          7033 => x"74",
          7034 => x"76",
          7035 => x"84",
          7036 => x"70",
          7037 => x"33",
          7038 => x"71",
          7039 => x"83",
          7040 => x"05",
          7041 => x"87",
          7042 => x"88",
          7043 => x"88",
          7044 => x"5f",
          7045 => x"57",
          7046 => x"1a",
          7047 => x"1a",
          7048 => x"f4",
          7049 => x"33",
          7050 => x"71",
          7051 => x"81",
          7052 => x"70",
          7053 => x"57",
          7054 => x"77",
          7055 => x"18",
          7056 => x"f4",
          7057 => x"05",
          7058 => x"39",
          7059 => x"79",
          7060 => x"08",
          7061 => x"80",
          7062 => x"77",
          7063 => x"38",
          7064 => x"84",
          7065 => x"0d",
          7066 => x"fb",
          7067 => x"bb",
          7068 => x"bb",
          7069 => x"3d",
          7070 => x"ff",
          7071 => x"ba",
          7072 => x"80",
          7073 => x"f0",
          7074 => x"80",
          7075 => x"84",
          7076 => x"fe",
          7077 => x"84",
          7078 => x"55",
          7079 => x"81",
          7080 => x"34",
          7081 => x"08",
          7082 => x"15",
          7083 => x"85",
          7084 => x"ba",
          7085 => x"76",
          7086 => x"81",
          7087 => x"34",
          7088 => x"08",
          7089 => x"22",
          7090 => x"80",
          7091 => x"83",
          7092 => x"70",
          7093 => x"51",
          7094 => x"88",
          7095 => x"89",
          7096 => x"ba",
          7097 => x"10",
          7098 => x"ba",
          7099 => x"f8",
          7100 => x"76",
          7101 => x"81",
          7102 => x"34",
          7103 => x"80",
          7104 => x"38",
          7105 => x"ed",
          7106 => x"67",
          7107 => x"70",
          7108 => x"08",
          7109 => x"76",
          7110 => x"aa",
          7111 => x"2e",
          7112 => x"7f",
          7113 => x"d7",
          7114 => x"84",
          7115 => x"38",
          7116 => x"83",
          7117 => x"70",
          7118 => x"06",
          7119 => x"83",
          7120 => x"7f",
          7121 => x"2a",
          7122 => x"ff",
          7123 => x"2b",
          7124 => x"33",
          7125 => x"71",
          7126 => x"70",
          7127 => x"83",
          7128 => x"70",
          7129 => x"fc",
          7130 => x"2b",
          7131 => x"33",
          7132 => x"71",
          7133 => x"70",
          7134 => x"90",
          7135 => x"45",
          7136 => x"54",
          7137 => x"48",
          7138 => x"5f",
          7139 => x"24",
          7140 => x"82",
          7141 => x"16",
          7142 => x"2b",
          7143 => x"10",
          7144 => x"33",
          7145 => x"71",
          7146 => x"90",
          7147 => x"5c",
          7148 => x"56",
          7149 => x"85",
          7150 => x"62",
          7151 => x"38",
          7152 => x"77",
          7153 => x"a2",
          7154 => x"2e",
          7155 => x"60",
          7156 => x"62",
          7157 => x"38",
          7158 => x"61",
          7159 => x"f7",
          7160 => x"70",
          7161 => x"33",
          7162 => x"71",
          7163 => x"7a",
          7164 => x"81",
          7165 => x"98",
          7166 => x"2b",
          7167 => x"59",
          7168 => x"5b",
          7169 => x"24",
          7170 => x"76",
          7171 => x"33",
          7172 => x"71",
          7173 => x"83",
          7174 => x"11",
          7175 => x"87",
          7176 => x"8b",
          7177 => x"2b",
          7178 => x"84",
          7179 => x"15",
          7180 => x"2b",
          7181 => x"2a",
          7182 => x"52",
          7183 => x"53",
          7184 => x"77",
          7185 => x"79",
          7186 => x"84",
          7187 => x"70",
          7188 => x"33",
          7189 => x"71",
          7190 => x"83",
          7191 => x"05",
          7192 => x"87",
          7193 => x"88",
          7194 => x"88",
          7195 => x"5e",
          7196 => x"41",
          7197 => x"16",
          7198 => x"16",
          7199 => x"f4",
          7200 => x"33",
          7201 => x"71",
          7202 => x"81",
          7203 => x"70",
          7204 => x"5c",
          7205 => x"79",
          7206 => x"1a",
          7207 => x"f4",
          7208 => x"82",
          7209 => x"12",
          7210 => x"2b",
          7211 => x"07",
          7212 => x"33",
          7213 => x"71",
          7214 => x"70",
          7215 => x"5c",
          7216 => x"5a",
          7217 => x"79",
          7218 => x"1a",
          7219 => x"f4",
          7220 => x"70",
          7221 => x"33",
          7222 => x"71",
          7223 => x"74",
          7224 => x"33",
          7225 => x"71",
          7226 => x"70",
          7227 => x"5c",
          7228 => x"5a",
          7229 => x"82",
          7230 => x"83",
          7231 => x"ba",
          7232 => x"1f",
          7233 => x"83",
          7234 => x"88",
          7235 => x"57",
          7236 => x"83",
          7237 => x"5a",
          7238 => x"84",
          7239 => x"c3",
          7240 => x"ba",
          7241 => x"84",
          7242 => x"05",
          7243 => x"ff",
          7244 => x"44",
          7245 => x"26",
          7246 => x"7e",
          7247 => x"bb",
          7248 => x"3d",
          7249 => x"ff",
          7250 => x"ba",
          7251 => x"80",
          7252 => x"f0",
          7253 => x"80",
          7254 => x"84",
          7255 => x"fe",
          7256 => x"84",
          7257 => x"5e",
          7258 => x"81",
          7259 => x"34",
          7260 => x"08",
          7261 => x"1e",
          7262 => x"85",
          7263 => x"ba",
          7264 => x"60",
          7265 => x"81",
          7266 => x"34",
          7267 => x"08",
          7268 => x"22",
          7269 => x"80",
          7270 => x"83",
          7271 => x"70",
          7272 => x"5a",
          7273 => x"88",
          7274 => x"89",
          7275 => x"ba",
          7276 => x"10",
          7277 => x"ba",
          7278 => x"f8",
          7279 => x"60",
          7280 => x"81",
          7281 => x"34",
          7282 => x"08",
          7283 => x"d3",
          7284 => x"2e",
          7285 => x"7e",
          7286 => x"2e",
          7287 => x"7f",
          7288 => x"3f",
          7289 => x"08",
          7290 => x"0c",
          7291 => x"04",
          7292 => x"ba",
          7293 => x"83",
          7294 => x"5e",
          7295 => x"70",
          7296 => x"33",
          7297 => x"07",
          7298 => x"06",
          7299 => x"48",
          7300 => x"40",
          7301 => x"60",
          7302 => x"61",
          7303 => x"08",
          7304 => x"2a",
          7305 => x"82",
          7306 => x"83",
          7307 => x"ba",
          7308 => x"1f",
          7309 => x"12",
          7310 => x"2b",
          7311 => x"2b",
          7312 => x"06",
          7313 => x"83",
          7314 => x"70",
          7315 => x"5c",
          7316 => x"5b",
          7317 => x"82",
          7318 => x"81",
          7319 => x"60",
          7320 => x"34",
          7321 => x"08",
          7322 => x"7b",
          7323 => x"1c",
          7324 => x"ba",
          7325 => x"84",
          7326 => x"88",
          7327 => x"fd",
          7328 => x"75",
          7329 => x"ff",
          7330 => x"54",
          7331 => x"77",
          7332 => x"06",
          7333 => x"83",
          7334 => x"82",
          7335 => x"18",
          7336 => x"2b",
          7337 => x"10",
          7338 => x"33",
          7339 => x"71",
          7340 => x"90",
          7341 => x"5e",
          7342 => x"58",
          7343 => x"80",
          7344 => x"38",
          7345 => x"61",
          7346 => x"83",
          7347 => x"24",
          7348 => x"77",
          7349 => x"06",
          7350 => x"27",
          7351 => x"fe",
          7352 => x"ff",
          7353 => x"ba",
          7354 => x"80",
          7355 => x"f0",
          7356 => x"80",
          7357 => x"84",
          7358 => x"fe",
          7359 => x"84",
          7360 => x"5a",
          7361 => x"81",
          7362 => x"34",
          7363 => x"08",
          7364 => x"1a",
          7365 => x"85",
          7366 => x"ba",
          7367 => x"7e",
          7368 => x"81",
          7369 => x"34",
          7370 => x"08",
          7371 => x"22",
          7372 => x"80",
          7373 => x"83",
          7374 => x"70",
          7375 => x"56",
          7376 => x"64",
          7377 => x"73",
          7378 => x"34",
          7379 => x"22",
          7380 => x"10",
          7381 => x"08",
          7382 => x"42",
          7383 => x"82",
          7384 => x"61",
          7385 => x"fc",
          7386 => x"7a",
          7387 => x"38",
          7388 => x"ff",
          7389 => x"7b",
          7390 => x"38",
          7391 => x"76",
          7392 => x"bd",
          7393 => x"ea",
          7394 => x"54",
          7395 => x"84",
          7396 => x"0d",
          7397 => x"82",
          7398 => x"12",
          7399 => x"2b",
          7400 => x"07",
          7401 => x"11",
          7402 => x"33",
          7403 => x"71",
          7404 => x"7e",
          7405 => x"33",
          7406 => x"71",
          7407 => x"70",
          7408 => x"44",
          7409 => x"46",
          7410 => x"45",
          7411 => x"84",
          7412 => x"64",
          7413 => x"84",
          7414 => x"70",
          7415 => x"33",
          7416 => x"71",
          7417 => x"83",
          7418 => x"05",
          7419 => x"87",
          7420 => x"88",
          7421 => x"88",
          7422 => x"42",
          7423 => x"5d",
          7424 => x"86",
          7425 => x"64",
          7426 => x"84",
          7427 => x"16",
          7428 => x"12",
          7429 => x"2b",
          7430 => x"ff",
          7431 => x"2a",
          7432 => x"5d",
          7433 => x"79",
          7434 => x"84",
          7435 => x"70",
          7436 => x"33",
          7437 => x"71",
          7438 => x"83",
          7439 => x"05",
          7440 => x"15",
          7441 => x"2b",
          7442 => x"2a",
          7443 => x"40",
          7444 => x"54",
          7445 => x"75",
          7446 => x"84",
          7447 => x"70",
          7448 => x"81",
          7449 => x"8b",
          7450 => x"2b",
          7451 => x"82",
          7452 => x"15",
          7453 => x"2b",
          7454 => x"2a",
          7455 => x"5b",
          7456 => x"55",
          7457 => x"34",
          7458 => x"34",
          7459 => x"08",
          7460 => x"11",
          7461 => x"33",
          7462 => x"07",
          7463 => x"56",
          7464 => x"42",
          7465 => x"7e",
          7466 => x"51",
          7467 => x"3f",
          7468 => x"08",
          7469 => x"78",
          7470 => x"06",
          7471 => x"99",
          7472 => x"f4",
          7473 => x"f4",
          7474 => x"0b",
          7475 => x"23",
          7476 => x"53",
          7477 => x"ff",
          7478 => x"bf",
          7479 => x"ba",
          7480 => x"7f",
          7481 => x"0b",
          7482 => x"84",
          7483 => x"55",
          7484 => x"34",
          7485 => x"16",
          7486 => x"f4",
          7487 => x"86",
          7488 => x"0b",
          7489 => x"84",
          7490 => x"84",
          7491 => x"ff",
          7492 => x"80",
          7493 => x"ff",
          7494 => x"88",
          7495 => x"44",
          7496 => x"1f",
          7497 => x"1f",
          7498 => x"f0",
          7499 => x"10",
          7500 => x"f4",
          7501 => x"05",
          7502 => x"82",
          7503 => x"0b",
          7504 => x"7e",
          7505 => x"3f",
          7506 => x"c0",
          7507 => x"33",
          7508 => x"71",
          7509 => x"83",
          7510 => x"05",
          7511 => x"85",
          7512 => x"88",
          7513 => x"88",
          7514 => x"5e",
          7515 => x"76",
          7516 => x"34",
          7517 => x"05",
          7518 => x"f4",
          7519 => x"84",
          7520 => x"12",
          7521 => x"2b",
          7522 => x"07",
          7523 => x"14",
          7524 => x"33",
          7525 => x"07",
          7526 => x"41",
          7527 => x"59",
          7528 => x"79",
          7529 => x"34",
          7530 => x"05",
          7531 => x"f4",
          7532 => x"33",
          7533 => x"71",
          7534 => x"81",
          7535 => x"70",
          7536 => x"42",
          7537 => x"78",
          7538 => x"19",
          7539 => x"f4",
          7540 => x"70",
          7541 => x"33",
          7542 => x"71",
          7543 => x"74",
          7544 => x"81",
          7545 => x"88",
          7546 => x"83",
          7547 => x"f8",
          7548 => x"63",
          7549 => x"5d",
          7550 => x"40",
          7551 => x"7f",
          7552 => x"7b",
          7553 => x"84",
          7554 => x"70",
          7555 => x"81",
          7556 => x"8b",
          7557 => x"2b",
          7558 => x"70",
          7559 => x"33",
          7560 => x"07",
          7561 => x"06",
          7562 => x"48",
          7563 => x"46",
          7564 => x"60",
          7565 => x"60",
          7566 => x"61",
          7567 => x"06",
          7568 => x"39",
          7569 => x"87",
          7570 => x"8b",
          7571 => x"2b",
          7572 => x"84",
          7573 => x"19",
          7574 => x"2b",
          7575 => x"2a",
          7576 => x"52",
          7577 => x"84",
          7578 => x"85",
          7579 => x"ba",
          7580 => x"19",
          7581 => x"85",
          7582 => x"8b",
          7583 => x"2b",
          7584 => x"86",
          7585 => x"15",
          7586 => x"2b",
          7587 => x"2a",
          7588 => x"52",
          7589 => x"56",
          7590 => x"05",
          7591 => x"87",
          7592 => x"ba",
          7593 => x"70",
          7594 => x"33",
          7595 => x"07",
          7596 => x"06",
          7597 => x"5b",
          7598 => x"77",
          7599 => x"81",
          7600 => x"ba",
          7601 => x"1f",
          7602 => x"12",
          7603 => x"2b",
          7604 => x"07",
          7605 => x"33",
          7606 => x"71",
          7607 => x"70",
          7608 => x"ff",
          7609 => x"05",
          7610 => x"56",
          7611 => x"58",
          7612 => x"55",
          7613 => x"34",
          7614 => x"34",
          7615 => x"08",
          7616 => x"33",
          7617 => x"71",
          7618 => x"83",
          7619 => x"05",
          7620 => x"12",
          7621 => x"2b",
          7622 => x"ff",
          7623 => x"2a",
          7624 => x"58",
          7625 => x"55",
          7626 => x"76",
          7627 => x"84",
          7628 => x"70",
          7629 => x"33",
          7630 => x"71",
          7631 => x"83",
          7632 => x"11",
          7633 => x"87",
          7634 => x"8b",
          7635 => x"2b",
          7636 => x"84",
          7637 => x"15",
          7638 => x"2b",
          7639 => x"2a",
          7640 => x"52",
          7641 => x"53",
          7642 => x"57",
          7643 => x"34",
          7644 => x"34",
          7645 => x"08",
          7646 => x"11",
          7647 => x"33",
          7648 => x"71",
          7649 => x"74",
          7650 => x"33",
          7651 => x"71",
          7652 => x"70",
          7653 => x"42",
          7654 => x"57",
          7655 => x"86",
          7656 => x"87",
          7657 => x"ba",
          7658 => x"70",
          7659 => x"33",
          7660 => x"07",
          7661 => x"06",
          7662 => x"5a",
          7663 => x"76",
          7664 => x"81",
          7665 => x"ba",
          7666 => x"1f",
          7667 => x"83",
          7668 => x"8b",
          7669 => x"2b",
          7670 => x"73",
          7671 => x"33",
          7672 => x"07",
          7673 => x"41",
          7674 => x"5f",
          7675 => x"79",
          7676 => x"81",
          7677 => x"ba",
          7678 => x"1f",
          7679 => x"12",
          7680 => x"2b",
          7681 => x"07",
          7682 => x"14",
          7683 => x"33",
          7684 => x"07",
          7685 => x"41",
          7686 => x"5f",
          7687 => x"79",
          7688 => x"75",
          7689 => x"84",
          7690 => x"70",
          7691 => x"33",
          7692 => x"71",
          7693 => x"66",
          7694 => x"70",
          7695 => x"52",
          7696 => x"05",
          7697 => x"fe",
          7698 => x"84",
          7699 => x"1e",
          7700 => x"65",
          7701 => x"83",
          7702 => x"5d",
          7703 => x"d5",
          7704 => x"33",
          7705 => x"71",
          7706 => x"83",
          7707 => x"05",
          7708 => x"85",
          7709 => x"88",
          7710 => x"88",
          7711 => x"5d",
          7712 => x"7a",
          7713 => x"34",
          7714 => x"05",
          7715 => x"f4",
          7716 => x"84",
          7717 => x"12",
          7718 => x"2b",
          7719 => x"07",
          7720 => x"14",
          7721 => x"33",
          7722 => x"07",
          7723 => x"5b",
          7724 => x"5c",
          7725 => x"73",
          7726 => x"34",
          7727 => x"05",
          7728 => x"f4",
          7729 => x"33",
          7730 => x"71",
          7731 => x"81",
          7732 => x"70",
          7733 => x"5f",
          7734 => x"75",
          7735 => x"16",
          7736 => x"f4",
          7737 => x"70",
          7738 => x"33",
          7739 => x"71",
          7740 => x"74",
          7741 => x"81",
          7742 => x"88",
          7743 => x"83",
          7744 => x"f8",
          7745 => x"63",
          7746 => x"44",
          7747 => x"5e",
          7748 => x"74",
          7749 => x"7b",
          7750 => x"84",
          7751 => x"70",
          7752 => x"81",
          7753 => x"8b",
          7754 => x"2b",
          7755 => x"70",
          7756 => x"33",
          7757 => x"07",
          7758 => x"06",
          7759 => x"47",
          7760 => x"46",
          7761 => x"7f",
          7762 => x"81",
          7763 => x"83",
          7764 => x"5b",
          7765 => x"7e",
          7766 => x"e5",
          7767 => x"bb",
          7768 => x"84",
          7769 => x"80",
          7770 => x"62",
          7771 => x"84",
          7772 => x"51",
          7773 => x"3f",
          7774 => x"88",
          7775 => x"61",
          7776 => x"b7",
          7777 => x"39",
          7778 => x"7a",
          7779 => x"ba",
          7780 => x"58",
          7781 => x"b7",
          7782 => x"77",
          7783 => x"84",
          7784 => x"89",
          7785 => x"77",
          7786 => x"3f",
          7787 => x"08",
          7788 => x"84",
          7789 => x"e6",
          7790 => x"80",
          7791 => x"84",
          7792 => x"b5",
          7793 => x"84",
          7794 => x"89",
          7795 => x"84",
          7796 => x"84",
          7797 => x"a0",
          7798 => x"ba",
          7799 => x"80",
          7800 => x"52",
          7801 => x"51",
          7802 => x"3f",
          7803 => x"08",
          7804 => x"34",
          7805 => x"16",
          7806 => x"f4",
          7807 => x"84",
          7808 => x"0b",
          7809 => x"84",
          7810 => x"56",
          7811 => x"34",
          7812 => x"17",
          7813 => x"f4",
          7814 => x"f0",
          7815 => x"fe",
          7816 => x"70",
          7817 => x"06",
          7818 => x"58",
          7819 => x"74",
          7820 => x"73",
          7821 => x"84",
          7822 => x"70",
          7823 => x"84",
          7824 => x"05",
          7825 => x"55",
          7826 => x"34",
          7827 => x"15",
          7828 => x"77",
          7829 => x"c6",
          7830 => x"39",
          7831 => x"02",
          7832 => x"51",
          7833 => x"72",
          7834 => x"84",
          7835 => x"33",
          7836 => x"bb",
          7837 => x"3d",
          7838 => x"3d",
          7839 => x"05",
          7840 => x"53",
          7841 => x"9d",
          7842 => x"d4",
          7843 => x"bb",
          7844 => x"ff",
          7845 => x"87",
          7846 => x"bb",
          7847 => x"84",
          7848 => x"33",
          7849 => x"bb",
          7850 => x"3d",
          7851 => x"3d",
          7852 => x"60",
          7853 => x"af",
          7854 => x"5c",
          7855 => x"54",
          7856 => x"87",
          7857 => x"80",
          7858 => x"73",
          7859 => x"83",
          7860 => x"38",
          7861 => x"0b",
          7862 => x"8c",
          7863 => x"75",
          7864 => x"d5",
          7865 => x"bb",
          7866 => x"ff",
          7867 => x"80",
          7868 => x"87",
          7869 => x"08",
          7870 => x"38",
          7871 => x"d6",
          7872 => x"80",
          7873 => x"73",
          7874 => x"38",
          7875 => x"55",
          7876 => x"84",
          7877 => x"0d",
          7878 => x"16",
          7879 => x"81",
          7880 => x"55",
          7881 => x"26",
          7882 => x"d5",
          7883 => x"0d",
          7884 => x"02",
          7885 => x"05",
          7886 => x"57",
          7887 => x"76",
          7888 => x"38",
          7889 => x"17",
          7890 => x"81",
          7891 => x"55",
          7892 => x"73",
          7893 => x"87",
          7894 => x"0c",
          7895 => x"52",
          7896 => x"8e",
          7897 => x"84",
          7898 => x"06",
          7899 => x"2e",
          7900 => x"c0",
          7901 => x"54",
          7902 => x"79",
          7903 => x"38",
          7904 => x"80",
          7905 => x"80",
          7906 => x"81",
          7907 => x"74",
          7908 => x"0c",
          7909 => x"04",
          7910 => x"81",
          7911 => x"ff",
          7912 => x"56",
          7913 => x"ff",
          7914 => x"39",
          7915 => x"78",
          7916 => x"9b",
          7917 => x"88",
          7918 => x"33",
          7919 => x"81",
          7920 => x"26",
          7921 => x"bb",
          7922 => x"53",
          7923 => x"54",
          7924 => x"9b",
          7925 => x"87",
          7926 => x"0c",
          7927 => x"73",
          7928 => x"72",
          7929 => x"38",
          7930 => x"9a",
          7931 => x"72",
          7932 => x"0c",
          7933 => x"04",
          7934 => x"75",
          7935 => x"bb",
          7936 => x"3d",
          7937 => x"80",
          7938 => x"0b",
          7939 => x"0c",
          7940 => x"04",
          7941 => x"87",
          7942 => x"11",
          7943 => x"cd",
          7944 => x"70",
          7945 => x"06",
          7946 => x"80",
          7947 => x"87",
          7948 => x"08",
          7949 => x"38",
          7950 => x"8c",
          7951 => x"ca",
          7952 => x"0c",
          7953 => x"8c",
          7954 => x"08",
          7955 => x"73",
          7956 => x"9b",
          7957 => x"82",
          7958 => x"ee",
          7959 => x"39",
          7960 => x"7c",
          7961 => x"83",
          7962 => x"5b",
          7963 => x"77",
          7964 => x"06",
          7965 => x"33",
          7966 => x"2e",
          7967 => x"80",
          7968 => x"81",
          7969 => x"fe",
          7970 => x"bb",
          7971 => x"2e",
          7972 => x"59",
          7973 => x"84",
          7974 => x"0d",
          7975 => x"b4",
          7976 => x"b8",
          7977 => x"81",
          7978 => x"5a",
          7979 => x"81",
          7980 => x"84",
          7981 => x"09",
          7982 => x"38",
          7983 => x"08",
          7984 => x"b4",
          7985 => x"a8",
          7986 => x"a0",
          7987 => x"bb",
          7988 => x"58",
          7989 => x"76",
          7990 => x"38",
          7991 => x"55",
          7992 => x"09",
          7993 => x"8e",
          7994 => x"75",
          7995 => x"52",
          7996 => x"51",
          7997 => x"76",
          7998 => x"59",
          7999 => x"09",
          8000 => x"fb",
          8001 => x"33",
          8002 => x"2e",
          8003 => x"fe",
          8004 => x"18",
          8005 => x"7a",
          8006 => x"75",
          8007 => x"57",
          8008 => x"57",
          8009 => x"80",
          8010 => x"b6",
          8011 => x"aa",
          8012 => x"19",
          8013 => x"7a",
          8014 => x"0b",
          8015 => x"80",
          8016 => x"19",
          8017 => x"0b",
          8018 => x"80",
          8019 => x"9c",
          8020 => x"f2",
          8021 => x"19",
          8022 => x"0b",
          8023 => x"34",
          8024 => x"84",
          8025 => x"94",
          8026 => x"74",
          8027 => x"34",
          8028 => x"5b",
          8029 => x"19",
          8030 => x"2a",
          8031 => x"a2",
          8032 => x"98",
          8033 => x"84",
          8034 => x"90",
          8035 => x"7a",
          8036 => x"34",
          8037 => x"55",
          8038 => x"19",
          8039 => x"2a",
          8040 => x"a6",
          8041 => x"98",
          8042 => x"84",
          8043 => x"a4",
          8044 => x"05",
          8045 => x"0c",
          8046 => x"7a",
          8047 => x"81",
          8048 => x"fa",
          8049 => x"84",
          8050 => x"53",
          8051 => x"18",
          8052 => x"d8",
          8053 => x"84",
          8054 => x"fd",
          8055 => x"b2",
          8056 => x"0d",
          8057 => x"08",
          8058 => x"81",
          8059 => x"38",
          8060 => x"76",
          8061 => x"81",
          8062 => x"bb",
          8063 => x"3d",
          8064 => x"77",
          8065 => x"74",
          8066 => x"cc",
          8067 => x"24",
          8068 => x"74",
          8069 => x"81",
          8070 => x"75",
          8071 => x"70",
          8072 => x"19",
          8073 => x"5a",
          8074 => x"17",
          8075 => x"b0",
          8076 => x"33",
          8077 => x"2e",
          8078 => x"83",
          8079 => x"54",
          8080 => x"17",
          8081 => x"33",
          8082 => x"3f",
          8083 => x"08",
          8084 => x"38",
          8085 => x"5b",
          8086 => x"0c",
          8087 => x"38",
          8088 => x"06",
          8089 => x"33",
          8090 => x"89",
          8091 => x"08",
          8092 => x"5d",
          8093 => x"08",
          8094 => x"38",
          8095 => x"18",
          8096 => x"56",
          8097 => x"2e",
          8098 => x"84",
          8099 => x"54",
          8100 => x"17",
          8101 => x"33",
          8102 => x"3f",
          8103 => x"08",
          8104 => x"38",
          8105 => x"5a",
          8106 => x"0c",
          8107 => x"38",
          8108 => x"06",
          8109 => x"33",
          8110 => x"7e",
          8111 => x"06",
          8112 => x"53",
          8113 => x"5d",
          8114 => x"38",
          8115 => x"06",
          8116 => x"0c",
          8117 => x"04",
          8118 => x"a8",
          8119 => x"59",
          8120 => x"79",
          8121 => x"80",
          8122 => x"33",
          8123 => x"5b",
          8124 => x"09",
          8125 => x"c2",
          8126 => x"78",
          8127 => x"52",
          8128 => x"51",
          8129 => x"84",
          8130 => x"80",
          8131 => x"ff",
          8132 => x"78",
          8133 => x"79",
          8134 => x"75",
          8135 => x"06",
          8136 => x"05",
          8137 => x"71",
          8138 => x"2b",
          8139 => x"84",
          8140 => x"8f",
          8141 => x"74",
          8142 => x"81",
          8143 => x"38",
          8144 => x"a8",
          8145 => x"59",
          8146 => x"79",
          8147 => x"80",
          8148 => x"33",
          8149 => x"5b",
          8150 => x"09",
          8151 => x"81",
          8152 => x"78",
          8153 => x"52",
          8154 => x"51",
          8155 => x"84",
          8156 => x"80",
          8157 => x"ff",
          8158 => x"78",
          8159 => x"79",
          8160 => x"75",
          8161 => x"fc",
          8162 => x"b8",
          8163 => x"33",
          8164 => x"71",
          8165 => x"88",
          8166 => x"14",
          8167 => x"07",
          8168 => x"33",
          8169 => x"ff",
          8170 => x"07",
          8171 => x"0c",
          8172 => x"59",
          8173 => x"3d",
          8174 => x"54",
          8175 => x"53",
          8176 => x"53",
          8177 => x"52",
          8178 => x"3f",
          8179 => x"bb",
          8180 => x"2e",
          8181 => x"fe",
          8182 => x"bb",
          8183 => x"18",
          8184 => x"08",
          8185 => x"31",
          8186 => x"08",
          8187 => x"a0",
          8188 => x"fe",
          8189 => x"17",
          8190 => x"82",
          8191 => x"06",
          8192 => x"81",
          8193 => x"08",
          8194 => x"05",
          8195 => x"81",
          8196 => x"f6",
          8197 => x"5a",
          8198 => x"81",
          8199 => x"08",
          8200 => x"70",
          8201 => x"33",
          8202 => x"81",
          8203 => x"84",
          8204 => x"09",
          8205 => x"81",
          8206 => x"84",
          8207 => x"34",
          8208 => x"a8",
          8209 => x"5d",
          8210 => x"08",
          8211 => x"82",
          8212 => x"7d",
          8213 => x"cb",
          8214 => x"84",
          8215 => x"de",
          8216 => x"b4",
          8217 => x"b8",
          8218 => x"81",
          8219 => x"5c",
          8220 => x"81",
          8221 => x"84",
          8222 => x"09",
          8223 => x"ff",
          8224 => x"84",
          8225 => x"34",
          8226 => x"a8",
          8227 => x"84",
          8228 => x"5b",
          8229 => x"18",
          8230 => x"c5",
          8231 => x"33",
          8232 => x"2e",
          8233 => x"fd",
          8234 => x"54",
          8235 => x"a0",
          8236 => x"53",
          8237 => x"17",
          8238 => x"f1",
          8239 => x"fd",
          8240 => x"54",
          8241 => x"53",
          8242 => x"53",
          8243 => x"52",
          8244 => x"3f",
          8245 => x"bb",
          8246 => x"2e",
          8247 => x"fb",
          8248 => x"bb",
          8249 => x"18",
          8250 => x"08",
          8251 => x"31",
          8252 => x"08",
          8253 => x"a0",
          8254 => x"fb",
          8255 => x"17",
          8256 => x"82",
          8257 => x"06",
          8258 => x"81",
          8259 => x"08",
          8260 => x"05",
          8261 => x"81",
          8262 => x"f4",
          8263 => x"5a",
          8264 => x"81",
          8265 => x"08",
          8266 => x"05",
          8267 => x"81",
          8268 => x"f3",
          8269 => x"86",
          8270 => x"7a",
          8271 => x"fa",
          8272 => x"3d",
          8273 => x"64",
          8274 => x"82",
          8275 => x"27",
          8276 => x"9c",
          8277 => x"95",
          8278 => x"55",
          8279 => x"96",
          8280 => x"24",
          8281 => x"74",
          8282 => x"8a",
          8283 => x"bb",
          8284 => x"3d",
          8285 => x"88",
          8286 => x"08",
          8287 => x"0b",
          8288 => x"58",
          8289 => x"2e",
          8290 => x"83",
          8291 => x"5b",
          8292 => x"2e",
          8293 => x"83",
          8294 => x"54",
          8295 => x"19",
          8296 => x"33",
          8297 => x"3f",
          8298 => x"08",
          8299 => x"38",
          8300 => x"5a",
          8301 => x"0c",
          8302 => x"ff",
          8303 => x"10",
          8304 => x"79",
          8305 => x"ff",
          8306 => x"5e",
          8307 => x"34",
          8308 => x"5a",
          8309 => x"34",
          8310 => x"1a",
          8311 => x"bb",
          8312 => x"3d",
          8313 => x"83",
          8314 => x"06",
          8315 => x"75",
          8316 => x"1a",
          8317 => x"80",
          8318 => x"08",
          8319 => x"78",
          8320 => x"38",
          8321 => x"7c",
          8322 => x"7c",
          8323 => x"06",
          8324 => x"81",
          8325 => x"b8",
          8326 => x"19",
          8327 => x"8e",
          8328 => x"84",
          8329 => x"85",
          8330 => x"81",
          8331 => x"1a",
          8332 => x"79",
          8333 => x"75",
          8334 => x"fc",
          8335 => x"b8",
          8336 => x"33",
          8337 => x"8f",
          8338 => x"f0",
          8339 => x"41",
          8340 => x"7d",
          8341 => x"88",
          8342 => x"b9",
          8343 => x"90",
          8344 => x"ba",
          8345 => x"98",
          8346 => x"bb",
          8347 => x"0b",
          8348 => x"fe",
          8349 => x"81",
          8350 => x"89",
          8351 => x"08",
          8352 => x"08",
          8353 => x"76",
          8354 => x"38",
          8355 => x"1a",
          8356 => x"56",
          8357 => x"2e",
          8358 => x"82",
          8359 => x"54",
          8360 => x"19",
          8361 => x"33",
          8362 => x"3f",
          8363 => x"08",
          8364 => x"38",
          8365 => x"5c",
          8366 => x"0c",
          8367 => x"fd",
          8368 => x"83",
          8369 => x"b8",
          8370 => x"77",
          8371 => x"5f",
          8372 => x"7c",
          8373 => x"38",
          8374 => x"9f",
          8375 => x"33",
          8376 => x"07",
          8377 => x"77",
          8378 => x"83",
          8379 => x"89",
          8380 => x"08",
          8381 => x"0b",
          8382 => x"56",
          8383 => x"2e",
          8384 => x"81",
          8385 => x"b8",
          8386 => x"81",
          8387 => x"57",
          8388 => x"81",
          8389 => x"84",
          8390 => x"09",
          8391 => x"c7",
          8392 => x"84",
          8393 => x"34",
          8394 => x"70",
          8395 => x"31",
          8396 => x"84",
          8397 => x"5b",
          8398 => x"74",
          8399 => x"38",
          8400 => x"55",
          8401 => x"82",
          8402 => x"54",
          8403 => x"52",
          8404 => x"51",
          8405 => x"84",
          8406 => x"80",
          8407 => x"ff",
          8408 => x"75",
          8409 => x"77",
          8410 => x"7d",
          8411 => x"19",
          8412 => x"84",
          8413 => x"7c",
          8414 => x"88",
          8415 => x"81",
          8416 => x"8f",
          8417 => x"5c",
          8418 => x"81",
          8419 => x"34",
          8420 => x"81",
          8421 => x"b8",
          8422 => x"81",
          8423 => x"5d",
          8424 => x"81",
          8425 => x"84",
          8426 => x"09",
          8427 => x"88",
          8428 => x"84",
          8429 => x"34",
          8430 => x"70",
          8431 => x"31",
          8432 => x"84",
          8433 => x"5d",
          8434 => x"7e",
          8435 => x"ca",
          8436 => x"33",
          8437 => x"2e",
          8438 => x"fb",
          8439 => x"54",
          8440 => x"7c",
          8441 => x"33",
          8442 => x"3f",
          8443 => x"aa",
          8444 => x"76",
          8445 => x"70",
          8446 => x"33",
          8447 => x"ad",
          8448 => x"84",
          8449 => x"7d",
          8450 => x"06",
          8451 => x"84",
          8452 => x"83",
          8453 => x"19",
          8454 => x"1b",
          8455 => x"1b",
          8456 => x"84",
          8457 => x"56",
          8458 => x"27",
          8459 => x"82",
          8460 => x"74",
          8461 => x"81",
          8462 => x"38",
          8463 => x"1f",
          8464 => x"81",
          8465 => x"ed",
          8466 => x"5c",
          8467 => x"81",
          8468 => x"b8",
          8469 => x"81",
          8470 => x"57",
          8471 => x"81",
          8472 => x"84",
          8473 => x"09",
          8474 => x"c5",
          8475 => x"84",
          8476 => x"34",
          8477 => x"70",
          8478 => x"31",
          8479 => x"84",
          8480 => x"5d",
          8481 => x"7e",
          8482 => x"87",
          8483 => x"33",
          8484 => x"2e",
          8485 => x"fa",
          8486 => x"54",
          8487 => x"76",
          8488 => x"33",
          8489 => x"3f",
          8490 => x"e7",
          8491 => x"79",
          8492 => x"52",
          8493 => x"51",
          8494 => x"7e",
          8495 => x"39",
          8496 => x"83",
          8497 => x"05",
          8498 => x"ff",
          8499 => x"58",
          8500 => x"34",
          8501 => x"5a",
          8502 => x"34",
          8503 => x"7e",
          8504 => x"39",
          8505 => x"2b",
          8506 => x"7a",
          8507 => x"83",
          8508 => x"98",
          8509 => x"06",
          8510 => x"06",
          8511 => x"5f",
          8512 => x"7d",
          8513 => x"2a",
          8514 => x"1d",
          8515 => x"2a",
          8516 => x"1d",
          8517 => x"2a",
          8518 => x"1d",
          8519 => x"39",
          8520 => x"7c",
          8521 => x"5b",
          8522 => x"81",
          8523 => x"19",
          8524 => x"80",
          8525 => x"38",
          8526 => x"08",
          8527 => x"38",
          8528 => x"70",
          8529 => x"80",
          8530 => x"38",
          8531 => x"81",
          8532 => x"56",
          8533 => x"9c",
          8534 => x"26",
          8535 => x"56",
          8536 => x"82",
          8537 => x"52",
          8538 => x"f5",
          8539 => x"84",
          8540 => x"81",
          8541 => x"58",
          8542 => x"08",
          8543 => x"38",
          8544 => x"08",
          8545 => x"70",
          8546 => x"25",
          8547 => x"51",
          8548 => x"73",
          8549 => x"75",
          8550 => x"81",
          8551 => x"38",
          8552 => x"84",
          8553 => x"8c",
          8554 => x"81",
          8555 => x"39",
          8556 => x"08",
          8557 => x"7a",
          8558 => x"f0",
          8559 => x"55",
          8560 => x"84",
          8561 => x"38",
          8562 => x"08",
          8563 => x"84",
          8564 => x"ce",
          8565 => x"08",
          8566 => x"08",
          8567 => x"7a",
          8568 => x"39",
          8569 => x"9c",
          8570 => x"26",
          8571 => x"56",
          8572 => x"51",
          8573 => x"80",
          8574 => x"84",
          8575 => x"81",
          8576 => x"bb",
          8577 => x"70",
          8578 => x"07",
          8579 => x"7b",
          8580 => x"84",
          8581 => x"51",
          8582 => x"ff",
          8583 => x"bb",
          8584 => x"2e",
          8585 => x"19",
          8586 => x"74",
          8587 => x"38",
          8588 => x"08",
          8589 => x"38",
          8590 => x"57",
          8591 => x"75",
          8592 => x"8e",
          8593 => x"75",
          8594 => x"f5",
          8595 => x"bb",
          8596 => x"bb",
          8597 => x"70",
          8598 => x"08",
          8599 => x"56",
          8600 => x"80",
          8601 => x"80",
          8602 => x"90",
          8603 => x"19",
          8604 => x"94",
          8605 => x"58",
          8606 => x"86",
          8607 => x"94",
          8608 => x"19",
          8609 => x"5a",
          8610 => x"34",
          8611 => x"84",
          8612 => x"8c",
          8613 => x"80",
          8614 => x"84",
          8615 => x"0d",
          8616 => x"84",
          8617 => x"da",
          8618 => x"2e",
          8619 => x"75",
          8620 => x"78",
          8621 => x"3f",
          8622 => x"08",
          8623 => x"39",
          8624 => x"08",
          8625 => x"0c",
          8626 => x"04",
          8627 => x"81",
          8628 => x"38",
          8629 => x"b6",
          8630 => x"0d",
          8631 => x"08",
          8632 => x"73",
          8633 => x"26",
          8634 => x"73",
          8635 => x"72",
          8636 => x"73",
          8637 => x"88",
          8638 => x"74",
          8639 => x"76",
          8640 => x"82",
          8641 => x"38",
          8642 => x"53",
          8643 => x"18",
          8644 => x"72",
          8645 => x"38",
          8646 => x"98",
          8647 => x"94",
          8648 => x"18",
          8649 => x"56",
          8650 => x"94",
          8651 => x"2a",
          8652 => x"0c",
          8653 => x"06",
          8654 => x"9c",
          8655 => x"56",
          8656 => x"84",
          8657 => x"0d",
          8658 => x"84",
          8659 => x"8a",
          8660 => x"ac",
          8661 => x"74",
          8662 => x"ac",
          8663 => x"22",
          8664 => x"57",
          8665 => x"27",
          8666 => x"17",
          8667 => x"15",
          8668 => x"56",
          8669 => x"73",
          8670 => x"8a",
          8671 => x"71",
          8672 => x"08",
          8673 => x"78",
          8674 => x"ff",
          8675 => x"52",
          8676 => x"cd",
          8677 => x"84",
          8678 => x"bb",
          8679 => x"2e",
          8680 => x"0b",
          8681 => x"08",
          8682 => x"38",
          8683 => x"53",
          8684 => x"08",
          8685 => x"91",
          8686 => x"31",
          8687 => x"27",
          8688 => x"aa",
          8689 => x"84",
          8690 => x"8a",
          8691 => x"f3",
          8692 => x"70",
          8693 => x"08",
          8694 => x"5a",
          8695 => x"0a",
          8696 => x"38",
          8697 => x"18",
          8698 => x"08",
          8699 => x"74",
          8700 => x"38",
          8701 => x"06",
          8702 => x"38",
          8703 => x"18",
          8704 => x"75",
          8705 => x"85",
          8706 => x"22",
          8707 => x"76",
          8708 => x"38",
          8709 => x"0c",
          8710 => x"0c",
          8711 => x"05",
          8712 => x"80",
          8713 => x"bb",
          8714 => x"3d",
          8715 => x"98",
          8716 => x"19",
          8717 => x"7a",
          8718 => x"5c",
          8719 => x"75",
          8720 => x"eb",
          8721 => x"bb",
          8722 => x"82",
          8723 => x"84",
          8724 => x"27",
          8725 => x"56",
          8726 => x"08",
          8727 => x"38",
          8728 => x"84",
          8729 => x"26",
          8730 => x"60",
          8731 => x"98",
          8732 => x"08",
          8733 => x"f9",
          8734 => x"bb",
          8735 => x"87",
          8736 => x"84",
          8737 => x"ff",
          8738 => x"56",
          8739 => x"08",
          8740 => x"91",
          8741 => x"84",
          8742 => x"ff",
          8743 => x"38",
          8744 => x"08",
          8745 => x"5f",
          8746 => x"ea",
          8747 => x"9c",
          8748 => x"05",
          8749 => x"5c",
          8750 => x"8d",
          8751 => x"22",
          8752 => x"b0",
          8753 => x"5d",
          8754 => x"1a",
          8755 => x"58",
          8756 => x"57",
          8757 => x"70",
          8758 => x"34",
          8759 => x"74",
          8760 => x"56",
          8761 => x"55",
          8762 => x"81",
          8763 => x"54",
          8764 => x"77",
          8765 => x"33",
          8766 => x"3f",
          8767 => x"08",
          8768 => x"81",
          8769 => x"39",
          8770 => x"0c",
          8771 => x"bb",
          8772 => x"3d",
          8773 => x"54",
          8774 => x"53",
          8775 => x"53",
          8776 => x"52",
          8777 => x"3f",
          8778 => x"08",
          8779 => x"84",
          8780 => x"83",
          8781 => x"19",
          8782 => x"08",
          8783 => x"a0",
          8784 => x"fe",
          8785 => x"19",
          8786 => x"82",
          8787 => x"06",
          8788 => x"81",
          8789 => x"08",
          8790 => x"05",
          8791 => x"81",
          8792 => x"e3",
          8793 => x"c5",
          8794 => x"22",
          8795 => x"ff",
          8796 => x"74",
          8797 => x"81",
          8798 => x"7c",
          8799 => x"fe",
          8800 => x"08",
          8801 => x"56",
          8802 => x"7d",
          8803 => x"38",
          8804 => x"76",
          8805 => x"1b",
          8806 => x"19",
          8807 => x"f8",
          8808 => x"84",
          8809 => x"8f",
          8810 => x"ee",
          8811 => x"66",
          8812 => x"7c",
          8813 => x"81",
          8814 => x"1e",
          8815 => x"5e",
          8816 => x"82",
          8817 => x"19",
          8818 => x"80",
          8819 => x"08",
          8820 => x"d1",
          8821 => x"33",
          8822 => x"74",
          8823 => x"81",
          8824 => x"38",
          8825 => x"53",
          8826 => x"81",
          8827 => x"e1",
          8828 => x"bb",
          8829 => x"2e",
          8830 => x"5a",
          8831 => x"b4",
          8832 => x"5b",
          8833 => x"38",
          8834 => x"70",
          8835 => x"76",
          8836 => x"81",
          8837 => x"33",
          8838 => x"81",
          8839 => x"41",
          8840 => x"34",
          8841 => x"32",
          8842 => x"ae",
          8843 => x"72",
          8844 => x"80",
          8845 => x"45",
          8846 => x"74",
          8847 => x"7a",
          8848 => x"56",
          8849 => x"81",
          8850 => x"60",
          8851 => x"38",
          8852 => x"80",
          8853 => x"fa",
          8854 => x"bb",
          8855 => x"84",
          8856 => x"81",
          8857 => x"1c",
          8858 => x"fe",
          8859 => x"84",
          8860 => x"94",
          8861 => x"81",
          8862 => x"08",
          8863 => x"81",
          8864 => x"e1",
          8865 => x"57",
          8866 => x"08",
          8867 => x"81",
          8868 => x"38",
          8869 => x"08",
          8870 => x"b4",
          8871 => x"1a",
          8872 => x"bb",
          8873 => x"5b",
          8874 => x"08",
          8875 => x"38",
          8876 => x"41",
          8877 => x"09",
          8878 => x"a8",
          8879 => x"b4",
          8880 => x"1a",
          8881 => x"7e",
          8882 => x"33",
          8883 => x"3f",
          8884 => x"90",
          8885 => x"2e",
          8886 => x"81",
          8887 => x"86",
          8888 => x"5b",
          8889 => x"93",
          8890 => x"33",
          8891 => x"06",
          8892 => x"08",
          8893 => x"0c",
          8894 => x"76",
          8895 => x"38",
          8896 => x"74",
          8897 => x"39",
          8898 => x"60",
          8899 => x"06",
          8900 => x"c1",
          8901 => x"80",
          8902 => x"0c",
          8903 => x"84",
          8904 => x"0d",
          8905 => x"fd",
          8906 => x"18",
          8907 => x"77",
          8908 => x"06",
          8909 => x"19",
          8910 => x"33",
          8911 => x"71",
          8912 => x"58",
          8913 => x"ff",
          8914 => x"33",
          8915 => x"06",
          8916 => x"05",
          8917 => x"76",
          8918 => x"e7",
          8919 => x"78",
          8920 => x"33",
          8921 => x"88",
          8922 => x"44",
          8923 => x"2e",
          8924 => x"79",
          8925 => x"ff",
          8926 => x"10",
          8927 => x"5c",
          8928 => x"23",
          8929 => x"81",
          8930 => x"77",
          8931 => x"77",
          8932 => x"2a",
          8933 => x"57",
          8934 => x"90",
          8935 => x"fe",
          8936 => x"38",
          8937 => x"05",
          8938 => x"23",
          8939 => x"81",
          8940 => x"41",
          8941 => x"75",
          8942 => x"2e",
          8943 => x"ff",
          8944 => x"39",
          8945 => x"7c",
          8946 => x"74",
          8947 => x"81",
          8948 => x"78",
          8949 => x"5a",
          8950 => x"05",
          8951 => x"06",
          8952 => x"56",
          8953 => x"38",
          8954 => x"fd",
          8955 => x"0b",
          8956 => x"7a",
          8957 => x"0c",
          8958 => x"04",
          8959 => x"63",
          8960 => x"5c",
          8961 => x"51",
          8962 => x"84",
          8963 => x"5a",
          8964 => x"08",
          8965 => x"81",
          8966 => x"5d",
          8967 => x"1d",
          8968 => x"5e",
          8969 => x"56",
          8970 => x"1b",
          8971 => x"82",
          8972 => x"1b",
          8973 => x"55",
          8974 => x"09",
          8975 => x"df",
          8976 => x"75",
          8977 => x"52",
          8978 => x"51",
          8979 => x"84",
          8980 => x"80",
          8981 => x"ff",
          8982 => x"75",
          8983 => x"76",
          8984 => x"b2",
          8985 => x"08",
          8986 => x"59",
          8987 => x"84",
          8988 => x"19",
          8989 => x"70",
          8990 => x"57",
          8991 => x"1d",
          8992 => x"e5",
          8993 => x"38",
          8994 => x"81",
          8995 => x"8f",
          8996 => x"38",
          8997 => x"38",
          8998 => x"81",
          8999 => x"aa",
          9000 => x"56",
          9001 => x"74",
          9002 => x"81",
          9003 => x"78",
          9004 => x"5a",
          9005 => x"05",
          9006 => x"06",
          9007 => x"56",
          9008 => x"38",
          9009 => x"80",
          9010 => x"1c",
          9011 => x"57",
          9012 => x"8b",
          9013 => x"59",
          9014 => x"81",
          9015 => x"78",
          9016 => x"5a",
          9017 => x"31",
          9018 => x"58",
          9019 => x"80",
          9020 => x"38",
          9021 => x"e1",
          9022 => x"5d",
          9023 => x"1d",
          9024 => x"7b",
          9025 => x"3f",
          9026 => x"08",
          9027 => x"84",
          9028 => x"fe",
          9029 => x"84",
          9030 => x"93",
          9031 => x"81",
          9032 => x"08",
          9033 => x"81",
          9034 => x"dc",
          9035 => x"57",
          9036 => x"08",
          9037 => x"81",
          9038 => x"38",
          9039 => x"08",
          9040 => x"b4",
          9041 => x"1c",
          9042 => x"bb",
          9043 => x"59",
          9044 => x"08",
          9045 => x"38",
          9046 => x"5a",
          9047 => x"09",
          9048 => x"dd",
          9049 => x"b4",
          9050 => x"1c",
          9051 => x"7d",
          9052 => x"33",
          9053 => x"3f",
          9054 => x"c5",
          9055 => x"fd",
          9056 => x"1c",
          9057 => x"2a",
          9058 => x"55",
          9059 => x"38",
          9060 => x"81",
          9061 => x"80",
          9062 => x"8d",
          9063 => x"81",
          9064 => x"90",
          9065 => x"ac",
          9066 => x"5e",
          9067 => x"2e",
          9068 => x"ff",
          9069 => x"80",
          9070 => x"f4",
          9071 => x"bb",
          9072 => x"84",
          9073 => x"80",
          9074 => x"38",
          9075 => x"75",
          9076 => x"c2",
          9077 => x"5d",
          9078 => x"1d",
          9079 => x"39",
          9080 => x"57",
          9081 => x"09",
          9082 => x"38",
          9083 => x"9b",
          9084 => x"1b",
          9085 => x"2b",
          9086 => x"40",
          9087 => x"38",
          9088 => x"bf",
          9089 => x"f3",
          9090 => x"81",
          9091 => x"83",
          9092 => x"33",
          9093 => x"11",
          9094 => x"71",
          9095 => x"52",
          9096 => x"80",
          9097 => x"38",
          9098 => x"26",
          9099 => x"76",
          9100 => x"d1",
          9101 => x"84",
          9102 => x"61",
          9103 => x"53",
          9104 => x"5b",
          9105 => x"bd",
          9106 => x"bb",
          9107 => x"09",
          9108 => x"de",
          9109 => x"81",
          9110 => x"78",
          9111 => x"38",
          9112 => x"86",
          9113 => x"56",
          9114 => x"2e",
          9115 => x"80",
          9116 => x"79",
          9117 => x"70",
          9118 => x"7f",
          9119 => x"ff",
          9120 => x"ff",
          9121 => x"fe",
          9122 => x"0b",
          9123 => x"0c",
          9124 => x"04",
          9125 => x"ff",
          9126 => x"38",
          9127 => x"fe",
          9128 => x"3d",
          9129 => x"08",
          9130 => x"33",
          9131 => x"58",
          9132 => x"86",
          9133 => x"b5",
          9134 => x"1d",
          9135 => x"57",
          9136 => x"80",
          9137 => x"81",
          9138 => x"17",
          9139 => x"56",
          9140 => x"38",
          9141 => x"1f",
          9142 => x"60",
          9143 => x"55",
          9144 => x"05",
          9145 => x"70",
          9146 => x"34",
          9147 => x"74",
          9148 => x"80",
          9149 => x"70",
          9150 => x"56",
          9151 => x"82",
          9152 => x"c0",
          9153 => x"34",
          9154 => x"3d",
          9155 => x"1c",
          9156 => x"59",
          9157 => x"5a",
          9158 => x"70",
          9159 => x"33",
          9160 => x"05",
          9161 => x"15",
          9162 => x"38",
          9163 => x"80",
          9164 => x"79",
          9165 => x"74",
          9166 => x"38",
          9167 => x"5a",
          9168 => x"75",
          9169 => x"10",
          9170 => x"2a",
          9171 => x"ff",
          9172 => x"2a",
          9173 => x"58",
          9174 => x"80",
          9175 => x"76",
          9176 => x"32",
          9177 => x"58",
          9178 => x"d7",
          9179 => x"55",
          9180 => x"87",
          9181 => x"80",
          9182 => x"58",
          9183 => x"bf",
          9184 => x"75",
          9185 => x"87",
          9186 => x"76",
          9187 => x"ff",
          9188 => x"2a",
          9189 => x"76",
          9190 => x"1f",
          9191 => x"79",
          9192 => x"58",
          9193 => x"27",
          9194 => x"33",
          9195 => x"2e",
          9196 => x"16",
          9197 => x"27",
          9198 => x"75",
          9199 => x"56",
          9200 => x"2e",
          9201 => x"ea",
          9202 => x"56",
          9203 => x"87",
          9204 => x"98",
          9205 => x"ec",
          9206 => x"71",
          9207 => x"41",
          9208 => x"87",
          9209 => x"f4",
          9210 => x"f8",
          9211 => x"bb",
          9212 => x"38",
          9213 => x"80",
          9214 => x"fe",
          9215 => x"56",
          9216 => x"2e",
          9217 => x"84",
          9218 => x"56",
          9219 => x"08",
          9220 => x"81",
          9221 => x"38",
          9222 => x"05",
          9223 => x"34",
          9224 => x"84",
          9225 => x"05",
          9226 => x"75",
          9227 => x"06",
          9228 => x"7e",
          9229 => x"38",
          9230 => x"1d",
          9231 => x"e8",
          9232 => x"84",
          9233 => x"80",
          9234 => x"ed",
          9235 => x"bb",
          9236 => x"84",
          9237 => x"81",
          9238 => x"bb",
          9239 => x"19",
          9240 => x"1e",
          9241 => x"57",
          9242 => x"76",
          9243 => x"38",
          9244 => x"40",
          9245 => x"09",
          9246 => x"a3",
          9247 => x"75",
          9248 => x"52",
          9249 => x"51",
          9250 => x"84",
          9251 => x"80",
          9252 => x"ff",
          9253 => x"75",
          9254 => x"76",
          9255 => x"38",
          9256 => x"70",
          9257 => x"74",
          9258 => x"81",
          9259 => x"30",
          9260 => x"78",
          9261 => x"74",
          9262 => x"c9",
          9263 => x"59",
          9264 => x"86",
          9265 => x"52",
          9266 => x"83",
          9267 => x"84",
          9268 => x"bb",
          9269 => x"2e",
          9270 => x"87",
          9271 => x"2e",
          9272 => x"75",
          9273 => x"83",
          9274 => x"40",
          9275 => x"38",
          9276 => x"57",
          9277 => x"77",
          9278 => x"83",
          9279 => x"57",
          9280 => x"82",
          9281 => x"76",
          9282 => x"52",
          9283 => x"51",
          9284 => x"84",
          9285 => x"80",
          9286 => x"ff",
          9287 => x"76",
          9288 => x"75",
          9289 => x"c3",
          9290 => x"9c",
          9291 => x"55",
          9292 => x"81",
          9293 => x"ff",
          9294 => x"f4",
          9295 => x"9c",
          9296 => x"58",
          9297 => x"70",
          9298 => x"33",
          9299 => x"05",
          9300 => x"15",
          9301 => x"38",
          9302 => x"ab",
          9303 => x"06",
          9304 => x"8c",
          9305 => x"0b",
          9306 => x"77",
          9307 => x"bb",
          9308 => x"3d",
          9309 => x"75",
          9310 => x"25",
          9311 => x"40",
          9312 => x"b9",
          9313 => x"81",
          9314 => x"ec",
          9315 => x"bb",
          9316 => x"84",
          9317 => x"80",
          9318 => x"38",
          9319 => x"81",
          9320 => x"08",
          9321 => x"81",
          9322 => x"d3",
          9323 => x"bb",
          9324 => x"2e",
          9325 => x"83",
          9326 => x"bb",
          9327 => x"19",
          9328 => x"08",
          9329 => x"31",
          9330 => x"19",
          9331 => x"38",
          9332 => x"41",
          9333 => x"84",
          9334 => x"bb",
          9335 => x"fd",
          9336 => x"85",
          9337 => x"08",
          9338 => x"58",
          9339 => x"e9",
          9340 => x"84",
          9341 => x"bb",
          9342 => x"ef",
          9343 => x"bb",
          9344 => x"58",
          9345 => x"81",
          9346 => x"80",
          9347 => x"70",
          9348 => x"33",
          9349 => x"70",
          9350 => x"ff",
          9351 => x"5d",
          9352 => x"74",
          9353 => x"b8",
          9354 => x"98",
          9355 => x"80",
          9356 => x"08",
          9357 => x"38",
          9358 => x"5b",
          9359 => x"09",
          9360 => x"c9",
          9361 => x"76",
          9362 => x"52",
          9363 => x"51",
          9364 => x"84",
          9365 => x"80",
          9366 => x"ff",
          9367 => x"76",
          9368 => x"75",
          9369 => x"83",
          9370 => x"08",
          9371 => x"61",
          9372 => x"5f",
          9373 => x"8d",
          9374 => x"0b",
          9375 => x"75",
          9376 => x"75",
          9377 => x"75",
          9378 => x"7c",
          9379 => x"05",
          9380 => x"58",
          9381 => x"ff",
          9382 => x"38",
          9383 => x"70",
          9384 => x"5b",
          9385 => x"e7",
          9386 => x"7b",
          9387 => x"75",
          9388 => x"57",
          9389 => x"2a",
          9390 => x"34",
          9391 => x"83",
          9392 => x"81",
          9393 => x"78",
          9394 => x"76",
          9395 => x"2e",
          9396 => x"78",
          9397 => x"22",
          9398 => x"80",
          9399 => x"38",
          9400 => x"81",
          9401 => x"34",
          9402 => x"51",
          9403 => x"84",
          9404 => x"58",
          9405 => x"08",
          9406 => x"7f",
          9407 => x"7f",
          9408 => x"fb",
          9409 => x"54",
          9410 => x"53",
          9411 => x"53",
          9412 => x"52",
          9413 => x"3f",
          9414 => x"bb",
          9415 => x"83",
          9416 => x"84",
          9417 => x"34",
          9418 => x"a8",
          9419 => x"84",
          9420 => x"57",
          9421 => x"1d",
          9422 => x"c9",
          9423 => x"33",
          9424 => x"2e",
          9425 => x"fb",
          9426 => x"54",
          9427 => x"a0",
          9428 => x"53",
          9429 => x"1c",
          9430 => x"d1",
          9431 => x"fb",
          9432 => x"9c",
          9433 => x"33",
          9434 => x"74",
          9435 => x"09",
          9436 => x"ba",
          9437 => x"39",
          9438 => x"57",
          9439 => x"fa",
          9440 => x"d7",
          9441 => x"c0",
          9442 => x"d4",
          9443 => x"b4",
          9444 => x"61",
          9445 => x"33",
          9446 => x"3f",
          9447 => x"08",
          9448 => x"81",
          9449 => x"84",
          9450 => x"83",
          9451 => x"1c",
          9452 => x"08",
          9453 => x"a0",
          9454 => x"8a",
          9455 => x"33",
          9456 => x"2e",
          9457 => x"bb",
          9458 => x"fc",
          9459 => x"ff",
          9460 => x"7f",
          9461 => x"98",
          9462 => x"39",
          9463 => x"f7",
          9464 => x"70",
          9465 => x"80",
          9466 => x"38",
          9467 => x"81",
          9468 => x"08",
          9469 => x"05",
          9470 => x"81",
          9471 => x"ce",
          9472 => x"c1",
          9473 => x"b4",
          9474 => x"19",
          9475 => x"7c",
          9476 => x"33",
          9477 => x"3f",
          9478 => x"f3",
          9479 => x"61",
          9480 => x"5e",
          9481 => x"96",
          9482 => x"1c",
          9483 => x"82",
          9484 => x"1c",
          9485 => x"80",
          9486 => x"70",
          9487 => x"05",
          9488 => x"57",
          9489 => x"58",
          9490 => x"bc",
          9491 => x"74",
          9492 => x"81",
          9493 => x"56",
          9494 => x"38",
          9495 => x"14",
          9496 => x"ff",
          9497 => x"76",
          9498 => x"82",
          9499 => x"79",
          9500 => x"70",
          9501 => x"55",
          9502 => x"38",
          9503 => x"80",
          9504 => x"7a",
          9505 => x"5e",
          9506 => x"05",
          9507 => x"82",
          9508 => x"70",
          9509 => x"57",
          9510 => x"08",
          9511 => x"81",
          9512 => x"53",
          9513 => x"b2",
          9514 => x"2e",
          9515 => x"75",
          9516 => x"30",
          9517 => x"80",
          9518 => x"54",
          9519 => x"90",
          9520 => x"2e",
          9521 => x"77",
          9522 => x"59",
          9523 => x"58",
          9524 => x"81",
          9525 => x"81",
          9526 => x"76",
          9527 => x"38",
          9528 => x"05",
          9529 => x"81",
          9530 => x"1d",
          9531 => x"a5",
          9532 => x"f3",
          9533 => x"96",
          9534 => x"57",
          9535 => x"05",
          9536 => x"82",
          9537 => x"1c",
          9538 => x"33",
          9539 => x"89",
          9540 => x"1e",
          9541 => x"08",
          9542 => x"33",
          9543 => x"9c",
          9544 => x"11",
          9545 => x"82",
          9546 => x"90",
          9547 => x"2b",
          9548 => x"33",
          9549 => x"88",
          9550 => x"71",
          9551 => x"59",
          9552 => x"96",
          9553 => x"88",
          9554 => x"41",
          9555 => x"56",
          9556 => x"86",
          9557 => x"15",
          9558 => x"33",
          9559 => x"07",
          9560 => x"84",
          9561 => x"3d",
          9562 => x"e5",
          9563 => x"39",
          9564 => x"11",
          9565 => x"31",
          9566 => x"83",
          9567 => x"90",
          9568 => x"51",
          9569 => x"3f",
          9570 => x"08",
          9571 => x"06",
          9572 => x"75",
          9573 => x"81",
          9574 => x"b3",
          9575 => x"2a",
          9576 => x"34",
          9577 => x"34",
          9578 => x"58",
          9579 => x"1f",
          9580 => x"78",
          9581 => x"70",
          9582 => x"54",
          9583 => x"38",
          9584 => x"74",
          9585 => x"70",
          9586 => x"25",
          9587 => x"07",
          9588 => x"75",
          9589 => x"74",
          9590 => x"78",
          9591 => x"0b",
          9592 => x"56",
          9593 => x"72",
          9594 => x"33",
          9595 => x"77",
          9596 => x"88",
          9597 => x"1e",
          9598 => x"54",
          9599 => x"ff",
          9600 => x"54",
          9601 => x"a4",
          9602 => x"08",
          9603 => x"54",
          9604 => x"27",
          9605 => x"84",
          9606 => x"81",
          9607 => x"80",
          9608 => x"a0",
          9609 => x"ff",
          9610 => x"53",
          9611 => x"81",
          9612 => x"81",
          9613 => x"81",
          9614 => x"13",
          9615 => x"59",
          9616 => x"ff",
          9617 => x"b4",
          9618 => x"2a",
          9619 => x"80",
          9620 => x"80",
          9621 => x"73",
          9622 => x"5f",
          9623 => x"39",
          9624 => x"63",
          9625 => x"42",
          9626 => x"65",
          9627 => x"55",
          9628 => x"2e",
          9629 => x"53",
          9630 => x"2e",
          9631 => x"72",
          9632 => x"d9",
          9633 => x"08",
          9634 => x"73",
          9635 => x"94",
          9636 => x"55",
          9637 => x"82",
          9638 => x"42",
          9639 => x"58",
          9640 => x"70",
          9641 => x"52",
          9642 => x"73",
          9643 => x"72",
          9644 => x"ff",
          9645 => x"38",
          9646 => x"74",
          9647 => x"76",
          9648 => x"80",
          9649 => x"17",
          9650 => x"ff",
          9651 => x"af",
          9652 => x"9f",
          9653 => x"80",
          9654 => x"5b",
          9655 => x"82",
          9656 => x"80",
          9657 => x"89",
          9658 => x"ff",
          9659 => x"83",
          9660 => x"83",
          9661 => x"70",
          9662 => x"56",
          9663 => x"80",
          9664 => x"38",
          9665 => x"8f",
          9666 => x"70",
          9667 => x"ff",
          9668 => x"56",
          9669 => x"72",
          9670 => x"5b",
          9671 => x"38",
          9672 => x"26",
          9673 => x"76",
          9674 => x"74",
          9675 => x"17",
          9676 => x"81",
          9677 => x"56",
          9678 => x"80",
          9679 => x"38",
          9680 => x"81",
          9681 => x"32",
          9682 => x"80",
          9683 => x"51",
          9684 => x"72",
          9685 => x"38",
          9686 => x"46",
          9687 => x"33",
          9688 => x"af",
          9689 => x"72",
          9690 => x"70",
          9691 => x"25",
          9692 => x"54",
          9693 => x"38",
          9694 => x"0c",
          9695 => x"3d",
          9696 => x"42",
          9697 => x"26",
          9698 => x"b4",
          9699 => x"52",
          9700 => x"8d",
          9701 => x"bb",
          9702 => x"ff",
          9703 => x"73",
          9704 => x"86",
          9705 => x"bb",
          9706 => x"3d",
          9707 => x"e6",
          9708 => x"81",
          9709 => x"53",
          9710 => x"fe",
          9711 => x"39",
          9712 => x"ab",
          9713 => x"52",
          9714 => x"8d",
          9715 => x"84",
          9716 => x"84",
          9717 => x"0d",
          9718 => x"80",
          9719 => x"30",
          9720 => x"73",
          9721 => x"5a",
          9722 => x"2e",
          9723 => x"14",
          9724 => x"70",
          9725 => x"56",
          9726 => x"dd",
          9727 => x"dc",
          9728 => x"70",
          9729 => x"07",
          9730 => x"7d",
          9731 => x"61",
          9732 => x"27",
          9733 => x"76",
          9734 => x"f8",
          9735 => x"2e",
          9736 => x"76",
          9737 => x"80",
          9738 => x"76",
          9739 => x"fe",
          9740 => x"70",
          9741 => x"30",
          9742 => x"52",
          9743 => x"56",
          9744 => x"2e",
          9745 => x"89",
          9746 => x"57",
          9747 => x"76",
          9748 => x"56",
          9749 => x"76",
          9750 => x"c7",
          9751 => x"22",
          9752 => x"ff",
          9753 => x"5d",
          9754 => x"a0",
          9755 => x"38",
          9756 => x"ff",
          9757 => x"ae",
          9758 => x"38",
          9759 => x"aa",
          9760 => x"fe",
          9761 => x"5a",
          9762 => x"2e",
          9763 => x"10",
          9764 => x"54",
          9765 => x"76",
          9766 => x"38",
          9767 => x"22",
          9768 => x"ae",
          9769 => x"06",
          9770 => x"0b",
          9771 => x"53",
          9772 => x"81",
          9773 => x"ff",
          9774 => x"f4",
          9775 => x"5c",
          9776 => x"16",
          9777 => x"19",
          9778 => x"5d",
          9779 => x"80",
          9780 => x"a0",
          9781 => x"38",
          9782 => x"70",
          9783 => x"25",
          9784 => x"75",
          9785 => x"ce",
          9786 => x"bb",
          9787 => x"7c",
          9788 => x"38",
          9789 => x"77",
          9790 => x"70",
          9791 => x"25",
          9792 => x"51",
          9793 => x"72",
          9794 => x"e0",
          9795 => x"2e",
          9796 => x"75",
          9797 => x"38",
          9798 => x"5a",
          9799 => x"9e",
          9800 => x"88",
          9801 => x"82",
          9802 => x"06",
          9803 => x"5f",
          9804 => x"70",
          9805 => x"58",
          9806 => x"ff",
          9807 => x"1c",
          9808 => x"81",
          9809 => x"84",
          9810 => x"2e",
          9811 => x"7d",
          9812 => x"77",
          9813 => x"ed",
          9814 => x"06",
          9815 => x"2e",
          9816 => x"79",
          9817 => x"06",
          9818 => x"38",
          9819 => x"5d",
          9820 => x"85",
          9821 => x"07",
          9822 => x"2a",
          9823 => x"7d",
          9824 => x"38",
          9825 => x"5a",
          9826 => x"34",
          9827 => x"ec",
          9828 => x"84",
          9829 => x"33",
          9830 => x"bb",
          9831 => x"2e",
          9832 => x"84",
          9833 => x"84",
          9834 => x"06",
          9835 => x"74",
          9836 => x"06",
          9837 => x"2e",
          9838 => x"74",
          9839 => x"06",
          9840 => x"98",
          9841 => x"65",
          9842 => x"42",
          9843 => x"58",
          9844 => x"ce",
          9845 => x"70",
          9846 => x"70",
          9847 => x"56",
          9848 => x"2e",
          9849 => x"80",
          9850 => x"38",
          9851 => x"5a",
          9852 => x"82",
          9853 => x"75",
          9854 => x"81",
          9855 => x"38",
          9856 => x"73",
          9857 => x"81",
          9858 => x"38",
          9859 => x"5b",
          9860 => x"80",
          9861 => x"56",
          9862 => x"76",
          9863 => x"38",
          9864 => x"75",
          9865 => x"57",
          9866 => x"53",
          9867 => x"e9",
          9868 => x"07",
          9869 => x"1d",
          9870 => x"e3",
          9871 => x"bb",
          9872 => x"1d",
          9873 => x"84",
          9874 => x"fe",
          9875 => x"82",
          9876 => x"58",
          9877 => x"38",
          9878 => x"70",
          9879 => x"06",
          9880 => x"80",
          9881 => x"38",
          9882 => x"83",
          9883 => x"05",
          9884 => x"33",
          9885 => x"33",
          9886 => x"07",
          9887 => x"57",
          9888 => x"83",
          9889 => x"38",
          9890 => x"0c",
          9891 => x"55",
          9892 => x"39",
          9893 => x"74",
          9894 => x"f0",
          9895 => x"59",
          9896 => x"38",
          9897 => x"79",
          9898 => x"17",
          9899 => x"81",
          9900 => x"2b",
          9901 => x"70",
          9902 => x"5e",
          9903 => x"09",
          9904 => x"95",
          9905 => x"07",
          9906 => x"39",
          9907 => x"1d",
          9908 => x"2e",
          9909 => x"fc",
          9910 => x"39",
          9911 => x"ab",
          9912 => x"0b",
          9913 => x"0c",
          9914 => x"04",
          9915 => x"26",
          9916 => x"ff",
          9917 => x"c9",
          9918 => x"59",
          9919 => x"81",
          9920 => x"83",
          9921 => x"18",
          9922 => x"fc",
          9923 => x"82",
          9924 => x"b5",
          9925 => x"81",
          9926 => x"84",
          9927 => x"83",
          9928 => x"70",
          9929 => x"06",
          9930 => x"80",
          9931 => x"74",
          9932 => x"83",
          9933 => x"33",
          9934 => x"81",
          9935 => x"b9",
          9936 => x"2e",
          9937 => x"83",
          9938 => x"83",
          9939 => x"70",
          9940 => x"56",
          9941 => x"80",
          9942 => x"38",
          9943 => x"8f",
          9944 => x"70",
          9945 => x"ff",
          9946 => x"59",
          9947 => x"72",
          9948 => x"59",
          9949 => x"38",
          9950 => x"54",
          9951 => x"8a",
          9952 => x"07",
          9953 => x"06",
          9954 => x"9f",
          9955 => x"99",
          9956 => x"7d",
          9957 => x"81",
          9958 => x"17",
          9959 => x"ff",
          9960 => x"5f",
          9961 => x"a0",
          9962 => x"79",
          9963 => x"5b",
          9964 => x"fa",
          9965 => x"53",
          9966 => x"83",
          9967 => x"70",
          9968 => x"5a",
          9969 => x"2e",
          9970 => x"80",
          9971 => x"07",
          9972 => x"05",
          9973 => x"74",
          9974 => x"1b",
          9975 => x"80",
          9976 => x"80",
          9977 => x"71",
          9978 => x"90",
          9979 => x"07",
          9980 => x"5a",
          9981 => x"39",
          9982 => x"05",
          9983 => x"54",
          9984 => x"34",
          9985 => x"11",
          9986 => x"5b",
          9987 => x"81",
          9988 => x"9c",
          9989 => x"07",
          9990 => x"58",
          9991 => x"e5",
          9992 => x"06",
          9993 => x"fd",
          9994 => x"82",
          9995 => x"5c",
          9996 => x"38",
          9997 => x"bb",
          9998 => x"3d",
          9999 => x"3d",
         10000 => x"02",
         10001 => x"e7",
         10002 => x"42",
         10003 => x"0c",
         10004 => x"70",
         10005 => x"79",
         10006 => x"d7",
         10007 => x"81",
         10008 => x"70",
         10009 => x"56",
         10010 => x"85",
         10011 => x"ed",
         10012 => x"2e",
         10013 => x"84",
         10014 => x"56",
         10015 => x"85",
         10016 => x"10",
         10017 => x"cc",
         10018 => x"58",
         10019 => x"76",
         10020 => x"96",
         10021 => x"0c",
         10022 => x"06",
         10023 => x"59",
         10024 => x"9b",
         10025 => x"33",
         10026 => x"b0",
         10027 => x"84",
         10028 => x"06",
         10029 => x"5e",
         10030 => x"2e",
         10031 => x"80",
         10032 => x"16",
         10033 => x"f8",
         10034 => x"18",
         10035 => x"81",
         10036 => x"ff",
         10037 => x"84",
         10038 => x"81",
         10039 => x"81",
         10040 => x"83",
         10041 => x"c2",
         10042 => x"2e",
         10043 => x"82",
         10044 => x"41",
         10045 => x"84",
         10046 => x"5b",
         10047 => x"34",
         10048 => x"18",
         10049 => x"5a",
         10050 => x"7a",
         10051 => x"70",
         10052 => x"33",
         10053 => x"bb",
         10054 => x"bb",
         10055 => x"2e",
         10056 => x"55",
         10057 => x"b4",
         10058 => x"56",
         10059 => x"84",
         10060 => x"84",
         10061 => x"71",
         10062 => x"56",
         10063 => x"74",
         10064 => x"2e",
         10065 => x"75",
         10066 => x"38",
         10067 => x"1d",
         10068 => x"85",
         10069 => x"58",
         10070 => x"83",
         10071 => x"58",
         10072 => x"83",
         10073 => x"c4",
         10074 => x"c3",
         10075 => x"88",
         10076 => x"59",
         10077 => x"2e",
         10078 => x"83",
         10079 => x"cf",
         10080 => x"ce",
         10081 => x"88",
         10082 => x"5a",
         10083 => x"80",
         10084 => x"11",
         10085 => x"33",
         10086 => x"71",
         10087 => x"81",
         10088 => x"72",
         10089 => x"75",
         10090 => x"56",
         10091 => x"5e",
         10092 => x"a0",
         10093 => x"c8",
         10094 => x"18",
         10095 => x"17",
         10096 => x"70",
         10097 => x"5f",
         10098 => x"58",
         10099 => x"82",
         10100 => x"81",
         10101 => x"71",
         10102 => x"19",
         10103 => x"5a",
         10104 => x"23",
         10105 => x"80",
         10106 => x"38",
         10107 => x"06",
         10108 => x"bb",
         10109 => x"17",
         10110 => x"18",
         10111 => x"2b",
         10112 => x"74",
         10113 => x"74",
         10114 => x"5e",
         10115 => x"7c",
         10116 => x"80",
         10117 => x"80",
         10118 => x"71",
         10119 => x"56",
         10120 => x"38",
         10121 => x"83",
         10122 => x"12",
         10123 => x"2b",
         10124 => x"07",
         10125 => x"70",
         10126 => x"2b",
         10127 => x"07",
         10128 => x"58",
         10129 => x"80",
         10130 => x"80",
         10131 => x"71",
         10132 => x"5d",
         10133 => x"7b",
         10134 => x"ce",
         10135 => x"7a",
         10136 => x"5a",
         10137 => x"81",
         10138 => x"52",
         10139 => x"51",
         10140 => x"3f",
         10141 => x"08",
         10142 => x"84",
         10143 => x"81",
         10144 => x"bb",
         10145 => x"ff",
         10146 => x"26",
         10147 => x"5d",
         10148 => x"f5",
         10149 => x"82",
         10150 => x"f5",
         10151 => x"38",
         10152 => x"16",
         10153 => x"0c",
         10154 => x"0c",
         10155 => x"a8",
         10156 => x"1d",
         10157 => x"57",
         10158 => x"2e",
         10159 => x"88",
         10160 => x"8d",
         10161 => x"2e",
         10162 => x"7d",
         10163 => x"0c",
         10164 => x"7c",
         10165 => x"38",
         10166 => x"70",
         10167 => x"81",
         10168 => x"5a",
         10169 => x"89",
         10170 => x"58",
         10171 => x"08",
         10172 => x"ff",
         10173 => x"0c",
         10174 => x"18",
         10175 => x"0b",
         10176 => x"7c",
         10177 => x"96",
         10178 => x"34",
         10179 => x"22",
         10180 => x"7c",
         10181 => x"23",
         10182 => x"23",
         10183 => x"0b",
         10184 => x"80",
         10185 => x"0c",
         10186 => x"84",
         10187 => x"97",
         10188 => x"8b",
         10189 => x"84",
         10190 => x"0d",
         10191 => x"d0",
         10192 => x"ff",
         10193 => x"58",
         10194 => x"91",
         10195 => x"78",
         10196 => x"d0",
         10197 => x"78",
         10198 => x"fe",
         10199 => x"08",
         10200 => x"5f",
         10201 => x"08",
         10202 => x"7a",
         10203 => x"5c",
         10204 => x"81",
         10205 => x"ff",
         10206 => x"58",
         10207 => x"26",
         10208 => x"16",
         10209 => x"06",
         10210 => x"9f",
         10211 => x"99",
         10212 => x"e0",
         10213 => x"ff",
         10214 => x"75",
         10215 => x"2a",
         10216 => x"77",
         10217 => x"06",
         10218 => x"ff",
         10219 => x"7a",
         10220 => x"70",
         10221 => x"2a",
         10222 => x"58",
         10223 => x"2e",
         10224 => x"81",
         10225 => x"5e",
         10226 => x"25",
         10227 => x"61",
         10228 => x"39",
         10229 => x"fe",
         10230 => x"82",
         10231 => x"5e",
         10232 => x"fe",
         10233 => x"58",
         10234 => x"7a",
         10235 => x"59",
         10236 => x"2e",
         10237 => x"83",
         10238 => x"75",
         10239 => x"70",
         10240 => x"25",
         10241 => x"5b",
         10242 => x"ad",
         10243 => x"e8",
         10244 => x"38",
         10245 => x"57",
         10246 => x"83",
         10247 => x"70",
         10248 => x"80",
         10249 => x"84",
         10250 => x"84",
         10251 => x"71",
         10252 => x"88",
         10253 => x"ff",
         10254 => x"72",
         10255 => x"83",
         10256 => x"71",
         10257 => x"5b",
         10258 => x"77",
         10259 => x"05",
         10260 => x"19",
         10261 => x"59",
         10262 => x"ff",
         10263 => x"ba",
         10264 => x"70",
         10265 => x"2a",
         10266 => x"9b",
         10267 => x"10",
         10268 => x"84",
         10269 => x"5d",
         10270 => x"42",
         10271 => x"83",
         10272 => x"2e",
         10273 => x"80",
         10274 => x"34",
         10275 => x"18",
         10276 => x"80",
         10277 => x"2e",
         10278 => x"54",
         10279 => x"17",
         10280 => x"33",
         10281 => x"86",
         10282 => x"84",
         10283 => x"85",
         10284 => x"81",
         10285 => x"18",
         10286 => x"75",
         10287 => x"1f",
         10288 => x"71",
         10289 => x"5d",
         10290 => x"7b",
         10291 => x"2e",
         10292 => x"a8",
         10293 => x"b8",
         10294 => x"58",
         10295 => x"2e",
         10296 => x"75",
         10297 => x"70",
         10298 => x"25",
         10299 => x"42",
         10300 => x"38",
         10301 => x"2e",
         10302 => x"58",
         10303 => x"06",
         10304 => x"84",
         10305 => x"33",
         10306 => x"78",
         10307 => x"06",
         10308 => x"58",
         10309 => x"f8",
         10310 => x"80",
         10311 => x"38",
         10312 => x"1a",
         10313 => x"7a",
         10314 => x"38",
         10315 => x"83",
         10316 => x"18",
         10317 => x"40",
         10318 => x"70",
         10319 => x"33",
         10320 => x"05",
         10321 => x"71",
         10322 => x"5b",
         10323 => x"77",
         10324 => x"c5",
         10325 => x"2e",
         10326 => x"0b",
         10327 => x"83",
         10328 => x"5d",
         10329 => x"81",
         10330 => x"7e",
         10331 => x"40",
         10332 => x"31",
         10333 => x"58",
         10334 => x"80",
         10335 => x"38",
         10336 => x"e1",
         10337 => x"fe",
         10338 => x"58",
         10339 => x"38",
         10340 => x"84",
         10341 => x"0d",
         10342 => x"75",
         10343 => x"dc",
         10344 => x"81",
         10345 => x"e6",
         10346 => x"58",
         10347 => x"8d",
         10348 => x"84",
         10349 => x"0d",
         10350 => x"80",
         10351 => x"e6",
         10352 => x"58",
         10353 => x"05",
         10354 => x"70",
         10355 => x"33",
         10356 => x"ff",
         10357 => x"5f",
         10358 => x"2e",
         10359 => x"74",
         10360 => x"38",
         10361 => x"8a",
         10362 => x"b8",
         10363 => x"78",
         10364 => x"5a",
         10365 => x"81",
         10366 => x"71",
         10367 => x"1b",
         10368 => x"40",
         10369 => x"84",
         10370 => x"80",
         10371 => x"93",
         10372 => x"5a",
         10373 => x"83",
         10374 => x"fd",
         10375 => x"e9",
         10376 => x"e8",
         10377 => x"88",
         10378 => x"55",
         10379 => x"09",
         10380 => x"d5",
         10381 => x"58",
         10382 => x"17",
         10383 => x"b1",
         10384 => x"33",
         10385 => x"2e",
         10386 => x"82",
         10387 => x"54",
         10388 => x"17",
         10389 => x"33",
         10390 => x"d2",
         10391 => x"84",
         10392 => x"85",
         10393 => x"81",
         10394 => x"18",
         10395 => x"99",
         10396 => x"18",
         10397 => x"17",
         10398 => x"18",
         10399 => x"2b",
         10400 => x"75",
         10401 => x"2e",
         10402 => x"f8",
         10403 => x"17",
         10404 => x"82",
         10405 => x"90",
         10406 => x"2b",
         10407 => x"33",
         10408 => x"88",
         10409 => x"71",
         10410 => x"59",
         10411 => x"59",
         10412 => x"85",
         10413 => x"09",
         10414 => x"cd",
         10415 => x"17",
         10416 => x"82",
         10417 => x"90",
         10418 => x"2b",
         10419 => x"33",
         10420 => x"88",
         10421 => x"71",
         10422 => x"40",
         10423 => x"5e",
         10424 => x"85",
         10425 => x"09",
         10426 => x"9d",
         10427 => x"17",
         10428 => x"82",
         10429 => x"90",
         10430 => x"2b",
         10431 => x"33",
         10432 => x"88",
         10433 => x"71",
         10434 => x"0c",
         10435 => x"1c",
         10436 => x"82",
         10437 => x"90",
         10438 => x"2b",
         10439 => x"33",
         10440 => x"88",
         10441 => x"71",
         10442 => x"05",
         10443 => x"49",
         10444 => x"40",
         10445 => x"5a",
         10446 => x"84",
         10447 => x"81",
         10448 => x"84",
         10449 => x"7c",
         10450 => x"84",
         10451 => x"8c",
         10452 => x"0b",
         10453 => x"f7",
         10454 => x"83",
         10455 => x"38",
         10456 => x"0c",
         10457 => x"39",
         10458 => x"17",
         10459 => x"17",
         10460 => x"18",
         10461 => x"ff",
         10462 => x"84",
         10463 => x"7a",
         10464 => x"06",
         10465 => x"84",
         10466 => x"83",
         10467 => x"17",
         10468 => x"08",
         10469 => x"a0",
         10470 => x"8b",
         10471 => x"33",
         10472 => x"2e",
         10473 => x"84",
         10474 => x"5a",
         10475 => x"74",
         10476 => x"2e",
         10477 => x"85",
         10478 => x"18",
         10479 => x"5c",
         10480 => x"ab",
         10481 => x"17",
         10482 => x"18",
         10483 => x"2b",
         10484 => x"8d",
         10485 => x"d2",
         10486 => x"22",
         10487 => x"ca",
         10488 => x"17",
         10489 => x"82",
         10490 => x"90",
         10491 => x"2b",
         10492 => x"33",
         10493 => x"88",
         10494 => x"71",
         10495 => x"0c",
         10496 => x"2b",
         10497 => x"40",
         10498 => x"d8",
         10499 => x"75",
         10500 => x"e8",
         10501 => x"f9",
         10502 => x"80",
         10503 => x"38",
         10504 => x"57",
         10505 => x"f7",
         10506 => x"5a",
         10507 => x"38",
         10508 => x"75",
         10509 => x"08",
         10510 => x"05",
         10511 => x"81",
         10512 => x"ff",
         10513 => x"fc",
         10514 => x"3d",
         10515 => x"d3",
         10516 => x"70",
         10517 => x"41",
         10518 => x"76",
         10519 => x"80",
         10520 => x"38",
         10521 => x"05",
         10522 => x"9f",
         10523 => x"74",
         10524 => x"e2",
         10525 => x"38",
         10526 => x"80",
         10527 => x"e2",
         10528 => x"80",
         10529 => x"c4",
         10530 => x"10",
         10531 => x"05",
         10532 => x"55",
         10533 => x"84",
         10534 => x"34",
         10535 => x"80",
         10536 => x"80",
         10537 => x"54",
         10538 => x"7c",
         10539 => x"2e",
         10540 => x"53",
         10541 => x"53",
         10542 => x"ef",
         10543 => x"bb",
         10544 => x"73",
         10545 => x"0c",
         10546 => x"04",
         10547 => x"bb",
         10548 => x"3d",
         10549 => x"33",
         10550 => x"81",
         10551 => x"56",
         10552 => x"26",
         10553 => x"16",
         10554 => x"06",
         10555 => x"58",
         10556 => x"80",
         10557 => x"7f",
         10558 => x"f4",
         10559 => x"7b",
         10560 => x"5a",
         10561 => x"05",
         10562 => x"70",
         10563 => x"33",
         10564 => x"59",
         10565 => x"99",
         10566 => x"e0",
         10567 => x"ff",
         10568 => x"ff",
         10569 => x"76",
         10570 => x"38",
         10571 => x"81",
         10572 => x"54",
         10573 => x"9f",
         10574 => x"74",
         10575 => x"81",
         10576 => x"76",
         10577 => x"77",
         10578 => x"30",
         10579 => x"9f",
         10580 => x"5c",
         10581 => x"80",
         10582 => x"81",
         10583 => x"5d",
         10584 => x"25",
         10585 => x"7f",
         10586 => x"39",
         10587 => x"f7",
         10588 => x"60",
         10589 => x"8b",
         10590 => x"0d",
         10591 => x"05",
         10592 => x"33",
         10593 => x"56",
         10594 => x"a6",
         10595 => x"06",
         10596 => x"3d",
         10597 => x"9e",
         10598 => x"52",
         10599 => x"3f",
         10600 => x"08",
         10601 => x"84",
         10602 => x"8f",
         10603 => x"0c",
         10604 => x"84",
         10605 => x"9c",
         10606 => x"7e",
         10607 => x"90",
         10608 => x"5c",
         10609 => x"84",
         10610 => x"57",
         10611 => x"08",
         10612 => x"ba",
         10613 => x"06",
         10614 => x"2e",
         10615 => x"76",
         10616 => x"e0",
         10617 => x"2e",
         10618 => x"78",
         10619 => x"76",
         10620 => x"78",
         10621 => x"06",
         10622 => x"2e",
         10623 => x"66",
         10624 => x"9a",
         10625 => x"88",
         10626 => x"70",
         10627 => x"5d",
         10628 => x"83",
         10629 => x"38",
         10630 => x"17",
         10631 => x"8f",
         10632 => x"0b",
         10633 => x"80",
         10634 => x"17",
         10635 => x"a0",
         10636 => x"34",
         10637 => x"5e",
         10638 => x"17",
         10639 => x"9b",
         10640 => x"33",
         10641 => x"2e",
         10642 => x"66",
         10643 => x"9c",
         10644 => x"0b",
         10645 => x"80",
         10646 => x"34",
         10647 => x"19",
         10648 => x"81",
         10649 => x"34",
         10650 => x"80",
         10651 => x"b4",
         10652 => x"7e",
         10653 => x"5f",
         10654 => x"27",
         10655 => x"16",
         10656 => x"83",
         10657 => x"57",
         10658 => x"fe",
         10659 => x"80",
         10660 => x"70",
         10661 => x"58",
         10662 => x"fe",
         10663 => x"79",
         10664 => x"57",
         10665 => x"38",
         10666 => x"38",
         10667 => x"05",
         10668 => x"2a",
         10669 => x"56",
         10670 => x"38",
         10671 => x"81",
         10672 => x"80",
         10673 => x"75",
         10674 => x"77",
         10675 => x"78",
         10676 => x"06",
         10677 => x"2e",
         10678 => x"80",
         10679 => x"7e",
         10680 => x"a0",
         10681 => x"a4",
         10682 => x"9b",
         10683 => x"12",
         10684 => x"2b",
         10685 => x"40",
         10686 => x"5b",
         10687 => x"81",
         10688 => x"88",
         10689 => x"16",
         10690 => x"82",
         10691 => x"90",
         10692 => x"2b",
         10693 => x"33",
         10694 => x"88",
         10695 => x"71",
         10696 => x"05",
         10697 => x"7f",
         10698 => x"5e",
         10699 => x"1b",
         10700 => x"23",
         10701 => x"34",
         10702 => x"1b",
         10703 => x"9c",
         10704 => x"0b",
         10705 => x"a8",
         10706 => x"80",
         10707 => x"80",
         10708 => x"05",
         10709 => x"15",
         10710 => x"38",
         10711 => x"81",
         10712 => x"80",
         10713 => x"38",
         10714 => x"55",
         10715 => x"fc",
         10716 => x"94",
         10717 => x"1b",
         10718 => x"2b",
         10719 => x"77",
         10720 => x"5b",
         10721 => x"78",
         10722 => x"51",
         10723 => x"27",
         10724 => x"81",
         10725 => x"5e",
         10726 => x"2e",
         10727 => x"77",
         10728 => x"ff",
         10729 => x"84",
         10730 => x"58",
         10731 => x"08",
         10732 => x"38",
         10733 => x"bb",
         10734 => x"2e",
         10735 => x"79",
         10736 => x"39",
         10737 => x"05",
         10738 => x"5e",
         10739 => x"78",
         10740 => x"06",
         10741 => x"2e",
         10742 => x"88",
         10743 => x"0c",
         10744 => x"87",
         10745 => x"0c",
         10746 => x"84",
         10747 => x"0c",
         10748 => x"7a",
         10749 => x"57",
         10750 => x"39",
         10751 => x"94",
         10752 => x"98",
         10753 => x"2b",
         10754 => x"88",
         10755 => x"18",
         10756 => x"82",
         10757 => x"90",
         10758 => x"2b",
         10759 => x"33",
         10760 => x"88",
         10761 => x"71",
         10762 => x"05",
         10763 => x"61",
         10764 => x"54",
         10765 => x"5c",
         10766 => x"84",
         10767 => x"90",
         10768 => x"0b",
         10769 => x"80",
         10770 => x"0c",
         10771 => x"1b",
         10772 => x"5c",
         10773 => x"57",
         10774 => x"39",
         10775 => x"c2",
         10776 => x"84",
         10777 => x"07",
         10778 => x"fa",
         10779 => x"83",
         10780 => x"7b",
         10781 => x"e9",
         10782 => x"84",
         10783 => x"bb",
         10784 => x"2e",
         10785 => x"84",
         10786 => x"81",
         10787 => x"38",
         10788 => x"08",
         10789 => x"b7",
         10790 => x"74",
         10791 => x"ff",
         10792 => x"84",
         10793 => x"83",
         10794 => x"16",
         10795 => x"94",
         10796 => x"56",
         10797 => x"27",
         10798 => x"17",
         10799 => x"84",
         10800 => x"07",
         10801 => x"17",
         10802 => x"77",
         10803 => x"a1",
         10804 => x"7f",
         10805 => x"57",
         10806 => x"08",
         10807 => x"38",
         10808 => x"58",
         10809 => x"09",
         10810 => x"eb",
         10811 => x"7d",
         10812 => x"52",
         10813 => x"51",
         10814 => x"3f",
         10815 => x"08",
         10816 => x"38",
         10817 => x"5c",
         10818 => x"0c",
         10819 => x"ff",
         10820 => x"0c",
         10821 => x"2e",
         10822 => x"80",
         10823 => x"90",
         10824 => x"94",
         10825 => x"0b",
         10826 => x"fa",
         10827 => x"16",
         10828 => x"33",
         10829 => x"71",
         10830 => x"7d",
         10831 => x"58",
         10832 => x"17",
         10833 => x"8f",
         10834 => x"0b",
         10835 => x"80",
         10836 => x"17",
         10837 => x"a0",
         10838 => x"34",
         10839 => x"5e",
         10840 => x"17",
         10841 => x"9b",
         10842 => x"33",
         10843 => x"2e",
         10844 => x"f9",
         10845 => x"a9",
         10846 => x"1b",
         10847 => x"ad",
         10848 => x"ff",
         10849 => x"80",
         10850 => x"38",
         10851 => x"9c",
         10852 => x"05",
         10853 => x"77",
         10854 => x"ea",
         10855 => x"22",
         10856 => x"b0",
         10857 => x"56",
         10858 => x"2e",
         10859 => x"75",
         10860 => x"70",
         10861 => x"58",
         10862 => x"53",
         10863 => x"19",
         10864 => x"a1",
         10865 => x"bb",
         10866 => x"2e",
         10867 => x"81",
         10868 => x"0c",
         10869 => x"81",
         10870 => x"08",
         10871 => x"70",
         10872 => x"33",
         10873 => x"a2",
         10874 => x"bb",
         10875 => x"2e",
         10876 => x"80",
         10877 => x"bb",
         10878 => x"17",
         10879 => x"08",
         10880 => x"31",
         10881 => x"08",
         10882 => x"a0",
         10883 => x"fd",
         10884 => x"16",
         10885 => x"82",
         10886 => x"06",
         10887 => x"81",
         10888 => x"08",
         10889 => x"05",
         10890 => x"81",
         10891 => x"ff",
         10892 => x"7c",
         10893 => x"39",
         10894 => x"08",
         10895 => x"0c",
         10896 => x"81",
         10897 => x"39",
         10898 => x"60",
         10899 => x"40",
         10900 => x"80",
         10901 => x"57",
         10902 => x"9f",
         10903 => x"56",
         10904 => x"97",
         10905 => x"55",
         10906 => x"8f",
         10907 => x"22",
         10908 => x"59",
         10909 => x"2e",
         10910 => x"80",
         10911 => x"76",
         10912 => x"e7",
         10913 => x"33",
         10914 => x"df",
         10915 => x"33",
         10916 => x"87",
         10917 => x"2e",
         10918 => x"94",
         10919 => x"1a",
         10920 => x"56",
         10921 => x"26",
         10922 => x"79",
         10923 => x"b0",
         10924 => x"ff",
         10925 => x"82",
         10926 => x"8a",
         10927 => x"05",
         10928 => x"06",
         10929 => x"9b",
         10930 => x"d0",
         10931 => x"08",
         10932 => x"27",
         10933 => x"74",
         10934 => x"ae",
         10935 => x"1a",
         10936 => x"98",
         10937 => x"05",
         10938 => x"fe",
         10939 => x"76",
         10940 => x"a5",
         10941 => x"22",
         10942 => x"b0",
         10943 => x"56",
         10944 => x"2e",
         10945 => x"7b",
         10946 => x"2a",
         10947 => x"80",
         10948 => x"38",
         10949 => x"75",
         10950 => x"38",
         10951 => x"5b",
         10952 => x"53",
         10953 => x"18",
         10954 => x"9f",
         10955 => x"bb",
         10956 => x"d6",
         10957 => x"33",
         10958 => x"59",
         10959 => x"24",
         10960 => x"7a",
         10961 => x"79",
         10962 => x"08",
         10963 => x"77",
         10964 => x"08",
         10965 => x"94",
         10966 => x"5a",
         10967 => x"38",
         10968 => x"84",
         10969 => x"90",
         10970 => x"74",
         10971 => x"0c",
         10972 => x"04",
         10973 => x"b3",
         10974 => x"08",
         10975 => x"2e",
         10976 => x"90",
         10977 => x"98",
         10978 => x"52",
         10979 => x"80",
         10980 => x"81",
         10981 => x"7a",
         10982 => x"33",
         10983 => x"8d",
         10984 => x"84",
         10985 => x"38",
         10986 => x"80",
         10987 => x"74",
         10988 => x"7e",
         10989 => x"76",
         10990 => x"81",
         10991 => x"ff",
         10992 => x"84",
         10993 => x"81",
         10994 => x"9c",
         10995 => x"19",
         10996 => x"83",
         10997 => x"80",
         10998 => x"55",
         10999 => x"83",
         11000 => x"76",
         11001 => x"a8",
         11002 => x"56",
         11003 => x"fe",
         11004 => x"70",
         11005 => x"33",
         11006 => x"05",
         11007 => x"16",
         11008 => x"2e",
         11009 => x"74",
         11010 => x"56",
         11011 => x"81",
         11012 => x"ff",
         11013 => x"da",
         11014 => x"39",
         11015 => x"52",
         11016 => x"a3",
         11017 => x"bb",
         11018 => x"fd",
         11019 => x"16",
         11020 => x"9c",
         11021 => x"bb",
         11022 => x"06",
         11023 => x"bb",
         11024 => x"08",
         11025 => x"b5",
         11026 => x"08",
         11027 => x"75",
         11028 => x"ef",
         11029 => x"76",
         11030 => x"a8",
         11031 => x"55",
         11032 => x"05",
         11033 => x"70",
         11034 => x"34",
         11035 => x"74",
         11036 => x"cf",
         11037 => x"81",
         11038 => x"77",
         11039 => x"59",
         11040 => x"55",
         11041 => x"fd",
         11042 => x"0b",
         11043 => x"81",
         11044 => x"84",
         11045 => x"0d",
         11046 => x"91",
         11047 => x"0b",
         11048 => x"0c",
         11049 => x"04",
         11050 => x"61",
         11051 => x"41",
         11052 => x"80",
         11053 => x"57",
         11054 => x"9f",
         11055 => x"56",
         11056 => x"97",
         11057 => x"55",
         11058 => x"8f",
         11059 => x"22",
         11060 => x"59",
         11061 => x"2e",
         11062 => x"80",
         11063 => x"76",
         11064 => x"cc",
         11065 => x"33",
         11066 => x"c4",
         11067 => x"33",
         11068 => x"81",
         11069 => x"87",
         11070 => x"2e",
         11071 => x"94",
         11072 => x"11",
         11073 => x"77",
         11074 => x"76",
         11075 => x"80",
         11076 => x"38",
         11077 => x"06",
         11078 => x"cd",
         11079 => x"11",
         11080 => x"78",
         11081 => x"5e",
         11082 => x"38",
         11083 => x"38",
         11084 => x"55",
         11085 => x"83",
         11086 => x"81",
         11087 => x"38",
         11088 => x"83",
         11089 => x"98",
         11090 => x"19",
         11091 => x"74",
         11092 => x"7f",
         11093 => x"33",
         11094 => x"5b",
         11095 => x"24",
         11096 => x"98",
         11097 => x"05",
         11098 => x"fe",
         11099 => x"76",
         11100 => x"b8",
         11101 => x"22",
         11102 => x"b0",
         11103 => x"56",
         11104 => x"2e",
         11105 => x"7c",
         11106 => x"2a",
         11107 => x"80",
         11108 => x"38",
         11109 => x"75",
         11110 => x"38",
         11111 => x"5a",
         11112 => x"53",
         11113 => x"18",
         11114 => x"9b",
         11115 => x"bb",
         11116 => x"e9",
         11117 => x"08",
         11118 => x"75",
         11119 => x"38",
         11120 => x"a8",
         11121 => x"29",
         11122 => x"58",
         11123 => x"81",
         11124 => x"77",
         11125 => x"59",
         11126 => x"55",
         11127 => x"90",
         11128 => x"ff",
         11129 => x"90",
         11130 => x"89",
         11131 => x"78",
         11132 => x"19",
         11133 => x"1f",
         11134 => x"1a",
         11135 => x"1e",
         11136 => x"08",
         11137 => x"5f",
         11138 => x"27",
         11139 => x"55",
         11140 => x"0c",
         11141 => x"38",
         11142 => x"58",
         11143 => x"07",
         11144 => x"1a",
         11145 => x"75",
         11146 => x"0c",
         11147 => x"04",
         11148 => x"84",
         11149 => x"0d",
         11150 => x"08",
         11151 => x"38",
         11152 => x"57",
         11153 => x"08",
         11154 => x"81",
         11155 => x"a8",
         11156 => x"18",
         11157 => x"98",
         11158 => x"bb",
         11159 => x"bd",
         11160 => x"08",
         11161 => x"1a",
         11162 => x"ff",
         11163 => x"71",
         11164 => x"7a",
         11165 => x"38",
         11166 => x"79",
         11167 => x"7f",
         11168 => x"77",
         11169 => x"38",
         11170 => x"05",
         11171 => x"70",
         11172 => x"34",
         11173 => x"75",
         11174 => x"19",
         11175 => x"07",
         11176 => x"1a",
         11177 => x"39",
         11178 => x"52",
         11179 => x"ac",
         11180 => x"bb",
         11181 => x"84",
         11182 => x"fc",
         11183 => x"19",
         11184 => x"d8",
         11185 => x"78",
         11186 => x"d4",
         11187 => x"84",
         11188 => x"bb",
         11189 => x"e2",
         11190 => x"81",
         11191 => x"08",
         11192 => x"52",
         11193 => x"51",
         11194 => x"3f",
         11195 => x"08",
         11196 => x"19",
         11197 => x"06",
         11198 => x"1a",
         11199 => x"fc",
         11200 => x"16",
         11201 => x"96",
         11202 => x"bb",
         11203 => x"06",
         11204 => x"c7",
         11205 => x"08",
         11206 => x"c1",
         11207 => x"91",
         11208 => x"0b",
         11209 => x"0c",
         11210 => x"04",
         11211 => x"1a",
         11212 => x"84",
         11213 => x"91",
         11214 => x"f5",
         11215 => x"58",
         11216 => x"80",
         11217 => x"77",
         11218 => x"80",
         11219 => x"75",
         11220 => x"80",
         11221 => x"86",
         11222 => x"19",
         11223 => x"79",
         11224 => x"d2",
         11225 => x"74",
         11226 => x"76",
         11227 => x"90",
         11228 => x"86",
         11229 => x"5c",
         11230 => x"2e",
         11231 => x"76",
         11232 => x"80",
         11233 => x"c9",
         11234 => x"19",
         11235 => x"b4",
         11236 => x"2e",
         11237 => x"0b",
         11238 => x"71",
         11239 => x"7a",
         11240 => x"81",
         11241 => x"38",
         11242 => x"53",
         11243 => x"81",
         11244 => x"ff",
         11245 => x"84",
         11246 => x"80",
         11247 => x"ff",
         11248 => x"76",
         11249 => x"78",
         11250 => x"90",
         11251 => x"08",
         11252 => x"a0",
         11253 => x"74",
         11254 => x"77",
         11255 => x"08",
         11256 => x"ff",
         11257 => x"56",
         11258 => x"34",
         11259 => x"5a",
         11260 => x"34",
         11261 => x"33",
         11262 => x"56",
         11263 => x"2e",
         11264 => x"8c",
         11265 => x"74",
         11266 => x"88",
         11267 => x"9d",
         11268 => x"90",
         11269 => x"9e",
         11270 => x"98",
         11271 => x"9f",
         11272 => x"7a",
         11273 => x"97",
         11274 => x"0b",
         11275 => x"80",
         11276 => x"18",
         11277 => x"92",
         11278 => x"0b",
         11279 => x"7b",
         11280 => x"83",
         11281 => x"51",
         11282 => x"3f",
         11283 => x"08",
         11284 => x"81",
         11285 => x"56",
         11286 => x"34",
         11287 => x"84",
         11288 => x"8d",
         11289 => x"81",
         11290 => x"08",
         11291 => x"70",
         11292 => x"33",
         11293 => x"95",
         11294 => x"59",
         11295 => x"08",
         11296 => x"81",
         11297 => x"38",
         11298 => x"08",
         11299 => x"b4",
         11300 => x"17",
         11301 => x"bb",
         11302 => x"55",
         11303 => x"08",
         11304 => x"38",
         11305 => x"55",
         11306 => x"09",
         11307 => x"f8",
         11308 => x"b4",
         11309 => x"17",
         11310 => x"7a",
         11311 => x"33",
         11312 => x"e9",
         11313 => x"fd",
         11314 => x"90",
         11315 => x"94",
         11316 => x"88",
         11317 => x"95",
         11318 => x"18",
         11319 => x"7b",
         11320 => x"2a",
         11321 => x"18",
         11322 => x"2a",
         11323 => x"18",
         11324 => x"2a",
         11325 => x"18",
         11326 => x"34",
         11327 => x"18",
         11328 => x"98",
         11329 => x"cc",
         11330 => x"34",
         11331 => x"18",
         11332 => x"93",
         11333 => x"5b",
         11334 => x"1c",
         11335 => x"ff",
         11336 => x"84",
         11337 => x"90",
         11338 => x"bf",
         11339 => x"79",
         11340 => x"fe",
         11341 => x"16",
         11342 => x"92",
         11343 => x"bb",
         11344 => x"06",
         11345 => x"9d",
         11346 => x"08",
         11347 => x"97",
         11348 => x"9c",
         11349 => x"a8",
         11350 => x"81",
         11351 => x"57",
         11352 => x"3f",
         11353 => x"bb",
         11354 => x"f2",
         11355 => x"33",
         11356 => x"59",
         11357 => x"34",
         11358 => x"08",
         11359 => x"16",
         11360 => x"09",
         11361 => x"8e",
         11362 => x"39",
         11363 => x"79",
         11364 => x"fb",
         11365 => x"bb",
         11366 => x"84",
         11367 => x"b1",
         11368 => x"74",
         11369 => x"38",
         11370 => x"72",
         11371 => x"38",
         11372 => x"71",
         11373 => x"38",
         11374 => x"84",
         11375 => x"52",
         11376 => x"96",
         11377 => x"71",
         11378 => x"75",
         11379 => x"75",
         11380 => x"bb",
         11381 => x"3d",
         11382 => x"13",
         11383 => x"90",
         11384 => x"bb",
         11385 => x"06",
         11386 => x"38",
         11387 => x"53",
         11388 => x"f6",
         11389 => x"7d",
         11390 => x"5b",
         11391 => x"b2",
         11392 => x"81",
         11393 => x"70",
         11394 => x"52",
         11395 => x"ac",
         11396 => x"38",
         11397 => x"a4",
         11398 => x"e0",
         11399 => x"71",
         11400 => x"70",
         11401 => x"34",
         11402 => x"bb",
         11403 => x"3d",
         11404 => x"0b",
         11405 => x"0c",
         11406 => x"04",
         11407 => x"11",
         11408 => x"06",
         11409 => x"70",
         11410 => x"38",
         11411 => x"81",
         11412 => x"05",
         11413 => x"76",
         11414 => x"38",
         11415 => x"e6",
         11416 => x"79",
         11417 => x"57",
         11418 => x"05",
         11419 => x"70",
         11420 => x"33",
         11421 => x"53",
         11422 => x"99",
         11423 => x"e0",
         11424 => x"ff",
         11425 => x"ff",
         11426 => x"70",
         11427 => x"38",
         11428 => x"81",
         11429 => x"54",
         11430 => x"9f",
         11431 => x"71",
         11432 => x"81",
         11433 => x"73",
         11434 => x"74",
         11435 => x"30",
         11436 => x"9f",
         11437 => x"59",
         11438 => x"80",
         11439 => x"81",
         11440 => x"5b",
         11441 => x"25",
         11442 => x"7a",
         11443 => x"39",
         11444 => x"f7",
         11445 => x"5e",
         11446 => x"39",
         11447 => x"80",
         11448 => x"cc",
         11449 => x"3d",
         11450 => x"3f",
         11451 => x"08",
         11452 => x"84",
         11453 => x"8a",
         11454 => x"bb",
         11455 => x"3d",
         11456 => x"5c",
         11457 => x"3d",
         11458 => x"c6",
         11459 => x"bb",
         11460 => x"84",
         11461 => x"80",
         11462 => x"80",
         11463 => x"70",
         11464 => x"5a",
         11465 => x"80",
         11466 => x"b2",
         11467 => x"84",
         11468 => x"57",
         11469 => x"2e",
         11470 => x"63",
         11471 => x"9a",
         11472 => x"88",
         11473 => x"33",
         11474 => x"57",
         11475 => x"2e",
         11476 => x"98",
         11477 => x"84",
         11478 => x"98",
         11479 => x"84",
         11480 => x"84",
         11481 => x"06",
         11482 => x"85",
         11483 => x"84",
         11484 => x"0d",
         11485 => x"33",
         11486 => x"71",
         11487 => x"90",
         11488 => x"07",
         11489 => x"5b",
         11490 => x"7a",
         11491 => x"0c",
         11492 => x"bb",
         11493 => x"3d",
         11494 => x"9e",
         11495 => x"e6",
         11496 => x"e6",
         11497 => x"40",
         11498 => x"80",
         11499 => x"3d",
         11500 => x"52",
         11501 => x"51",
         11502 => x"84",
         11503 => x"59",
         11504 => x"08",
         11505 => x"60",
         11506 => x"0c",
         11507 => x"11",
         11508 => x"3d",
         11509 => x"db",
         11510 => x"58",
         11511 => x"82",
         11512 => x"d8",
         11513 => x"40",
         11514 => x"7a",
         11515 => x"e9",
         11516 => x"84",
         11517 => x"bb",
         11518 => x"92",
         11519 => x"df",
         11520 => x"56",
         11521 => x"77",
         11522 => x"84",
         11523 => x"83",
         11524 => x"5d",
         11525 => x"38",
         11526 => x"53",
         11527 => x"81",
         11528 => x"ff",
         11529 => x"84",
         11530 => x"80",
         11531 => x"ff",
         11532 => x"76",
         11533 => x"78",
         11534 => x"80",
         11535 => x"9b",
         11536 => x"12",
         11537 => x"2b",
         11538 => x"33",
         11539 => x"56",
         11540 => x"2e",
         11541 => x"76",
         11542 => x"0c",
         11543 => x"51",
         11544 => x"3f",
         11545 => x"08",
         11546 => x"84",
         11547 => x"38",
         11548 => x"51",
         11549 => x"3f",
         11550 => x"08",
         11551 => x"84",
         11552 => x"80",
         11553 => x"9b",
         11554 => x"12",
         11555 => x"2b",
         11556 => x"33",
         11557 => x"5e",
         11558 => x"2e",
         11559 => x"76",
         11560 => x"38",
         11561 => x"08",
         11562 => x"ff",
         11563 => x"84",
         11564 => x"59",
         11565 => x"08",
         11566 => x"b4",
         11567 => x"2e",
         11568 => x"78",
         11569 => x"80",
         11570 => x"b8",
         11571 => x"51",
         11572 => x"3f",
         11573 => x"05",
         11574 => x"79",
         11575 => x"38",
         11576 => x"81",
         11577 => x"70",
         11578 => x"57",
         11579 => x"81",
         11580 => x"78",
         11581 => x"38",
         11582 => x"9c",
         11583 => x"82",
         11584 => x"18",
         11585 => x"08",
         11586 => x"ff",
         11587 => x"56",
         11588 => x"75",
         11589 => x"38",
         11590 => x"e6",
         11591 => x"5f",
         11592 => x"34",
         11593 => x"08",
         11594 => x"bd",
         11595 => x"2e",
         11596 => x"80",
         11597 => x"e0",
         11598 => x"10",
         11599 => x"05",
         11600 => x"33",
         11601 => x"5e",
         11602 => x"2e",
         11603 => x"1a",
         11604 => x"33",
         11605 => x"74",
         11606 => x"1a",
         11607 => x"26",
         11608 => x"57",
         11609 => x"94",
         11610 => x"5f",
         11611 => x"70",
         11612 => x"34",
         11613 => x"79",
         11614 => x"38",
         11615 => x"81",
         11616 => x"76",
         11617 => x"81",
         11618 => x"38",
         11619 => x"7c",
         11620 => x"bb",
         11621 => x"e4",
         11622 => x"95",
         11623 => x"17",
         11624 => x"2b",
         11625 => x"07",
         11626 => x"56",
         11627 => x"39",
         11628 => x"94",
         11629 => x"98",
         11630 => x"2b",
         11631 => x"80",
         11632 => x"5a",
         11633 => x"7a",
         11634 => x"8d",
         11635 => x"84",
         11636 => x"bb",
         11637 => x"2e",
         11638 => x"ff",
         11639 => x"54",
         11640 => x"53",
         11641 => x"53",
         11642 => x"52",
         11643 => x"bd",
         11644 => x"84",
         11645 => x"fc",
         11646 => x"bb",
         11647 => x"17",
         11648 => x"08",
         11649 => x"31",
         11650 => x"08",
         11651 => x"a0",
         11652 => x"fc",
         11653 => x"16",
         11654 => x"82",
         11655 => x"06",
         11656 => x"81",
         11657 => x"08",
         11658 => x"05",
         11659 => x"81",
         11660 => x"ff",
         11661 => x"7c",
         11662 => x"39",
         11663 => x"e6",
         11664 => x"5c",
         11665 => x"34",
         11666 => x"e2",
         11667 => x"10",
         11668 => x"f4",
         11669 => x"70",
         11670 => x"59",
         11671 => x"7a",
         11672 => x"06",
         11673 => x"fd",
         11674 => x"e5",
         11675 => x"81",
         11676 => x"79",
         11677 => x"81",
         11678 => x"77",
         11679 => x"8e",
         11680 => x"3d",
         11681 => x"19",
         11682 => x"33",
         11683 => x"05",
         11684 => x"78",
         11685 => x"fd",
         11686 => x"59",
         11687 => x"78",
         11688 => x"0c",
         11689 => x"0d",
         11690 => x"0d",
         11691 => x"57",
         11692 => x"80",
         11693 => x"76",
         11694 => x"80",
         11695 => x"75",
         11696 => x"80",
         11697 => x"86",
         11698 => x"18",
         11699 => x"7a",
         11700 => x"ee",
         11701 => x"74",
         11702 => x"77",
         11703 => x"91",
         11704 => x"74",
         11705 => x"8c",
         11706 => x"78",
         11707 => x"f2",
         11708 => x"08",
         11709 => x"78",
         11710 => x"85",
         11711 => x"11",
         11712 => x"2b",
         11713 => x"75",
         11714 => x"fc",
         11715 => x"ff",
         11716 => x"bb",
         11717 => x"bb",
         11718 => x"17",
         11719 => x"53",
         11720 => x"bb",
         11721 => x"bb",
         11722 => x"26",
         11723 => x"77",
         11724 => x"70",
         11725 => x"79",
         11726 => x"19",
         11727 => x"5b",
         11728 => x"81",
         11729 => x"79",
         11730 => x"38",
         11731 => x"94",
         11732 => x"94",
         11733 => x"18",
         11734 => x"2a",
         11735 => x"5c",
         11736 => x"2e",
         11737 => x"75",
         11738 => x"ff",
         11739 => x"84",
         11740 => x"56",
         11741 => x"08",
         11742 => x"38",
         11743 => x"81",
         11744 => x"76",
         11745 => x"38",
         11746 => x"9c",
         11747 => x"82",
         11748 => x"98",
         11749 => x"ae",
         11750 => x"84",
         11751 => x"17",
         11752 => x"18",
         11753 => x"ff",
         11754 => x"80",
         11755 => x"7b",
         11756 => x"12",
         11757 => x"5c",
         11758 => x"7a",
         11759 => x"38",
         11760 => x"76",
         11761 => x"1a",
         11762 => x"89",
         11763 => x"5c",
         11764 => x"2e",
         11765 => x"8c",
         11766 => x"94",
         11767 => x"77",
         11768 => x"38",
         11769 => x"0c",
         11770 => x"80",
         11771 => x"78",
         11772 => x"75",
         11773 => x"5b",
         11774 => x"81",
         11775 => x"17",
         11776 => x"7a",
         11777 => x"38",
         11778 => x"70",
         11779 => x"19",
         11780 => x"74",
         11781 => x"38",
         11782 => x"53",
         11783 => x"81",
         11784 => x"56",
         11785 => x"3f",
         11786 => x"08",
         11787 => x"17",
         11788 => x"06",
         11789 => x"18",
         11790 => x"79",
         11791 => x"7b",
         11792 => x"52",
         11793 => x"e6",
         11794 => x"84",
         11795 => x"80",
         11796 => x"0b",
         11797 => x"81",
         11798 => x"bb",
         11799 => x"3d",
         11800 => x"17",
         11801 => x"2a",
         11802 => x"5a",
         11803 => x"38",
         11804 => x"08",
         11805 => x"5a",
         11806 => x"09",
         11807 => x"fd",
         11808 => x"18",
         11809 => x"39",
         11810 => x"18",
         11811 => x"08",
         11812 => x"2e",
         11813 => x"75",
         11814 => x"75",
         11815 => x"b7",
         11816 => x"39",
         11817 => x"0c",
         11818 => x"bb",
         11819 => x"3d",
         11820 => x"52",
         11821 => x"8a",
         11822 => x"bb",
         11823 => x"fd",
         11824 => x"16",
         11825 => x"83",
         11826 => x"bb",
         11827 => x"06",
         11828 => x"81",
         11829 => x"08",
         11830 => x"fb",
         11831 => x"76",
         11832 => x"bc",
         11833 => x"84",
         11834 => x"bb",
         11835 => x"2e",
         11836 => x"bb",
         11837 => x"2e",
         11838 => x"84",
         11839 => x"88",
         11840 => x"98",
         11841 => x"93",
         11842 => x"91",
         11843 => x"0b",
         11844 => x"0c",
         11845 => x"04",
         11846 => x"7c",
         11847 => x"75",
         11848 => x"38",
         11849 => x"3d",
         11850 => x"8d",
         11851 => x"51",
         11852 => x"84",
         11853 => x"55",
         11854 => x"08",
         11855 => x"38",
         11856 => x"74",
         11857 => x"bb",
         11858 => x"3d",
         11859 => x"76",
         11860 => x"75",
         11861 => x"88",
         11862 => x"84",
         11863 => x"bb",
         11864 => x"d1",
         11865 => x"33",
         11866 => x"59",
         11867 => x"24",
         11868 => x"16",
         11869 => x"2a",
         11870 => x"54",
         11871 => x"80",
         11872 => x"16",
         11873 => x"33",
         11874 => x"71",
         11875 => x"7d",
         11876 => x"5d",
         11877 => x"78",
         11878 => x"38",
         11879 => x"0c",
         11880 => x"18",
         11881 => x"23",
         11882 => x"51",
         11883 => x"3f",
         11884 => x"08",
         11885 => x"2e",
         11886 => x"80",
         11887 => x"38",
         11888 => x"fe",
         11889 => x"55",
         11890 => x"fe",
         11891 => x"17",
         11892 => x"33",
         11893 => x"71",
         11894 => x"7a",
         11895 => x"0c",
         11896 => x"bc",
         11897 => x"0d",
         11898 => x"54",
         11899 => x"9e",
         11900 => x"53",
         11901 => x"96",
         11902 => x"52",
         11903 => x"8e",
         11904 => x"22",
         11905 => x"57",
         11906 => x"2e",
         11907 => x"52",
         11908 => x"84",
         11909 => x"0c",
         11910 => x"84",
         11911 => x"0d",
         11912 => x"33",
         11913 => x"b4",
         11914 => x"84",
         11915 => x"52",
         11916 => x"71",
         11917 => x"54",
         11918 => x"3d",
         11919 => x"58",
         11920 => x"74",
         11921 => x"38",
         11922 => x"73",
         11923 => x"38",
         11924 => x"72",
         11925 => x"38",
         11926 => x"84",
         11927 => x"53",
         11928 => x"81",
         11929 => x"53",
         11930 => x"53",
         11931 => x"38",
         11932 => x"80",
         11933 => x"52",
         11934 => x"9e",
         11935 => x"bb",
         11936 => x"84",
         11937 => x"84",
         11938 => x"84",
         11939 => x"a6",
         11940 => x"74",
         11941 => x"83",
         11942 => x"74",
         11943 => x"af",
         11944 => x"84",
         11945 => x"70",
         11946 => x"07",
         11947 => x"bb",
         11948 => x"55",
         11949 => x"84",
         11950 => x"8a",
         11951 => x"75",
         11952 => x"52",
         11953 => x"d3",
         11954 => x"74",
         11955 => x"ff",
         11956 => x"84",
         11957 => x"70",
         11958 => x"07",
         11959 => x"bb",
         11960 => x"55",
         11961 => x"39",
         11962 => x"51",
         11963 => x"3f",
         11964 => x"08",
         11965 => x"0c",
         11966 => x"04",
         11967 => x"51",
         11968 => x"3f",
         11969 => x"08",
         11970 => x"72",
         11971 => x"72",
         11972 => x"56",
         11973 => x"ed",
         11974 => x"57",
         11975 => x"3d",
         11976 => x"3d",
         11977 => x"96",
         11978 => x"84",
         11979 => x"bb",
         11980 => x"2e",
         11981 => x"84",
         11982 => x"95",
         11983 => x"65",
         11984 => x"ff",
         11985 => x"84",
         11986 => x"55",
         11987 => x"08",
         11988 => x"80",
         11989 => x"70",
         11990 => x"58",
         11991 => x"97",
         11992 => x"2e",
         11993 => x"52",
         11994 => x"b1",
         11995 => x"84",
         11996 => x"95",
         11997 => x"86",
         11998 => x"84",
         11999 => x"0d",
         12000 => x"0d",
         12001 => x"5f",
         12002 => x"3d",
         12003 => x"96",
         12004 => x"aa",
         12005 => x"84",
         12006 => x"bb",
         12007 => x"38",
         12008 => x"74",
         12009 => x"08",
         12010 => x"13",
         12011 => x"59",
         12012 => x"26",
         12013 => x"7f",
         12014 => x"bb",
         12015 => x"3d",
         12016 => x"bb",
         12017 => x"33",
         12018 => x"81",
         12019 => x"38",
         12020 => x"08",
         12021 => x"08",
         12022 => x"77",
         12023 => x"7b",
         12024 => x"5c",
         12025 => x"17",
         12026 => x"82",
         12027 => x"17",
         12028 => x"5d",
         12029 => x"38",
         12030 => x"53",
         12031 => x"81",
         12032 => x"fe",
         12033 => x"84",
         12034 => x"80",
         12035 => x"ff",
         12036 => x"79",
         12037 => x"7f",
         12038 => x"7d",
         12039 => x"76",
         12040 => x"82",
         12041 => x"38",
         12042 => x"05",
         12043 => x"82",
         12044 => x"90",
         12045 => x"2b",
         12046 => x"33",
         12047 => x"88",
         12048 => x"71",
         12049 => x"fe",
         12050 => x"70",
         12051 => x"25",
         12052 => x"84",
         12053 => x"06",
         12054 => x"43",
         12055 => x"54",
         12056 => x"40",
         12057 => x"fe",
         12058 => x"7f",
         12059 => x"18",
         12060 => x"33",
         12061 => x"77",
         12062 => x"79",
         12063 => x"0c",
         12064 => x"04",
         12065 => x"17",
         12066 => x"17",
         12067 => x"18",
         12068 => x"fe",
         12069 => x"81",
         12070 => x"84",
         12071 => x"38",
         12072 => x"08",
         12073 => x"b4",
         12074 => x"18",
         12075 => x"bb",
         12076 => x"55",
         12077 => x"08",
         12078 => x"38",
         12079 => x"55",
         12080 => x"09",
         12081 => x"b0",
         12082 => x"b4",
         12083 => x"18",
         12084 => x"7c",
         12085 => x"33",
         12086 => x"d1",
         12087 => x"fe",
         12088 => x"77",
         12089 => x"59",
         12090 => x"77",
         12091 => x"f1",
         12092 => x"84",
         12093 => x"80",
         12094 => x"bb",
         12095 => x"2e",
         12096 => x"84",
         12097 => x"30",
         12098 => x"84",
         12099 => x"25",
         12100 => x"18",
         12101 => x"5c",
         12102 => x"08",
         12103 => x"38",
         12104 => x"7a",
         12105 => x"84",
         12106 => x"07",
         12107 => x"18",
         12108 => x"39",
         12109 => x"05",
         12110 => x"71",
         12111 => x"2b",
         12112 => x"70",
         12113 => x"82",
         12114 => x"06",
         12115 => x"5d",
         12116 => x"5f",
         12117 => x"83",
         12118 => x"39",
         12119 => x"bf",
         12120 => x"58",
         12121 => x"0c",
         12122 => x"0c",
         12123 => x"81",
         12124 => x"84",
         12125 => x"83",
         12126 => x"58",
         12127 => x"f6",
         12128 => x"58",
         12129 => x"80",
         12130 => x"77",
         12131 => x"80",
         12132 => x"75",
         12133 => x"80",
         12134 => x"86",
         12135 => x"19",
         12136 => x"79",
         12137 => x"81",
         12138 => x"74",
         12139 => x"83",
         12140 => x"33",
         12141 => x"fb",
         12142 => x"33",
         12143 => x"81",
         12144 => x"87",
         12145 => x"2e",
         12146 => x"94",
         12147 => x"74",
         12148 => x"27",
         12149 => x"74",
         12150 => x"88",
         12151 => x"08",
         12152 => x"75",
         12153 => x"9c",
         12154 => x"26",
         12155 => x"82",
         12156 => x"88",
         12157 => x"18",
         12158 => x"0c",
         12159 => x"07",
         12160 => x"19",
         12161 => x"38",
         12162 => x"5a",
         12163 => x"a3",
         12164 => x"9c",
         12165 => x"a8",
         12166 => x"81",
         12167 => x"59",
         12168 => x"3f",
         12169 => x"08",
         12170 => x"90",
         12171 => x"76",
         12172 => x"76",
         12173 => x"bb",
         12174 => x"3d",
         12175 => x"55",
         12176 => x"80",
         12177 => x"52",
         12178 => x"ff",
         12179 => x"bb",
         12180 => x"84",
         12181 => x"80",
         12182 => x"38",
         12183 => x"08",
         12184 => x"e8",
         12185 => x"84",
         12186 => x"82",
         12187 => x"53",
         12188 => x"51",
         12189 => x"3f",
         12190 => x"08",
         12191 => x"9c",
         12192 => x"11",
         12193 => x"58",
         12194 => x"75",
         12195 => x"38",
         12196 => x"18",
         12197 => x"33",
         12198 => x"74",
         12199 => x"79",
         12200 => x"26",
         12201 => x"9c",
         12202 => x"33",
         12203 => x"ac",
         12204 => x"84",
         12205 => x"55",
         12206 => x"38",
         12207 => x"56",
         12208 => x"39",
         12209 => x"19",
         12210 => x"74",
         12211 => x"88",
         12212 => x"a2",
         12213 => x"08",
         12214 => x"fe",
         12215 => x"84",
         12216 => x"ff",
         12217 => x"38",
         12218 => x"08",
         12219 => x"be",
         12220 => x"ae",
         12221 => x"84",
         12222 => x"9c",
         12223 => x"81",
         12224 => x"bb",
         12225 => x"19",
         12226 => x"59",
         12227 => x"0b",
         12228 => x"08",
         12229 => x"38",
         12230 => x"08",
         12231 => x"27",
         12232 => x"75",
         12233 => x"38",
         12234 => x"52",
         12235 => x"84",
         12236 => x"bb",
         12237 => x"84",
         12238 => x"80",
         12239 => x"52",
         12240 => x"fd",
         12241 => x"bb",
         12242 => x"84",
         12243 => x"80",
         12244 => x"38",
         12245 => x"08",
         12246 => x"dc",
         12247 => x"84",
         12248 => x"81",
         12249 => x"53",
         12250 => x"51",
         12251 => x"3f",
         12252 => x"08",
         12253 => x"9c",
         12254 => x"11",
         12255 => x"58",
         12256 => x"75",
         12257 => x"81",
         12258 => x"0c",
         12259 => x"81",
         12260 => x"84",
         12261 => x"55",
         12262 => x"ff",
         12263 => x"56",
         12264 => x"18",
         12265 => x"ce",
         12266 => x"fe",
         12267 => x"0b",
         12268 => x"5a",
         12269 => x"39",
         12270 => x"39",
         12271 => x"80",
         12272 => x"74",
         12273 => x"76",
         12274 => x"39",
         12275 => x"19",
         12276 => x"fd",
         12277 => x"bb",
         12278 => x"19",
         12279 => x"fd",
         12280 => x"0b",
         12281 => x"5a",
         12282 => x"39",
         12283 => x"08",
         12284 => x"39",
         12285 => x"aa",
         12286 => x"0d",
         12287 => x"3d",
         12288 => x"52",
         12289 => x"ff",
         12290 => x"84",
         12291 => x"56",
         12292 => x"08",
         12293 => x"38",
         12294 => x"84",
         12295 => x"0d",
         12296 => x"a8",
         12297 => x"9b",
         12298 => x"59",
         12299 => x"3f",
         12300 => x"08",
         12301 => x"84",
         12302 => x"02",
         12303 => x"33",
         12304 => x"81",
         12305 => x"86",
         12306 => x"38",
         12307 => x"5b",
         12308 => x"c4",
         12309 => x"ee",
         12310 => x"81",
         12311 => x"87",
         12312 => x"b4",
         12313 => x"3d",
         12314 => x"33",
         12315 => x"71",
         12316 => x"73",
         12317 => x"5c",
         12318 => x"83",
         12319 => x"38",
         12320 => x"81",
         12321 => x"80",
         12322 => x"38",
         12323 => x"18",
         12324 => x"ff",
         12325 => x"5f",
         12326 => x"bb",
         12327 => x"8f",
         12328 => x"55",
         12329 => x"3f",
         12330 => x"08",
         12331 => x"84",
         12332 => x"38",
         12333 => x"08",
         12334 => x"ff",
         12335 => x"84",
         12336 => x"56",
         12337 => x"08",
         12338 => x"0b",
         12339 => x"0c",
         12340 => x"04",
         12341 => x"94",
         12342 => x"98",
         12343 => x"2b",
         12344 => x"5d",
         12345 => x"98",
         12346 => x"84",
         12347 => x"88",
         12348 => x"84",
         12349 => x"38",
         12350 => x"a8",
         12351 => x"5d",
         12352 => x"2e",
         12353 => x"74",
         12354 => x"ff",
         12355 => x"84",
         12356 => x"56",
         12357 => x"08",
         12358 => x"38",
         12359 => x"77",
         12360 => x"56",
         12361 => x"2e",
         12362 => x"80",
         12363 => x"7a",
         12364 => x"55",
         12365 => x"89",
         12366 => x"08",
         12367 => x"fd",
         12368 => x"75",
         12369 => x"7d",
         12370 => x"94",
         12371 => x"84",
         12372 => x"84",
         12373 => x"0d",
         12374 => x"5d",
         12375 => x"56",
         12376 => x"17",
         12377 => x"82",
         12378 => x"17",
         12379 => x"55",
         12380 => x"09",
         12381 => x"dd",
         12382 => x"75",
         12383 => x"52",
         12384 => x"51",
         12385 => x"3f",
         12386 => x"08",
         12387 => x"38",
         12388 => x"58",
         12389 => x"0c",
         12390 => x"ab",
         12391 => x"08",
         12392 => x"34",
         12393 => x"18",
         12394 => x"08",
         12395 => x"ec",
         12396 => x"78",
         12397 => x"97",
         12398 => x"84",
         12399 => x"bb",
         12400 => x"2e",
         12401 => x"75",
         12402 => x"81",
         12403 => x"38",
         12404 => x"c8",
         12405 => x"b4",
         12406 => x"7c",
         12407 => x"33",
         12408 => x"c9",
         12409 => x"84",
         12410 => x"7a",
         12411 => x"06",
         12412 => x"84",
         12413 => x"83",
         12414 => x"17",
         12415 => x"08",
         12416 => x"84",
         12417 => x"74",
         12418 => x"27",
         12419 => x"82",
         12420 => x"74",
         12421 => x"81",
         12422 => x"38",
         12423 => x"17",
         12424 => x"08",
         12425 => x"52",
         12426 => x"51",
         12427 => x"3f",
         12428 => x"c5",
         12429 => x"79",
         12430 => x"e1",
         12431 => x"78",
         12432 => x"9d",
         12433 => x"84",
         12434 => x"bb",
         12435 => x"2e",
         12436 => x"84",
         12437 => x"81",
         12438 => x"38",
         12439 => x"08",
         12440 => x"cb",
         12441 => x"74",
         12442 => x"fe",
         12443 => x"84",
         12444 => x"b3",
         12445 => x"08",
         12446 => x"19",
         12447 => x"58",
         12448 => x"ff",
         12449 => x"16",
         12450 => x"84",
         12451 => x"07",
         12452 => x"18",
         12453 => x"77",
         12454 => x"a1",
         12455 => x"fd",
         12456 => x"56",
         12457 => x"84",
         12458 => x"56",
         12459 => x"81",
         12460 => x"39",
         12461 => x"82",
         12462 => x"ff",
         12463 => x"a0",
         12464 => x"b2",
         12465 => x"bb",
         12466 => x"84",
         12467 => x"80",
         12468 => x"75",
         12469 => x"0c",
         12470 => x"04",
         12471 => x"52",
         12472 => x"52",
         12473 => x"f8",
         12474 => x"84",
         12475 => x"bb",
         12476 => x"38",
         12477 => x"bb",
         12478 => x"3d",
         12479 => x"bb",
         12480 => x"2e",
         12481 => x"cb",
         12482 => x"f3",
         12483 => x"85",
         12484 => x"56",
         12485 => x"74",
         12486 => x"7d",
         12487 => x"8f",
         12488 => x"5d",
         12489 => x"3f",
         12490 => x"08",
         12491 => x"84",
         12492 => x"83",
         12493 => x"84",
         12494 => x"81",
         12495 => x"38",
         12496 => x"08",
         12497 => x"cb",
         12498 => x"c9",
         12499 => x"bb",
         12500 => x"12",
         12501 => x"57",
         12502 => x"38",
         12503 => x"18",
         12504 => x"5a",
         12505 => x"75",
         12506 => x"38",
         12507 => x"76",
         12508 => x"19",
         12509 => x"58",
         12510 => x"0c",
         12511 => x"84",
         12512 => x"55",
         12513 => x"81",
         12514 => x"ff",
         12515 => x"f4",
         12516 => x"8a",
         12517 => x"77",
         12518 => x"f9",
         12519 => x"77",
         12520 => x"52",
         12521 => x"51",
         12522 => x"3f",
         12523 => x"08",
         12524 => x"81",
         12525 => x"39",
         12526 => x"84",
         12527 => x"b4",
         12528 => x"b8",
         12529 => x"81",
         12530 => x"58",
         12531 => x"3f",
         12532 => x"bb",
         12533 => x"38",
         12534 => x"08",
         12535 => x"b4",
         12536 => x"18",
         12537 => x"74",
         12538 => x"27",
         12539 => x"82",
         12540 => x"7a",
         12541 => x"81",
         12542 => x"38",
         12543 => x"17",
         12544 => x"08",
         12545 => x"52",
         12546 => x"51",
         12547 => x"3f",
         12548 => x"81",
         12549 => x"08",
         12550 => x"7c",
         12551 => x"38",
         12552 => x"08",
         12553 => x"38",
         12554 => x"51",
         12555 => x"3f",
         12556 => x"08",
         12557 => x"84",
         12558 => x"fd",
         12559 => x"bb",
         12560 => x"2e",
         12561 => x"84",
         12562 => x"ff",
         12563 => x"38",
         12564 => x"52",
         12565 => x"f9",
         12566 => x"bb",
         12567 => x"f3",
         12568 => x"08",
         12569 => x"19",
         12570 => x"59",
         12571 => x"90",
         12572 => x"94",
         12573 => x"17",
         12574 => x"5c",
         12575 => x"34",
         12576 => x"7a",
         12577 => x"38",
         12578 => x"84",
         12579 => x"0d",
         12580 => x"22",
         12581 => x"ff",
         12582 => x"81",
         12583 => x"2e",
         12584 => x"fe",
         12585 => x"0b",
         12586 => x"56",
         12587 => x"81",
         12588 => x"ff",
         12589 => x"f4",
         12590 => x"ae",
         12591 => x"34",
         12592 => x"0b",
         12593 => x"34",
         12594 => x"80",
         12595 => x"75",
         12596 => x"34",
         12597 => x"d0",
         12598 => x"cc",
         12599 => x"1a",
         12600 => x"83",
         12601 => x"59",
         12602 => x"d2",
         12603 => x"88",
         12604 => x"80",
         12605 => x"75",
         12606 => x"83",
         12607 => x"38",
         12608 => x"0b",
         12609 => x"b8",
         12610 => x"56",
         12611 => x"05",
         12612 => x"70",
         12613 => x"34",
         12614 => x"75",
         12615 => x"56",
         12616 => x"d9",
         12617 => x"7e",
         12618 => x"ff",
         12619 => x"57",
         12620 => x"17",
         12621 => x"2a",
         12622 => x"f3",
         12623 => x"33",
         12624 => x"2e",
         12625 => x"7d",
         12626 => x"83",
         12627 => x"51",
         12628 => x"3f",
         12629 => x"08",
         12630 => x"84",
         12631 => x"38",
         12632 => x"bb",
         12633 => x"17",
         12634 => x"84",
         12635 => x"34",
         12636 => x"17",
         12637 => x"0b",
         12638 => x"7d",
         12639 => x"77",
         12640 => x"77",
         12641 => x"78",
         12642 => x"7c",
         12643 => x"83",
         12644 => x"38",
         12645 => x"0b",
         12646 => x"7d",
         12647 => x"83",
         12648 => x"51",
         12649 => x"3f",
         12650 => x"08",
         12651 => x"bb",
         12652 => x"3d",
         12653 => x"90",
         12654 => x"80",
         12655 => x"74",
         12656 => x"76",
         12657 => x"34",
         12658 => x"7b",
         12659 => x"7a",
         12660 => x"34",
         12661 => x"55",
         12662 => x"17",
         12663 => x"a0",
         12664 => x"1a",
         12665 => x"58",
         12666 => x"39",
         12667 => x"58",
         12668 => x"34",
         12669 => x"5c",
         12670 => x"34",
         12671 => x"0b",
         12672 => x"7d",
         12673 => x"83",
         12674 => x"51",
         12675 => x"3f",
         12676 => x"08",
         12677 => x"39",
         12678 => x"b3",
         12679 => x"08",
         12680 => x"5f",
         12681 => x"9b",
         12682 => x"81",
         12683 => x"70",
         12684 => x"56",
         12685 => x"81",
         12686 => x"ed",
         12687 => x"2e",
         12688 => x"82",
         12689 => x"fe",
         12690 => x"b2",
         12691 => x"ab",
         12692 => x"bb",
         12693 => x"84",
         12694 => x"80",
         12695 => x"75",
         12696 => x"0c",
         12697 => x"04",
         12698 => x"0c",
         12699 => x"52",
         12700 => x"52",
         12701 => x"e8",
         12702 => x"84",
         12703 => x"bb",
         12704 => x"38",
         12705 => x"05",
         12706 => x"06",
         12707 => x"7c",
         12708 => x"0b",
         12709 => x"3d",
         12710 => x"55",
         12711 => x"05",
         12712 => x"70",
         12713 => x"34",
         12714 => x"74",
         12715 => x"3d",
         12716 => x"7a",
         12717 => x"75",
         12718 => x"57",
         12719 => x"81",
         12720 => x"ff",
         12721 => x"ef",
         12722 => x"08",
         12723 => x"ff",
         12724 => x"84",
         12725 => x"56",
         12726 => x"08",
         12727 => x"6a",
         12728 => x"2e",
         12729 => x"88",
         12730 => x"84",
         12731 => x"0d",
         12732 => x"d0",
         12733 => x"ff",
         12734 => x"58",
         12735 => x"91",
         12736 => x"78",
         12737 => x"d0",
         12738 => x"78",
         12739 => x"fa",
         12740 => x"08",
         12741 => x"70",
         12742 => x"5e",
         12743 => x"7a",
         12744 => x"5c",
         12745 => x"81",
         12746 => x"ff",
         12747 => x"58",
         12748 => x"26",
         12749 => x"16",
         12750 => x"06",
         12751 => x"9f",
         12752 => x"99",
         12753 => x"e0",
         12754 => x"ff",
         12755 => x"75",
         12756 => x"2a",
         12757 => x"77",
         12758 => x"06",
         12759 => x"ff",
         12760 => x"7a",
         12761 => x"70",
         12762 => x"2a",
         12763 => x"58",
         12764 => x"2e",
         12765 => x"1c",
         12766 => x"5c",
         12767 => x"fd",
         12768 => x"08",
         12769 => x"ff",
         12770 => x"83",
         12771 => x"38",
         12772 => x"82",
         12773 => x"fe",
         12774 => x"b2",
         12775 => x"a9",
         12776 => x"bb",
         12777 => x"84",
         12778 => x"fd",
         12779 => x"b8",
         12780 => x"3d",
         12781 => x"81",
         12782 => x"38",
         12783 => x"8d",
         12784 => x"bb",
         12785 => x"84",
         12786 => x"fd",
         12787 => x"58",
         12788 => x"19",
         12789 => x"80",
         12790 => x"56",
         12791 => x"81",
         12792 => x"75",
         12793 => x"57",
         12794 => x"5a",
         12795 => x"02",
         12796 => x"33",
         12797 => x"8b",
         12798 => x"84",
         12799 => x"40",
         12800 => x"38",
         12801 => x"57",
         12802 => x"34",
         12803 => x"0b",
         12804 => x"8b",
         12805 => x"84",
         12806 => x"57",
         12807 => x"2e",
         12808 => x"a7",
         12809 => x"2e",
         12810 => x"7f",
         12811 => x"9a",
         12812 => x"88",
         12813 => x"33",
         12814 => x"57",
         12815 => x"82",
         12816 => x"16",
         12817 => x"fe",
         12818 => x"75",
         12819 => x"c7",
         12820 => x"22",
         12821 => x"b0",
         12822 => x"57",
         12823 => x"2e",
         12824 => x"75",
         12825 => x"b4",
         12826 => x"2e",
         12827 => x"17",
         12828 => x"83",
         12829 => x"54",
         12830 => x"17",
         12831 => x"33",
         12832 => x"aa",
         12833 => x"84",
         12834 => x"85",
         12835 => x"81",
         12836 => x"18",
         12837 => x"7b",
         12838 => x"56",
         12839 => x"bf",
         12840 => x"33",
         12841 => x"2e",
         12842 => x"bb",
         12843 => x"83",
         12844 => x"5d",
         12845 => x"f2",
         12846 => x"88",
         12847 => x"80",
         12848 => x"76",
         12849 => x"83",
         12850 => x"06",
         12851 => x"90",
         12852 => x"80",
         12853 => x"7d",
         12854 => x"75",
         12855 => x"34",
         12856 => x"0b",
         12857 => x"78",
         12858 => x"08",
         12859 => x"57",
         12860 => x"ff",
         12861 => x"74",
         12862 => x"fe",
         12863 => x"84",
         12864 => x"55",
         12865 => x"08",
         12866 => x"b8",
         12867 => x"19",
         12868 => x"5a",
         12869 => x"77",
         12870 => x"83",
         12871 => x"59",
         12872 => x"2e",
         12873 => x"81",
         12874 => x"54",
         12875 => x"16",
         12876 => x"33",
         12877 => x"f6",
         12878 => x"84",
         12879 => x"85",
         12880 => x"81",
         12881 => x"17",
         12882 => x"77",
         12883 => x"19",
         12884 => x"7a",
         12885 => x"83",
         12886 => x"19",
         12887 => x"a5",
         12888 => x"78",
         12889 => x"e7",
         12890 => x"84",
         12891 => x"bb",
         12892 => x"2e",
         12893 => x"82",
         12894 => x"2e",
         12895 => x"74",
         12896 => x"db",
         12897 => x"fe",
         12898 => x"84",
         12899 => x"84",
         12900 => x"b1",
         12901 => x"82",
         12902 => x"84",
         12903 => x"0d",
         12904 => x"33",
         12905 => x"71",
         12906 => x"90",
         12907 => x"07",
         12908 => x"fd",
         12909 => x"bb",
         12910 => x"2e",
         12911 => x"84",
         12912 => x"80",
         12913 => x"38",
         12914 => x"84",
         12915 => x"0d",
         12916 => x"b4",
         12917 => x"7b",
         12918 => x"33",
         12919 => x"cd",
         12920 => x"84",
         12921 => x"7a",
         12922 => x"06",
         12923 => x"84",
         12924 => x"83",
         12925 => x"16",
         12926 => x"08",
         12927 => x"84",
         12928 => x"74",
         12929 => x"27",
         12930 => x"82",
         12931 => x"7c",
         12932 => x"81",
         12933 => x"38",
         12934 => x"16",
         12935 => x"08",
         12936 => x"52",
         12937 => x"51",
         12938 => x"3f",
         12939 => x"fa",
         12940 => x"b4",
         12941 => x"b8",
         12942 => x"81",
         12943 => x"5b",
         12944 => x"3f",
         12945 => x"bb",
         12946 => x"c9",
         12947 => x"84",
         12948 => x"34",
         12949 => x"a8",
         12950 => x"84",
         12951 => x"5d",
         12952 => x"18",
         12953 => x"8e",
         12954 => x"33",
         12955 => x"2e",
         12956 => x"fc",
         12957 => x"54",
         12958 => x"a0",
         12959 => x"53",
         12960 => x"17",
         12961 => x"e1",
         12962 => x"5c",
         12963 => x"ec",
         12964 => x"80",
         12965 => x"02",
         12966 => x"e3",
         12967 => x"57",
         12968 => x"3d",
         12969 => x"97",
         12970 => x"a3",
         12971 => x"bb",
         12972 => x"84",
         12973 => x"80",
         12974 => x"75",
         12975 => x"0c",
         12976 => x"04",
         12977 => x"52",
         12978 => x"05",
         12979 => x"90",
         12980 => x"84",
         12981 => x"bb",
         12982 => x"38",
         12983 => x"05",
         12984 => x"06",
         12985 => x"73",
         12986 => x"a7",
         12987 => x"09",
         12988 => x"71",
         12989 => x"06",
         12990 => x"57",
         12991 => x"17",
         12992 => x"81",
         12993 => x"34",
         12994 => x"e2",
         12995 => x"bb",
         12996 => x"bb",
         12997 => x"3d",
         12998 => x"3d",
         12999 => x"82",
         13000 => x"cc",
         13001 => x"3d",
         13002 => x"92",
         13003 => x"84",
         13004 => x"bb",
         13005 => x"2e",
         13006 => x"84",
         13007 => x"96",
         13008 => x"78",
         13009 => x"96",
         13010 => x"51",
         13011 => x"3f",
         13012 => x"08",
         13013 => x"84",
         13014 => x"02",
         13015 => x"33",
         13016 => x"56",
         13017 => x"d2",
         13018 => x"18",
         13019 => x"22",
         13020 => x"07",
         13021 => x"76",
         13022 => x"76",
         13023 => x"74",
         13024 => x"76",
         13025 => x"77",
         13026 => x"76",
         13027 => x"73",
         13028 => x"78",
         13029 => x"83",
         13030 => x"51",
         13031 => x"3f",
         13032 => x"08",
         13033 => x"0c",
         13034 => x"04",
         13035 => x"6b",
         13036 => x"80",
         13037 => x"cc",
         13038 => x"3d",
         13039 => x"fe",
         13040 => x"84",
         13041 => x"84",
         13042 => x"84",
         13043 => x"07",
         13044 => x"56",
         13045 => x"2e",
         13046 => x"70",
         13047 => x"56",
         13048 => x"38",
         13049 => x"78",
         13050 => x"56",
         13051 => x"2e",
         13052 => x"81",
         13053 => x"5a",
         13054 => x"2e",
         13055 => x"7c",
         13056 => x"58",
         13057 => x"b4",
         13058 => x"2e",
         13059 => x"83",
         13060 => x"5a",
         13061 => x"2e",
         13062 => x"81",
         13063 => x"54",
         13064 => x"16",
         13065 => x"33",
         13066 => x"82",
         13067 => x"84",
         13068 => x"85",
         13069 => x"81",
         13070 => x"17",
         13071 => x"78",
         13072 => x"70",
         13073 => x"80",
         13074 => x"83",
         13075 => x"80",
         13076 => x"84",
         13077 => x"a7",
         13078 => x"b8",
         13079 => x"33",
         13080 => x"71",
         13081 => x"88",
         13082 => x"14",
         13083 => x"07",
         13084 => x"33",
         13085 => x"0c",
         13086 => x"57",
         13087 => x"84",
         13088 => x"9a",
         13089 => x"7c",
         13090 => x"80",
         13091 => x"70",
         13092 => x"f4",
         13093 => x"bb",
         13094 => x"84",
         13095 => x"80",
         13096 => x"38",
         13097 => x"09",
         13098 => x"b8",
         13099 => x"34",
         13100 => x"b0",
         13101 => x"b4",
         13102 => x"b8",
         13103 => x"81",
         13104 => x"5b",
         13105 => x"3f",
         13106 => x"bb",
         13107 => x"2e",
         13108 => x"fe",
         13109 => x"bb",
         13110 => x"17",
         13111 => x"08",
         13112 => x"31",
         13113 => x"08",
         13114 => x"a0",
         13115 => x"fe",
         13116 => x"16",
         13117 => x"82",
         13118 => x"06",
         13119 => x"77",
         13120 => x"08",
         13121 => x"05",
         13122 => x"81",
         13123 => x"fe",
         13124 => x"79",
         13125 => x"76",
         13126 => x"52",
         13127 => x"51",
         13128 => x"3f",
         13129 => x"08",
         13130 => x"8d",
         13131 => x"39",
         13132 => x"51",
         13133 => x"3f",
         13134 => x"08",
         13135 => x"84",
         13136 => x"38",
         13137 => x"08",
         13138 => x"08",
         13139 => x"59",
         13140 => x"19",
         13141 => x"59",
         13142 => x"75",
         13143 => x"59",
         13144 => x"ec",
         13145 => x"1c",
         13146 => x"76",
         13147 => x"2e",
         13148 => x"ff",
         13149 => x"70",
         13150 => x"58",
         13151 => x"ea",
         13152 => x"39",
         13153 => x"ba",
         13154 => x"0d",
         13155 => x"3d",
         13156 => x"52",
         13157 => x"ff",
         13158 => x"84",
         13159 => x"56",
         13160 => x"08",
         13161 => x"8f",
         13162 => x"7d",
         13163 => x"76",
         13164 => x"58",
         13165 => x"55",
         13166 => x"74",
         13167 => x"70",
         13168 => x"ff",
         13169 => x"58",
         13170 => x"27",
         13171 => x"a2",
         13172 => x"5c",
         13173 => x"ff",
         13174 => x"57",
         13175 => x"f5",
         13176 => x"0c",
         13177 => x"ff",
         13178 => x"38",
         13179 => x"95",
         13180 => x"52",
         13181 => x"08",
         13182 => x"3f",
         13183 => x"08",
         13184 => x"06",
         13185 => x"2e",
         13186 => x"83",
         13187 => x"83",
         13188 => x"70",
         13189 => x"5b",
         13190 => x"80",
         13191 => x"38",
         13192 => x"77",
         13193 => x"81",
         13194 => x"70",
         13195 => x"57",
         13196 => x"80",
         13197 => x"74",
         13198 => x"81",
         13199 => x"75",
         13200 => x"59",
         13201 => x"38",
         13202 => x"27",
         13203 => x"79",
         13204 => x"96",
         13205 => x"77",
         13206 => x"76",
         13207 => x"74",
         13208 => x"05",
         13209 => x"1a",
         13210 => x"70",
         13211 => x"34",
         13212 => x"3d",
         13213 => x"70",
         13214 => x"5b",
         13215 => x"77",
         13216 => x"d1",
         13217 => x"33",
         13218 => x"76",
         13219 => x"bc",
         13220 => x"2e",
         13221 => x"b7",
         13222 => x"16",
         13223 => x"5c",
         13224 => x"09",
         13225 => x"38",
         13226 => x"79",
         13227 => x"45",
         13228 => x"52",
         13229 => x"52",
         13230 => x"9d",
         13231 => x"84",
         13232 => x"bb",
         13233 => x"2e",
         13234 => x"56",
         13235 => x"84",
         13236 => x"0d",
         13237 => x"52",
         13238 => x"e7",
         13239 => x"84",
         13240 => x"ff",
         13241 => x"fd",
         13242 => x"56",
         13243 => x"84",
         13244 => x"0d",
         13245 => x"94",
         13246 => x"c3",
         13247 => x"75",
         13248 => x"a7",
         13249 => x"84",
         13250 => x"bb",
         13251 => x"c1",
         13252 => x"2e",
         13253 => x"8b",
         13254 => x"57",
         13255 => x"81",
         13256 => x"76",
         13257 => x"58",
         13258 => x"55",
         13259 => x"7d",
         13260 => x"83",
         13261 => x"51",
         13262 => x"3f",
         13263 => x"08",
         13264 => x"ff",
         13265 => x"7a",
         13266 => x"38",
         13267 => x"9c",
         13268 => x"84",
         13269 => x"09",
         13270 => x"ee",
         13271 => x"79",
         13272 => x"e6",
         13273 => x"75",
         13274 => x"58",
         13275 => x"3f",
         13276 => x"08",
         13277 => x"84",
         13278 => x"09",
         13279 => x"84",
         13280 => x"84",
         13281 => x"5c",
         13282 => x"08",
         13283 => x"b4",
         13284 => x"2e",
         13285 => x"18",
         13286 => x"79",
         13287 => x"06",
         13288 => x"81",
         13289 => x"b8",
         13290 => x"18",
         13291 => x"d5",
         13292 => x"bb",
         13293 => x"2e",
         13294 => x"57",
         13295 => x"b4",
         13296 => x"57",
         13297 => x"78",
         13298 => x"70",
         13299 => x"57",
         13300 => x"2e",
         13301 => x"74",
         13302 => x"25",
         13303 => x"5c",
         13304 => x"81",
         13305 => x"1a",
         13306 => x"2e",
         13307 => x"52",
         13308 => x"ef",
         13309 => x"bb",
         13310 => x"84",
         13311 => x"80",
         13312 => x"38",
         13313 => x"84",
         13314 => x"38",
         13315 => x"fd",
         13316 => x"6c",
         13317 => x"76",
         13318 => x"58",
         13319 => x"55",
         13320 => x"6b",
         13321 => x"8b",
         13322 => x"6c",
         13323 => x"55",
         13324 => x"05",
         13325 => x"70",
         13326 => x"34",
         13327 => x"74",
         13328 => x"eb",
         13329 => x"81",
         13330 => x"76",
         13331 => x"58",
         13332 => x"55",
         13333 => x"fd",
         13334 => x"5a",
         13335 => x"7d",
         13336 => x"83",
         13337 => x"51",
         13338 => x"3f",
         13339 => x"08",
         13340 => x"39",
         13341 => x"df",
         13342 => x"b4",
         13343 => x"7a",
         13344 => x"33",
         13345 => x"a5",
         13346 => x"84",
         13347 => x"09",
         13348 => x"c3",
         13349 => x"84",
         13350 => x"34",
         13351 => x"a8",
         13352 => x"5c",
         13353 => x"08",
         13354 => x"82",
         13355 => x"74",
         13356 => x"38",
         13357 => x"08",
         13358 => x"39",
         13359 => x"52",
         13360 => x"ee",
         13361 => x"bb",
         13362 => x"84",
         13363 => x"80",
         13364 => x"38",
         13365 => x"81",
         13366 => x"78",
         13367 => x"e7",
         13368 => x"39",
         13369 => x"18",
         13370 => x"08",
         13371 => x"52",
         13372 => x"51",
         13373 => x"3f",
         13374 => x"f2",
         13375 => x"62",
         13376 => x"80",
         13377 => x"5e",
         13378 => x"56",
         13379 => x"9f",
         13380 => x"55",
         13381 => x"97",
         13382 => x"54",
         13383 => x"8f",
         13384 => x"22",
         13385 => x"59",
         13386 => x"2e",
         13387 => x"80",
         13388 => x"75",
         13389 => x"91",
         13390 => x"75",
         13391 => x"79",
         13392 => x"a2",
         13393 => x"08",
         13394 => x"90",
         13395 => x"81",
         13396 => x"56",
         13397 => x"2e",
         13398 => x"7e",
         13399 => x"70",
         13400 => x"55",
         13401 => x"5c",
         13402 => x"bc",
         13403 => x"7a",
         13404 => x"70",
         13405 => x"2a",
         13406 => x"08",
         13407 => x"08",
         13408 => x"5f",
         13409 => x"78",
         13410 => x"9c",
         13411 => x"26",
         13412 => x"58",
         13413 => x"5b",
         13414 => x"52",
         13415 => x"d8",
         13416 => x"15",
         13417 => x"9c",
         13418 => x"26",
         13419 => x"55",
         13420 => x"08",
         13421 => x"dc",
         13422 => x"84",
         13423 => x"81",
         13424 => x"bb",
         13425 => x"c5",
         13426 => x"59",
         13427 => x"bb",
         13428 => x"2e",
         13429 => x"c2",
         13430 => x"75",
         13431 => x"bb",
         13432 => x"3d",
         13433 => x"0b",
         13434 => x"0c",
         13435 => x"04",
         13436 => x"51",
         13437 => x"3f",
         13438 => x"08",
         13439 => x"73",
         13440 => x"73",
         13441 => x"56",
         13442 => x"7b",
         13443 => x"8e",
         13444 => x"56",
         13445 => x"2e",
         13446 => x"18",
         13447 => x"2e",
         13448 => x"73",
         13449 => x"7e",
         13450 => x"96",
         13451 => x"84",
         13452 => x"bb",
         13453 => x"a3",
         13454 => x"19",
         13455 => x"59",
         13456 => x"38",
         13457 => x"12",
         13458 => x"80",
         13459 => x"38",
         13460 => x"0c",
         13461 => x"0c",
         13462 => x"80",
         13463 => x"7b",
         13464 => x"9c",
         13465 => x"05",
         13466 => x"58",
         13467 => x"26",
         13468 => x"76",
         13469 => x"16",
         13470 => x"33",
         13471 => x"7c",
         13472 => x"75",
         13473 => x"39",
         13474 => x"97",
         13475 => x"80",
         13476 => x"39",
         13477 => x"c5",
         13478 => x"fe",
         13479 => x"1b",
         13480 => x"39",
         13481 => x"08",
         13482 => x"a3",
         13483 => x"3d",
         13484 => x"05",
         13485 => x"33",
         13486 => x"ff",
         13487 => x"08",
         13488 => x"40",
         13489 => x"85",
         13490 => x"70",
         13491 => x"33",
         13492 => x"56",
         13493 => x"2e",
         13494 => x"74",
         13495 => x"ba",
         13496 => x"38",
         13497 => x"33",
         13498 => x"24",
         13499 => x"75",
         13500 => x"e2",
         13501 => x"08",
         13502 => x"80",
         13503 => x"80",
         13504 => x"16",
         13505 => x"11",
         13506 => x"f9",
         13507 => x"5b",
         13508 => x"79",
         13509 => x"e2",
         13510 => x"84",
         13511 => x"06",
         13512 => x"5d",
         13513 => x"7b",
         13514 => x"75",
         13515 => x"06",
         13516 => x"7f",
         13517 => x"9f",
         13518 => x"53",
         13519 => x"51",
         13520 => x"3f",
         13521 => x"08",
         13522 => x"6d",
         13523 => x"2e",
         13524 => x"74",
         13525 => x"26",
         13526 => x"ff",
         13527 => x"55",
         13528 => x"38",
         13529 => x"88",
         13530 => x"7f",
         13531 => x"38",
         13532 => x"0a",
         13533 => x"38",
         13534 => x"06",
         13535 => x"e7",
         13536 => x"2a",
         13537 => x"89",
         13538 => x"2b",
         13539 => x"47",
         13540 => x"2e",
         13541 => x"65",
         13542 => x"25",
         13543 => x"5f",
         13544 => x"83",
         13545 => x"80",
         13546 => x"38",
         13547 => x"53",
         13548 => x"51",
         13549 => x"3f",
         13550 => x"bb",
         13551 => x"95",
         13552 => x"ff",
         13553 => x"83",
         13554 => x"71",
         13555 => x"59",
         13556 => x"77",
         13557 => x"2e",
         13558 => x"82",
         13559 => x"90",
         13560 => x"83",
         13561 => x"44",
         13562 => x"2e",
         13563 => x"83",
         13564 => x"11",
         13565 => x"33",
         13566 => x"71",
         13567 => x"81",
         13568 => x"72",
         13569 => x"75",
         13570 => x"83",
         13571 => x"11",
         13572 => x"33",
         13573 => x"71",
         13574 => x"81",
         13575 => x"72",
         13576 => x"75",
         13577 => x"5c",
         13578 => x"42",
         13579 => x"a3",
         13580 => x"4e",
         13581 => x"4f",
         13582 => x"78",
         13583 => x"80",
         13584 => x"82",
         13585 => x"57",
         13586 => x"26",
         13587 => x"61",
         13588 => x"81",
         13589 => x"63",
         13590 => x"f9",
         13591 => x"06",
         13592 => x"2e",
         13593 => x"81",
         13594 => x"83",
         13595 => x"6e",
         13596 => x"46",
         13597 => x"62",
         13598 => x"c2",
         13599 => x"38",
         13600 => x"57",
         13601 => x"e8",
         13602 => x"58",
         13603 => x"9d",
         13604 => x"26",
         13605 => x"e8",
         13606 => x"10",
         13607 => x"22",
         13608 => x"74",
         13609 => x"38",
         13610 => x"ee",
         13611 => x"78",
         13612 => x"f4",
         13613 => x"84",
         13614 => x"05",
         13615 => x"84",
         13616 => x"26",
         13617 => x"0b",
         13618 => x"08",
         13619 => x"84",
         13620 => x"11",
         13621 => x"05",
         13622 => x"83",
         13623 => x"2a",
         13624 => x"a0",
         13625 => x"7d",
         13626 => x"66",
         13627 => x"70",
         13628 => x"31",
         13629 => x"44",
         13630 => x"89",
         13631 => x"1d",
         13632 => x"29",
         13633 => x"31",
         13634 => x"79",
         13635 => x"38",
         13636 => x"7d",
         13637 => x"70",
         13638 => x"56",
         13639 => x"3f",
         13640 => x"08",
         13641 => x"2e",
         13642 => x"62",
         13643 => x"81",
         13644 => x"38",
         13645 => x"0b",
         13646 => x"08",
         13647 => x"38",
         13648 => x"38",
         13649 => x"74",
         13650 => x"89",
         13651 => x"5b",
         13652 => x"8b",
         13653 => x"bb",
         13654 => x"3d",
         13655 => x"90",
         13656 => x"4e",
         13657 => x"93",
         13658 => x"84",
         13659 => x"0d",
         13660 => x"0c",
         13661 => x"d0",
         13662 => x"ff",
         13663 => x"57",
         13664 => x"91",
         13665 => x"77",
         13666 => x"d0",
         13667 => x"77",
         13668 => x"b2",
         13669 => x"83",
         13670 => x"5c",
         13671 => x"57",
         13672 => x"81",
         13673 => x"76",
         13674 => x"58",
         13675 => x"12",
         13676 => x"62",
         13677 => x"38",
         13678 => x"81",
         13679 => x"44",
         13680 => x"45",
         13681 => x"89",
         13682 => x"70",
         13683 => x"59",
         13684 => x"70",
         13685 => x"47",
         13686 => x"09",
         13687 => x"38",
         13688 => x"38",
         13689 => x"70",
         13690 => x"07",
         13691 => x"07",
         13692 => x"7a",
         13693 => x"ce",
         13694 => x"84",
         13695 => x"83",
         13696 => x"98",
         13697 => x"f9",
         13698 => x"3d",
         13699 => x"81",
         13700 => x"fe",
         13701 => x"81",
         13702 => x"84",
         13703 => x"38",
         13704 => x"77",
         13705 => x"84",
         13706 => x"75",
         13707 => x"5f",
         13708 => x"57",
         13709 => x"fe",
         13710 => x"7f",
         13711 => x"fb",
         13712 => x"fa",
         13713 => x"83",
         13714 => x"38",
         13715 => x"3d",
         13716 => x"95",
         13717 => x"06",
         13718 => x"67",
         13719 => x"f5",
         13720 => x"70",
         13721 => x"43",
         13722 => x"84",
         13723 => x"9f",
         13724 => x"38",
         13725 => x"77",
         13726 => x"80",
         13727 => x"f5",
         13728 => x"76",
         13729 => x"0c",
         13730 => x"84",
         13731 => x"04",
         13732 => x"81",
         13733 => x"38",
         13734 => x"27",
         13735 => x"81",
         13736 => x"57",
         13737 => x"38",
         13738 => x"57",
         13739 => x"70",
         13740 => x"34",
         13741 => x"74",
         13742 => x"61",
         13743 => x"59",
         13744 => x"70",
         13745 => x"33",
         13746 => x"05",
         13747 => x"15",
         13748 => x"38",
         13749 => x"45",
         13750 => x"82",
         13751 => x"34",
         13752 => x"05",
         13753 => x"ff",
         13754 => x"6a",
         13755 => x"34",
         13756 => x"5c",
         13757 => x"05",
         13758 => x"90",
         13759 => x"83",
         13760 => x"5a",
         13761 => x"91",
         13762 => x"9e",
         13763 => x"49",
         13764 => x"05",
         13765 => x"75",
         13766 => x"26",
         13767 => x"75",
         13768 => x"06",
         13769 => x"93",
         13770 => x"88",
         13771 => x"61",
         13772 => x"f8",
         13773 => x"34",
         13774 => x"05",
         13775 => x"99",
         13776 => x"61",
         13777 => x"80",
         13778 => x"34",
         13779 => x"05",
         13780 => x"2a",
         13781 => x"9d",
         13782 => x"90",
         13783 => x"61",
         13784 => x"7e",
         13785 => x"bb",
         13786 => x"bb",
         13787 => x"9f",
         13788 => x"83",
         13789 => x"38",
         13790 => x"05",
         13791 => x"a8",
         13792 => x"61",
         13793 => x"80",
         13794 => x"05",
         13795 => x"ff",
         13796 => x"74",
         13797 => x"34",
         13798 => x"4b",
         13799 => x"05",
         13800 => x"61",
         13801 => x"a9",
         13802 => x"34",
         13803 => x"05",
         13804 => x"59",
         13805 => x"70",
         13806 => x"33",
         13807 => x"05",
         13808 => x"15",
         13809 => x"38",
         13810 => x"05",
         13811 => x"69",
         13812 => x"ff",
         13813 => x"aa",
         13814 => x"54",
         13815 => x"52",
         13816 => x"c6",
         13817 => x"57",
         13818 => x"08",
         13819 => x"60",
         13820 => x"83",
         13821 => x"38",
         13822 => x"55",
         13823 => x"81",
         13824 => x"ff",
         13825 => x"f4",
         13826 => x"41",
         13827 => x"2e",
         13828 => x"87",
         13829 => x"57",
         13830 => x"83",
         13831 => x"76",
         13832 => x"88",
         13833 => x"55",
         13834 => x"81",
         13835 => x"76",
         13836 => x"78",
         13837 => x"05",
         13838 => x"98",
         13839 => x"64",
         13840 => x"65",
         13841 => x"26",
         13842 => x"59",
         13843 => x"53",
         13844 => x"51",
         13845 => x"3f",
         13846 => x"08",
         13847 => x"84",
         13848 => x"55",
         13849 => x"81",
         13850 => x"ff",
         13851 => x"f4",
         13852 => x"77",
         13853 => x"5b",
         13854 => x"7f",
         13855 => x"7f",
         13856 => x"89",
         13857 => x"62",
         13858 => x"38",
         13859 => x"55",
         13860 => x"83",
         13861 => x"74",
         13862 => x"60",
         13863 => x"fe",
         13864 => x"84",
         13865 => x"85",
         13866 => x"1b",
         13867 => x"57",
         13868 => x"38",
         13869 => x"83",
         13870 => x"86",
         13871 => x"ff",
         13872 => x"38",
         13873 => x"82",
         13874 => x"81",
         13875 => x"c1",
         13876 => x"2a",
         13877 => x"7d",
         13878 => x"84",
         13879 => x"59",
         13880 => x"81",
         13881 => x"ff",
         13882 => x"f4",
         13883 => x"69",
         13884 => x"6b",
         13885 => x"be",
         13886 => x"67",
         13887 => x"81",
         13888 => x"67",
         13889 => x"78",
         13890 => x"34",
         13891 => x"05",
         13892 => x"80",
         13893 => x"62",
         13894 => x"f7",
         13895 => x"67",
         13896 => x"84",
         13897 => x"82",
         13898 => x"57",
         13899 => x"05",
         13900 => x"84",
         13901 => x"05",
         13902 => x"83",
         13903 => x"67",
         13904 => x"05",
         13905 => x"83",
         13906 => x"84",
         13907 => x"61",
         13908 => x"34",
         13909 => x"ca",
         13910 => x"88",
         13911 => x"61",
         13912 => x"34",
         13913 => x"58",
         13914 => x"cc",
         13915 => x"98",
         13916 => x"61",
         13917 => x"34",
         13918 => x"53",
         13919 => x"51",
         13920 => x"3f",
         13921 => x"bb",
         13922 => x"c9",
         13923 => x"80",
         13924 => x"fe",
         13925 => x"81",
         13926 => x"84",
         13927 => x"38",
         13928 => x"08",
         13929 => x"0c",
         13930 => x"84",
         13931 => x"04",
         13932 => x"e4",
         13933 => x"64",
         13934 => x"f6",
         13935 => x"ae",
         13936 => x"2a",
         13937 => x"83",
         13938 => x"56",
         13939 => x"2e",
         13940 => x"77",
         13941 => x"83",
         13942 => x"77",
         13943 => x"70",
         13944 => x"58",
         13945 => x"86",
         13946 => x"27",
         13947 => x"52",
         13948 => x"f5",
         13949 => x"bb",
         13950 => x"10",
         13951 => x"70",
         13952 => x"5c",
         13953 => x"0b",
         13954 => x"08",
         13955 => x"05",
         13956 => x"ff",
         13957 => x"27",
         13958 => x"8e",
         13959 => x"39",
         13960 => x"08",
         13961 => x"26",
         13962 => x"7a",
         13963 => x"77",
         13964 => x"7a",
         13965 => x"8e",
         13966 => x"39",
         13967 => x"44",
         13968 => x"f8",
         13969 => x"43",
         13970 => x"75",
         13971 => x"34",
         13972 => x"49",
         13973 => x"05",
         13974 => x"2a",
         13975 => x"a2",
         13976 => x"98",
         13977 => x"61",
         13978 => x"f9",
         13979 => x"61",
         13980 => x"34",
         13981 => x"c4",
         13982 => x"61",
         13983 => x"34",
         13984 => x"80",
         13985 => x"7c",
         13986 => x"34",
         13987 => x"5c",
         13988 => x"05",
         13989 => x"2a",
         13990 => x"a6",
         13991 => x"98",
         13992 => x"61",
         13993 => x"82",
         13994 => x"34",
         13995 => x"05",
         13996 => x"ae",
         13997 => x"61",
         13998 => x"81",
         13999 => x"34",
         14000 => x"05",
         14001 => x"b2",
         14002 => x"61",
         14003 => x"ff",
         14004 => x"c0",
         14005 => x"61",
         14006 => x"34",
         14007 => x"c7",
         14008 => x"e0",
         14009 => x"76",
         14010 => x"58",
         14011 => x"81",
         14012 => x"ff",
         14013 => x"80",
         14014 => x"38",
         14015 => x"05",
         14016 => x"70",
         14017 => x"34",
         14018 => x"74",
         14019 => x"b8",
         14020 => x"80",
         14021 => x"79",
         14022 => x"92",
         14023 => x"84",
         14024 => x"f4",
         14025 => x"90",
         14026 => x"42",
         14027 => x"b2",
         14028 => x"54",
         14029 => x"08",
         14030 => x"79",
         14031 => x"ed",
         14032 => x"39",
         14033 => x"bb",
         14034 => x"3d",
         14035 => x"90",
         14036 => x"61",
         14037 => x"ff",
         14038 => x"05",
         14039 => x"6a",
         14040 => x"4c",
         14041 => x"34",
         14042 => x"05",
         14043 => x"85",
         14044 => x"61",
         14045 => x"ff",
         14046 => x"34",
         14047 => x"05",
         14048 => x"89",
         14049 => x"61",
         14050 => x"8f",
         14051 => x"57",
         14052 => x"76",
         14053 => x"53",
         14054 => x"51",
         14055 => x"3f",
         14056 => x"56",
         14057 => x"70",
         14058 => x"34",
         14059 => x"76",
         14060 => x"5c",
         14061 => x"70",
         14062 => x"34",
         14063 => x"d2",
         14064 => x"05",
         14065 => x"e1",
         14066 => x"05",
         14067 => x"c1",
         14068 => x"f2",
         14069 => x"05",
         14070 => x"61",
         14071 => x"34",
         14072 => x"83",
         14073 => x"80",
         14074 => x"e7",
         14075 => x"ff",
         14076 => x"61",
         14077 => x"34",
         14078 => x"59",
         14079 => x"e9",
         14080 => x"90",
         14081 => x"61",
         14082 => x"34",
         14083 => x"40",
         14084 => x"eb",
         14085 => x"61",
         14086 => x"34",
         14087 => x"ed",
         14088 => x"61",
         14089 => x"34",
         14090 => x"ef",
         14091 => x"d5",
         14092 => x"aa",
         14093 => x"54",
         14094 => x"60",
         14095 => x"fe",
         14096 => x"81",
         14097 => x"53",
         14098 => x"51",
         14099 => x"3f",
         14100 => x"55",
         14101 => x"f4",
         14102 => x"61",
         14103 => x"7b",
         14104 => x"5a",
         14105 => x"78",
         14106 => x"8d",
         14107 => x"3d",
         14108 => x"81",
         14109 => x"79",
         14110 => x"cc",
         14111 => x"2e",
         14112 => x"9e",
         14113 => x"33",
         14114 => x"2e",
         14115 => x"76",
         14116 => x"58",
         14117 => x"57",
         14118 => x"86",
         14119 => x"24",
         14120 => x"76",
         14121 => x"76",
         14122 => x"55",
         14123 => x"84",
         14124 => x"0d",
         14125 => x"0d",
         14126 => x"05",
         14127 => x"59",
         14128 => x"2e",
         14129 => x"84",
         14130 => x"80",
         14131 => x"38",
         14132 => x"77",
         14133 => x"56",
         14134 => x"34",
         14135 => x"74",
         14136 => x"38",
         14137 => x"0c",
         14138 => x"18",
         14139 => x"0d",
         14140 => x"fc",
         14141 => x"53",
         14142 => x"76",
         14143 => x"9f",
         14144 => x"7a",
         14145 => x"70",
         14146 => x"2a",
         14147 => x"1b",
         14148 => x"88",
         14149 => x"56",
         14150 => x"8d",
         14151 => x"ff",
         14152 => x"a3",
         14153 => x"0d",
         14154 => x"05",
         14155 => x"58",
         14156 => x"77",
         14157 => x"76",
         14158 => x"58",
         14159 => x"55",
         14160 => x"a1",
         14161 => x"0c",
         14162 => x"80",
         14163 => x"56",
         14164 => x"80",
         14165 => x"77",
         14166 => x"56",
         14167 => x"34",
         14168 => x"74",
         14169 => x"38",
         14170 => x"0c",
         14171 => x"18",
         14172 => x"80",
         14173 => x"38",
         14174 => x"ac",
         14175 => x"54",
         14176 => x"76",
         14177 => x"9e",
         14178 => x"bb",
         14179 => x"38",
         14180 => x"ba",
         14181 => x"84",
         14182 => x"9f",
         14183 => x"9f",
         14184 => x"11",
         14185 => x"c0",
         14186 => x"08",
         14187 => x"f8",
         14188 => x"32",
         14189 => x"72",
         14190 => x"70",
         14191 => x"56",
         14192 => x"39",
         14193 => x"51",
         14194 => x"ff",
         14195 => x"84",
         14196 => x"9f",
         14197 => x"fd",
         14198 => x"02",
         14199 => x"05",
         14200 => x"80",
         14201 => x"ff",
         14202 => x"72",
         14203 => x"06",
         14204 => x"bb",
         14205 => x"3d",
         14206 => x"ff",
         14207 => x"54",
         14208 => x"2e",
         14209 => x"e9",
         14210 => x"2e",
         14211 => x"e8",
         14212 => x"72",
         14213 => x"38",
         14214 => x"83",
         14215 => x"53",
         14216 => x"ff",
         14217 => x"71",
         14218 => x"c8",
         14219 => x"51",
         14220 => x"81",
         14221 => x"81",
         14222 => x"bb",
         14223 => x"85",
         14224 => x"fe",
         14225 => x"92",
         14226 => x"84",
         14227 => x"22",
         14228 => x"53",
         14229 => x"26",
         14230 => x"53",
         14231 => x"84",
         14232 => x"0d",
         14233 => x"b5",
         14234 => x"06",
         14235 => x"81",
         14236 => x"38",
         14237 => x"e6",
         14238 => x"22",
         14239 => x"0c",
         14240 => x"0d",
         14241 => x"0d",
         14242 => x"83",
         14243 => x"80",
         14244 => x"83",
         14245 => x"83",
         14246 => x"56",
         14247 => x"26",
         14248 => x"74",
         14249 => x"56",
         14250 => x"30",
         14251 => x"73",
         14252 => x"54",
         14253 => x"70",
         14254 => x"70",
         14255 => x"22",
         14256 => x"2a",
         14257 => x"ff",
         14258 => x"52",
         14259 => x"24",
         14260 => x"cf",
         14261 => x"15",
         14262 => x"05",
         14263 => x"73",
         14264 => x"25",
         14265 => x"07",
         14266 => x"70",
         14267 => x"38",
         14268 => x"84",
         14269 => x"87",
         14270 => x"83",
         14271 => x"ff",
         14272 => x"88",
         14273 => x"71",
         14274 => x"ca",
         14275 => x"73",
         14276 => x"a0",
         14277 => x"ff",
         14278 => x"51",
         14279 => x"39",
         14280 => x"70",
         14281 => x"06",
         14282 => x"39",
         14283 => x"83",
         14284 => x"57",
         14285 => x"e6",
         14286 => x"ff",
         14287 => x"51",
         14288 => x"16",
         14289 => x"ff",
         14290 => x"d0",
         14291 => x"70",
         14292 => x"06",
         14293 => x"39",
         14294 => x"83",
         14295 => x"57",
         14296 => x"39",
         14297 => x"81",
         14298 => x"31",
         14299 => x"ff",
         14300 => x"55",
         14301 => x"75",
         14302 => x"75",
         14303 => x"52",
         14304 => x"39",
         14305 => x"00",
         14306 => x"ff",
         14307 => x"ff",
         14308 => x"ff",
         14309 => x"00",
         14310 => x"00",
         14311 => x"00",
         14312 => x"00",
         14313 => x"00",
         14314 => x"00",
         14315 => x"00",
         14316 => x"00",
         14317 => x"00",
         14318 => x"00",
         14319 => x"00",
         14320 => x"00",
         14321 => x"00",
         14322 => x"00",
         14323 => x"00",
         14324 => x"00",
         14325 => x"00",
         14326 => x"00",
         14327 => x"00",
         14328 => x"00",
         14329 => x"00",
         14330 => x"00",
         14331 => x"00",
         14332 => x"00",
         14333 => x"00",
         14334 => x"00",
         14335 => x"00",
         14336 => x"00",
         14337 => x"00",
         14338 => x"00",
         14339 => x"00",
         14340 => x"00",
         14341 => x"00",
         14342 => x"00",
         14343 => x"00",
         14344 => x"00",
         14345 => x"00",
         14346 => x"00",
         14347 => x"00",
         14348 => x"00",
         14349 => x"00",
         14350 => x"00",
         14351 => x"00",
         14352 => x"00",
         14353 => x"00",
         14354 => x"00",
         14355 => x"00",
         14356 => x"00",
         14357 => x"00",
         14358 => x"00",
         14359 => x"00",
         14360 => x"00",
         14361 => x"00",
         14362 => x"00",
         14363 => x"00",
         14364 => x"00",
         14365 => x"00",
         14366 => x"00",
         14367 => x"00",
         14368 => x"00",
         14369 => x"00",
         14370 => x"00",
         14371 => x"00",
         14372 => x"00",
         14373 => x"00",
         14374 => x"00",
         14375 => x"00",
         14376 => x"00",
         14377 => x"00",
         14378 => x"00",
         14379 => x"00",
         14380 => x"00",
         14381 => x"00",
         14382 => x"00",
         14383 => x"00",
         14384 => x"00",
         14385 => x"00",
         14386 => x"00",
         14387 => x"00",
         14388 => x"00",
         14389 => x"00",
         14390 => x"00",
         14391 => x"00",
         14392 => x"00",
         14393 => x"00",
         14394 => x"00",
         14395 => x"00",
         14396 => x"00",
         14397 => x"00",
         14398 => x"00",
         14399 => x"00",
         14400 => x"00",
         14401 => x"00",
         14402 => x"00",
         14403 => x"00",
         14404 => x"00",
         14405 => x"00",
         14406 => x"00",
         14407 => x"00",
         14408 => x"00",
         14409 => x"00",
         14410 => x"00",
         14411 => x"00",
         14412 => x"00",
         14413 => x"00",
         14414 => x"00",
         14415 => x"00",
         14416 => x"00",
         14417 => x"00",
         14418 => x"00",
         14419 => x"00",
         14420 => x"00",
         14421 => x"00",
         14422 => x"00",
         14423 => x"00",
         14424 => x"00",
         14425 => x"00",
         14426 => x"00",
         14427 => x"00",
         14428 => x"00",
         14429 => x"00",
         14430 => x"00",
         14431 => x"00",
         14432 => x"00",
         14433 => x"00",
         14434 => x"00",
         14435 => x"00",
         14436 => x"00",
         14437 => x"00",
         14438 => x"00",
         14439 => x"00",
         14440 => x"00",
         14441 => x"00",
         14442 => x"00",
         14443 => x"00",
         14444 => x"00",
         14445 => x"00",
         14446 => x"00",
         14447 => x"00",
         14448 => x"00",
         14449 => x"00",
         14450 => x"00",
         14451 => x"00",
         14452 => x"00",
         14453 => x"00",
         14454 => x"00",
         14455 => x"00",
         14456 => x"00",
         14457 => x"00",
         14458 => x"00",
         14459 => x"00",
         14460 => x"00",
         14461 => x"00",
         14462 => x"00",
         14463 => x"00",
         14464 => x"00",
         14465 => x"00",
         14466 => x"00",
         14467 => x"00",
         14468 => x"00",
         14469 => x"00",
         14470 => x"00",
         14471 => x"00",
         14472 => x"00",
         14473 => x"00",
         14474 => x"00",
         14475 => x"00",
         14476 => x"00",
         14477 => x"00",
         14478 => x"00",
         14479 => x"00",
         14480 => x"00",
         14481 => x"00",
         14482 => x"00",
         14483 => x"00",
         14484 => x"00",
         14485 => x"00",
         14486 => x"00",
         14487 => x"00",
         14488 => x"00",
         14489 => x"00",
         14490 => x"00",
         14491 => x"00",
         14492 => x"00",
         14493 => x"00",
         14494 => x"00",
         14495 => x"00",
         14496 => x"00",
         14497 => x"00",
         14498 => x"00",
         14499 => x"00",
         14500 => x"00",
         14501 => x"00",
         14502 => x"00",
         14503 => x"00",
         14504 => x"00",
         14505 => x"00",
         14506 => x"00",
         14507 => x"00",
         14508 => x"00",
         14509 => x"00",
         14510 => x"00",
         14511 => x"00",
         14512 => x"00",
         14513 => x"00",
         14514 => x"00",
         14515 => x"00",
         14516 => x"00",
         14517 => x"00",
         14518 => x"00",
         14519 => x"00",
         14520 => x"00",
         14521 => x"00",
         14522 => x"00",
         14523 => x"00",
         14524 => x"00",
         14525 => x"00",
         14526 => x"00",
         14527 => x"00",
         14528 => x"00",
         14529 => x"00",
         14530 => x"00",
         14531 => x"00",
         14532 => x"00",
         14533 => x"00",
         14534 => x"00",
         14535 => x"00",
         14536 => x"00",
         14537 => x"00",
         14538 => x"00",
         14539 => x"00",
         14540 => x"00",
         14541 => x"00",
         14542 => x"00",
         14543 => x"00",
         14544 => x"00",
         14545 => x"00",
         14546 => x"00",
         14547 => x"00",
         14548 => x"00",
         14549 => x"00",
         14550 => x"00",
         14551 => x"00",
         14552 => x"00",
         14553 => x"00",
         14554 => x"00",
         14555 => x"00",
         14556 => x"00",
         14557 => x"00",
         14558 => x"00",
         14559 => x"00",
         14560 => x"00",
         14561 => x"00",
         14562 => x"00",
         14563 => x"00",
         14564 => x"00",
         14565 => x"00",
         14566 => x"00",
         14567 => x"00",
         14568 => x"00",
         14569 => x"00",
         14570 => x"00",
         14571 => x"00",
         14572 => x"00",
         14573 => x"00",
         14574 => x"00",
         14575 => x"00",
         14576 => x"00",
         14577 => x"00",
         14578 => x"00",
         14579 => x"00",
         14580 => x"00",
         14581 => x"00",
         14582 => x"00",
         14583 => x"00",
         14584 => x"00",
         14585 => x"00",
         14586 => x"00",
         14587 => x"00",
         14588 => x"00",
         14589 => x"00",
         14590 => x"00",
         14591 => x"00",
         14592 => x"00",
         14593 => x"00",
         14594 => x"00",
         14595 => x"00",
         14596 => x"00",
         14597 => x"00",
         14598 => x"00",
         14599 => x"00",
         14600 => x"00",
         14601 => x"00",
         14602 => x"00",
         14603 => x"00",
         14604 => x"00",
         14605 => x"00",
         14606 => x"00",
         14607 => x"00",
         14608 => x"00",
         14609 => x"00",
         14610 => x"00",
         14611 => x"00",
         14612 => x"00",
         14613 => x"00",
         14614 => x"00",
         14615 => x"00",
         14616 => x"00",
         14617 => x"00",
         14618 => x"00",
         14619 => x"00",
         14620 => x"00",
         14621 => x"00",
         14622 => x"00",
         14623 => x"00",
         14624 => x"00",
         14625 => x"00",
         14626 => x"00",
         14627 => x"00",
         14628 => x"00",
         14629 => x"00",
         14630 => x"00",
         14631 => x"00",
         14632 => x"00",
         14633 => x"00",
         14634 => x"00",
         14635 => x"00",
         14636 => x"00",
         14637 => x"00",
         14638 => x"00",
         14639 => x"00",
         14640 => x"00",
         14641 => x"00",
         14642 => x"00",
         14643 => x"00",
         14644 => x"00",
         14645 => x"00",
         14646 => x"00",
         14647 => x"00",
         14648 => x"00",
         14649 => x"00",
         14650 => x"00",
         14651 => x"00",
         14652 => x"00",
         14653 => x"00",
         14654 => x"00",
         14655 => x"00",
         14656 => x"00",
         14657 => x"00",
         14658 => x"00",
         14659 => x"00",
         14660 => x"00",
         14661 => x"00",
         14662 => x"00",
         14663 => x"00",
         14664 => x"00",
         14665 => x"00",
         14666 => x"00",
         14667 => x"00",
         14668 => x"00",
         14669 => x"00",
         14670 => x"00",
         14671 => x"00",
         14672 => x"00",
         14673 => x"00",
         14674 => x"00",
         14675 => x"00",
         14676 => x"00",
         14677 => x"00",
         14678 => x"00",
         14679 => x"00",
         14680 => x"00",
         14681 => x"00",
         14682 => x"00",
         14683 => x"00",
         14684 => x"00",
         14685 => x"00",
         14686 => x"00",
         14687 => x"00",
         14688 => x"00",
         14689 => x"00",
         14690 => x"00",
         14691 => x"00",
         14692 => x"00",
         14693 => x"00",
         14694 => x"00",
         14695 => x"00",
         14696 => x"00",
         14697 => x"00",
         14698 => x"00",
         14699 => x"00",
         14700 => x"00",
         14701 => x"00",
         14702 => x"00",
         14703 => x"00",
         14704 => x"00",
         14705 => x"00",
         14706 => x"00",
         14707 => x"00",
         14708 => x"00",
         14709 => x"00",
         14710 => x"00",
         14711 => x"00",
         14712 => x"00",
         14713 => x"00",
         14714 => x"00",
         14715 => x"00",
         14716 => x"00",
         14717 => x"00",
         14718 => x"00",
         14719 => x"00",
         14720 => x"00",
         14721 => x"00",
         14722 => x"00",
         14723 => x"00",
         14724 => x"00",
         14725 => x"00",
         14726 => x"00",
         14727 => x"00",
         14728 => x"00",
         14729 => x"00",
         14730 => x"00",
         14731 => x"00",
         14732 => x"00",
         14733 => x"00",
         14734 => x"00",
         14735 => x"00",
         14736 => x"00",
         14737 => x"00",
         14738 => x"00",
         14739 => x"00",
         14740 => x"00",
         14741 => x"00",
         14742 => x"00",
         14743 => x"00",
         14744 => x"00",
         14745 => x"00",
         14746 => x"00",
         14747 => x"00",
         14748 => x"00",
         14749 => x"00",
         14750 => x"00",
         14751 => x"00",
         14752 => x"00",
         14753 => x"00",
         14754 => x"00",
         14755 => x"00",
         14756 => x"00",
         14757 => x"00",
         14758 => x"00",
         14759 => x"00",
         14760 => x"00",
         14761 => x"00",
         14762 => x"00",
         14763 => x"00",
         14764 => x"00",
         14765 => x"00",
         14766 => x"00",
         14767 => x"00",
         14768 => x"00",
         14769 => x"00",
         14770 => x"00",
         14771 => x"00",
         14772 => x"00",
         14773 => x"00",
         14774 => x"00",
         14775 => x"00",
         14776 => x"00",
         14777 => x"00",
         14778 => x"00",
         14779 => x"00",
         14780 => x"00",
         14781 => x"00",
         14782 => x"64",
         14783 => x"74",
         14784 => x"64",
         14785 => x"74",
         14786 => x"66",
         14787 => x"74",
         14788 => x"66",
         14789 => x"64",
         14790 => x"66",
         14791 => x"63",
         14792 => x"6d",
         14793 => x"61",
         14794 => x"6d",
         14795 => x"79",
         14796 => x"6d",
         14797 => x"66",
         14798 => x"6d",
         14799 => x"70",
         14800 => x"6d",
         14801 => x"6d",
         14802 => x"6d",
         14803 => x"68",
         14804 => x"68",
         14805 => x"68",
         14806 => x"68",
         14807 => x"63",
         14808 => x"00",
         14809 => x"6a",
         14810 => x"72",
         14811 => x"61",
         14812 => x"72",
         14813 => x"74",
         14814 => x"69",
         14815 => x"00",
         14816 => x"74",
         14817 => x"00",
         14818 => x"63",
         14819 => x"7a",
         14820 => x"74",
         14821 => x"69",
         14822 => x"6d",
         14823 => x"69",
         14824 => x"6b",
         14825 => x"00",
         14826 => x"65",
         14827 => x"55",
         14828 => x"6f",
         14829 => x"65",
         14830 => x"72",
         14831 => x"50",
         14832 => x"6d",
         14833 => x"72",
         14834 => x"6e",
         14835 => x"72",
         14836 => x"2e",
         14837 => x"54",
         14838 => x"6d",
         14839 => x"20",
         14840 => x"6e",
         14841 => x"6c",
         14842 => x"00",
         14843 => x"49",
         14844 => x"66",
         14845 => x"69",
         14846 => x"20",
         14847 => x"6f",
         14848 => x"00",
         14849 => x"46",
         14850 => x"20",
         14851 => x"6c",
         14852 => x"65",
         14853 => x"54",
         14854 => x"6f",
         14855 => x"20",
         14856 => x"72",
         14857 => x"6f",
         14858 => x"61",
         14859 => x"6c",
         14860 => x"2e",
         14861 => x"46",
         14862 => x"61",
         14863 => x"62",
         14864 => x"65",
         14865 => x"4e",
         14866 => x"6f",
         14867 => x"74",
         14868 => x"65",
         14869 => x"6c",
         14870 => x"73",
         14871 => x"20",
         14872 => x"6e",
         14873 => x"6e",
         14874 => x"73",
         14875 => x"44",
         14876 => x"20",
         14877 => x"20",
         14878 => x"62",
         14879 => x"2e",
         14880 => x"44",
         14881 => x"65",
         14882 => x"6d",
         14883 => x"20",
         14884 => x"69",
         14885 => x"6c",
         14886 => x"00",
         14887 => x"53",
         14888 => x"73",
         14889 => x"69",
         14890 => x"70",
         14891 => x"65",
         14892 => x"64",
         14893 => x"46",
         14894 => x"20",
         14895 => x"64",
         14896 => x"69",
         14897 => x"6c",
         14898 => x"00",
         14899 => x"46",
         14900 => x"20",
         14901 => x"65",
         14902 => x"20",
         14903 => x"73",
         14904 => x"00",
         14905 => x"41",
         14906 => x"73",
         14907 => x"65",
         14908 => x"64",
         14909 => x"49",
         14910 => x"6c",
         14911 => x"66",
         14912 => x"6e",
         14913 => x"2e",
         14914 => x"4e",
         14915 => x"61",
         14916 => x"66",
         14917 => x"64",
         14918 => x"4e",
         14919 => x"69",
         14920 => x"66",
         14921 => x"64",
         14922 => x"44",
         14923 => x"20",
         14924 => x"20",
         14925 => x"64",
         14926 => x"49",
         14927 => x"72",
         14928 => x"20",
         14929 => x"6f",
         14930 => x"44",
         14931 => x"20",
         14932 => x"6f",
         14933 => x"53",
         14934 => x"65",
         14935 => x"00",
         14936 => x"0a",
         14937 => x"20",
         14938 => x"65",
         14939 => x"73",
         14940 => x"20",
         14941 => x"20",
         14942 => x"65",
         14943 => x"65",
         14944 => x"00",
         14945 => x"72",
         14946 => x"00",
         14947 => x"25",
         14948 => x"58",
         14949 => x"3a",
         14950 => x"25",
         14951 => x"00",
         14952 => x"20",
         14953 => x"7c",
         14954 => x"20",
         14955 => x"25",
         14956 => x"00",
         14957 => x"20",
         14958 => x"20",
         14959 => x"00",
         14960 => x"7a",
         14961 => x"2a",
         14962 => x"73",
         14963 => x"32",
         14964 => x"37",
         14965 => x"32",
         14966 => x"76",
         14967 => x"32",
         14968 => x"20",
         14969 => x"2c",
         14970 => x"76",
         14971 => x"32",
         14972 => x"25",
         14973 => x"73",
         14974 => x"0a",
         14975 => x"4f",
         14976 => x"20",
         14977 => x"42",
         14978 => x"20",
         14979 => x"72",
         14980 => x"20",
         14981 => x"20",
         14982 => x"20",
         14983 => x"20",
         14984 => x"30",
         14985 => x"0a",
         14986 => x"20",
         14987 => x"41",
         14988 => x"41",
         14989 => x"65",
         14990 => x"20",
         14991 => x"20",
         14992 => x"20",
         14993 => x"20",
         14994 => x"30",
         14995 => x"0a",
         14996 => x"5a",
         14997 => x"49",
         14998 => x"72",
         14999 => x"74",
         15000 => x"6e",
         15001 => x"72",
         15002 => x"55",
         15003 => x"31",
         15004 => x"20",
         15005 => x"65",
         15006 => x"70",
         15007 => x"55",
         15008 => x"31",
         15009 => x"20",
         15010 => x"65",
         15011 => x"70",
         15012 => x"55",
         15013 => x"30",
         15014 => x"20",
         15015 => x"65",
         15016 => x"70",
         15017 => x"55",
         15018 => x"30",
         15019 => x"20",
         15020 => x"65",
         15021 => x"70",
         15022 => x"49",
         15023 => x"4c",
         15024 => x"20",
         15025 => x"65",
         15026 => x"70",
         15027 => x"49",
         15028 => x"4c",
         15029 => x"20",
         15030 => x"65",
         15031 => x"70",
         15032 => x"50",
         15033 => x"69",
         15034 => x"72",
         15035 => x"74",
         15036 => x"54",
         15037 => x"72",
         15038 => x"74",
         15039 => x"75",
         15040 => x"53",
         15041 => x"69",
         15042 => x"75",
         15043 => x"69",
         15044 => x"2e",
         15045 => x"45",
         15046 => x"6c",
         15047 => x"20",
         15048 => x"65",
         15049 => x"2e",
         15050 => x"61",
         15051 => x"65",
         15052 => x"2e",
         15053 => x"00",
         15054 => x"7a",
         15055 => x"7a",
         15056 => x"68",
         15057 => x"46",
         15058 => x"65",
         15059 => x"6f",
         15060 => x"69",
         15061 => x"6c",
         15062 => x"20",
         15063 => x"63",
         15064 => x"20",
         15065 => x"70",
         15066 => x"73",
         15067 => x"6e",
         15068 => x"6d",
         15069 => x"61",
         15070 => x"2e",
         15071 => x"2a",
         15072 => x"25",
         15073 => x"25",
         15074 => x"30",
         15075 => x"42",
         15076 => x"63",
         15077 => x"61",
         15078 => x"00",
         15079 => x"5a",
         15080 => x"62",
         15081 => x"25",
         15082 => x"25",
         15083 => x"73",
         15084 => x"00",
         15085 => x"43",
         15086 => x"20",
         15087 => x"6f",
         15088 => x"6e",
         15089 => x"2e",
         15090 => x"52",
         15091 => x"61",
         15092 => x"6e",
         15093 => x"70",
         15094 => x"63",
         15095 => x"6f",
         15096 => x"2e",
         15097 => x"43",
         15098 => x"69",
         15099 => x"63",
         15100 => x"20",
         15101 => x"30",
         15102 => x"20",
         15103 => x"0a",
         15104 => x"43",
         15105 => x"20",
         15106 => x"75",
         15107 => x"64",
         15108 => x"64",
         15109 => x"25",
         15110 => x"0a",
         15111 => x"45",
         15112 => x"75",
         15113 => x"67",
         15114 => x"64",
         15115 => x"20",
         15116 => x"6c",
         15117 => x"2e",
         15118 => x"25",
         15119 => x"58",
         15120 => x"38",
         15121 => x"00",
         15122 => x"25",
         15123 => x"58",
         15124 => x"34",
         15125 => x"43",
         15126 => x"61",
         15127 => x"67",
         15128 => x"00",
         15129 => x"25",
         15130 => x"78",
         15131 => x"38",
         15132 => x"3e",
         15133 => x"6c",
         15134 => x"30",
         15135 => x"0a",
         15136 => x"43",
         15137 => x"69",
         15138 => x"2e",
         15139 => x"25",
         15140 => x"58",
         15141 => x"32",
         15142 => x"43",
         15143 => x"72",
         15144 => x"2e",
         15145 => x"00",
         15146 => x"44",
         15147 => x"20",
         15148 => x"6f",
         15149 => x"0a",
         15150 => x"70",
         15151 => x"65",
         15152 => x"25",
         15153 => x"25",
         15154 => x"73",
         15155 => x"4d",
         15156 => x"72",
         15157 => x"78",
         15158 => x"73",
         15159 => x"2c",
         15160 => x"6e",
         15161 => x"20",
         15162 => x"63",
         15163 => x"20",
         15164 => x"6d",
         15165 => x"2e",
         15166 => x"3f",
         15167 => x"25",
         15168 => x"64",
         15169 => x"20",
         15170 => x"25",
         15171 => x"64",
         15172 => x"25",
         15173 => x"53",
         15174 => x"43",
         15175 => x"69",
         15176 => x"61",
         15177 => x"6e",
         15178 => x"3a",
         15179 => x"76",
         15180 => x"73",
         15181 => x"70",
         15182 => x"65",
         15183 => x"64",
         15184 => x"41",
         15185 => x"65",
         15186 => x"73",
         15187 => x"20",
         15188 => x"43",
         15189 => x"52",
         15190 => x"74",
         15191 => x"63",
         15192 => x"20",
         15193 => x"72",
         15194 => x"20",
         15195 => x"30",
         15196 => x"00",
         15197 => x"20",
         15198 => x"43",
         15199 => x"4d",
         15200 => x"72",
         15201 => x"74",
         15202 => x"20",
         15203 => x"72",
         15204 => x"20",
         15205 => x"30",
         15206 => x"00",
         15207 => x"20",
         15208 => x"53",
         15209 => x"6b",
         15210 => x"61",
         15211 => x"41",
         15212 => x"65",
         15213 => x"20",
         15214 => x"20",
         15215 => x"30",
         15216 => x"00",
         15217 => x"4d",
         15218 => x"3a",
         15219 => x"20",
         15220 => x"5a",
         15221 => x"49",
         15222 => x"20",
         15223 => x"20",
         15224 => x"20",
         15225 => x"20",
         15226 => x"20",
         15227 => x"30",
         15228 => x"00",
         15229 => x"20",
         15230 => x"53",
         15231 => x"65",
         15232 => x"6c",
         15233 => x"20",
         15234 => x"71",
         15235 => x"20",
         15236 => x"20",
         15237 => x"64",
         15238 => x"34",
         15239 => x"7a",
         15240 => x"20",
         15241 => x"57",
         15242 => x"62",
         15243 => x"20",
         15244 => x"41",
         15245 => x"6c",
         15246 => x"20",
         15247 => x"71",
         15248 => x"64",
         15249 => x"34",
         15250 => x"7a",
         15251 => x"20",
         15252 => x"53",
         15253 => x"4d",
         15254 => x"6f",
         15255 => x"46",
         15256 => x"20",
         15257 => x"20",
         15258 => x"20",
         15259 => x"64",
         15260 => x"34",
         15261 => x"7a",
         15262 => x"20",
         15263 => x"53",
         15264 => x"20",
         15265 => x"50",
         15266 => x"20",
         15267 => x"49",
         15268 => x"4c",
         15269 => x"20",
         15270 => x"57",
         15271 => x"32",
         15272 => x"20",
         15273 => x"57",
         15274 => x"42",
         15275 => x"20",
         15276 => x"00",
         15277 => x"20",
         15278 => x"49",
         15279 => x"20",
         15280 => x"4c",
         15281 => x"68",
         15282 => x"65",
         15283 => x"25",
         15284 => x"29",
         15285 => x"20",
         15286 => x"54",
         15287 => x"52",
         15288 => x"20",
         15289 => x"69",
         15290 => x"73",
         15291 => x"25",
         15292 => x"29",
         15293 => x"20",
         15294 => x"53",
         15295 => x"41",
         15296 => x"20",
         15297 => x"65",
         15298 => x"65",
         15299 => x"25",
         15300 => x"29",
         15301 => x"20",
         15302 => x"52",
         15303 => x"20",
         15304 => x"20",
         15305 => x"30",
         15306 => x"25",
         15307 => x"29",
         15308 => x"20",
         15309 => x"42",
         15310 => x"20",
         15311 => x"20",
         15312 => x"30",
         15313 => x"25",
         15314 => x"29",
         15315 => x"20",
         15316 => x"49",
         15317 => x"20",
         15318 => x"4d",
         15319 => x"30",
         15320 => x"25",
         15321 => x"29",
         15322 => x"20",
         15323 => x"53",
         15324 => x"4d",
         15325 => x"20",
         15326 => x"30",
         15327 => x"25",
         15328 => x"29",
         15329 => x"20",
         15330 => x"57",
         15331 => x"44",
         15332 => x"20",
         15333 => x"30",
         15334 => x"25",
         15335 => x"29",
         15336 => x"20",
         15337 => x"6f",
         15338 => x"6f",
         15339 => x"6f",
         15340 => x"67",
         15341 => x"55",
         15342 => x"6f",
         15343 => x"45",
         15344 => x"00",
         15345 => x"53",
         15346 => x"6c",
         15347 => x"4d",
         15348 => x"75",
         15349 => x"46",
         15350 => x"00",
         15351 => x"45",
         15352 => x"00",
         15353 => x"01",
         15354 => x"00",
         15355 => x"00",
         15356 => x"01",
         15357 => x"00",
         15358 => x"00",
         15359 => x"01",
         15360 => x"00",
         15361 => x"00",
         15362 => x"01",
         15363 => x"00",
         15364 => x"00",
         15365 => x"01",
         15366 => x"00",
         15367 => x"00",
         15368 => x"01",
         15369 => x"00",
         15370 => x"00",
         15371 => x"01",
         15372 => x"00",
         15373 => x"00",
         15374 => x"01",
         15375 => x"00",
         15376 => x"00",
         15377 => x"01",
         15378 => x"00",
         15379 => x"00",
         15380 => x"01",
         15381 => x"00",
         15382 => x"00",
         15383 => x"01",
         15384 => x"00",
         15385 => x"00",
         15386 => x"04",
         15387 => x"00",
         15388 => x"00",
         15389 => x"04",
         15390 => x"00",
         15391 => x"00",
         15392 => x"04",
         15393 => x"00",
         15394 => x"00",
         15395 => x"03",
         15396 => x"00",
         15397 => x"00",
         15398 => x"04",
         15399 => x"00",
         15400 => x"00",
         15401 => x"04",
         15402 => x"00",
         15403 => x"00",
         15404 => x"04",
         15405 => x"00",
         15406 => x"00",
         15407 => x"03",
         15408 => x"00",
         15409 => x"00",
         15410 => x"03",
         15411 => x"00",
         15412 => x"00",
         15413 => x"03",
         15414 => x"00",
         15415 => x"00",
         15416 => x"03",
         15417 => x"00",
         15418 => x"1b",
         15419 => x"1b",
         15420 => x"1b",
         15421 => x"1b",
         15422 => x"1b",
         15423 => x"1b",
         15424 => x"1b",
         15425 => x"1b",
         15426 => x"1b",
         15427 => x"1b",
         15428 => x"1b",
         15429 => x"10",
         15430 => x"0e",
         15431 => x"0d",
         15432 => x"0b",
         15433 => x"08",
         15434 => x"06",
         15435 => x"05",
         15436 => x"04",
         15437 => x"03",
         15438 => x"02",
         15439 => x"01",
         15440 => x"48",
         15441 => x"6f",
         15442 => x"68",
         15443 => x"3a",
         15444 => x"6c",
         15445 => x"43",
         15446 => x"6f",
         15447 => x"70",
         15448 => x"63",
         15449 => x"74",
         15450 => x"69",
         15451 => x"72",
         15452 => x"69",
         15453 => x"20",
         15454 => x"61",
         15455 => x"6e",
         15456 => x"68",
         15457 => x"6f",
         15458 => x"68",
         15459 => x"00",
         15460 => x"21",
         15461 => x"48",
         15462 => x"6f",
         15463 => x"62",
         15464 => x"65",
         15465 => x"30",
         15466 => x"0a",
         15467 => x"25",
         15468 => x"75",
         15469 => x"73",
         15470 => x"46",
         15471 => x"65",
         15472 => x"6f",
         15473 => x"73",
         15474 => x"74",
         15475 => x"68",
         15476 => x"6f",
         15477 => x"66",
         15478 => x"20",
         15479 => x"45",
         15480 => x"00",
         15481 => x"3e",
         15482 => x"00",
         15483 => x"1b",
         15484 => x"00",
         15485 => x"1b",
         15486 => x"1b",
         15487 => x"1b",
         15488 => x"1b",
         15489 => x"1b",
         15490 => x"7e",
         15491 => x"1b",
         15492 => x"7e",
         15493 => x"1b",
         15494 => x"7e",
         15495 => x"1b",
         15496 => x"7e",
         15497 => x"1b",
         15498 => x"7e",
         15499 => x"1b",
         15500 => x"7e",
         15501 => x"1b",
         15502 => x"7e",
         15503 => x"1b",
         15504 => x"7e",
         15505 => x"1b",
         15506 => x"7e",
         15507 => x"1b",
         15508 => x"7e",
         15509 => x"1b",
         15510 => x"00",
         15511 => x"1b",
         15512 => x"00",
         15513 => x"1b",
         15514 => x"1b",
         15515 => x"00",
         15516 => x"1b",
         15517 => x"00",
         15518 => x"58",
         15519 => x"2c",
         15520 => x"25",
         15521 => x"64",
         15522 => x"2c",
         15523 => x"25",
         15524 => x"00",
         15525 => x"44",
         15526 => x"2d",
         15527 => x"25",
         15528 => x"63",
         15529 => x"2c",
         15530 => x"25",
         15531 => x"25",
         15532 => x"4b",
         15533 => x"3a",
         15534 => x"25",
         15535 => x"2c",
         15536 => x"25",
         15537 => x"64",
         15538 => x"52",
         15539 => x"52",
         15540 => x"72",
         15541 => x"75",
         15542 => x"72",
         15543 => x"55",
         15544 => x"30",
         15545 => x"25",
         15546 => x"00",
         15547 => x"44",
         15548 => x"30",
         15549 => x"25",
         15550 => x"00",
         15551 => x"48",
         15552 => x"30",
         15553 => x"00",
         15554 => x"4e",
         15555 => x"65",
         15556 => x"64",
         15557 => x"6e",
         15558 => x"00",
         15559 => x"53",
         15560 => x"22",
         15561 => x"3e",
         15562 => x"00",
         15563 => x"2b",
         15564 => x"5b",
         15565 => x"46",
         15566 => x"46",
         15567 => x"32",
         15568 => x"eb",
         15569 => x"53",
         15570 => x"35",
         15571 => x"4e",
         15572 => x"41",
         15573 => x"20",
         15574 => x"41",
         15575 => x"20",
         15576 => x"4e",
         15577 => x"41",
         15578 => x"20",
         15579 => x"41",
         15580 => x"20",
         15581 => x"00",
         15582 => x"00",
         15583 => x"00",
         15584 => x"00",
         15585 => x"01",
         15586 => x"09",
         15587 => x"14",
         15588 => x"1e",
         15589 => x"80",
         15590 => x"8e",
         15591 => x"45",
         15592 => x"49",
         15593 => x"90",
         15594 => x"99",
         15595 => x"59",
         15596 => x"9c",
         15597 => x"41",
         15598 => x"a5",
         15599 => x"a8",
         15600 => x"ac",
         15601 => x"b0",
         15602 => x"b4",
         15603 => x"b8",
         15604 => x"bc",
         15605 => x"c0",
         15606 => x"c4",
         15607 => x"c8",
         15608 => x"cc",
         15609 => x"d0",
         15610 => x"d4",
         15611 => x"d8",
         15612 => x"dc",
         15613 => x"e0",
         15614 => x"e4",
         15615 => x"e8",
         15616 => x"ec",
         15617 => x"f0",
         15618 => x"f4",
         15619 => x"f8",
         15620 => x"fc",
         15621 => x"2b",
         15622 => x"3d",
         15623 => x"5c",
         15624 => x"3c",
         15625 => x"7f",
         15626 => x"00",
         15627 => x"00",
         15628 => x"01",
         15629 => x"00",
         15630 => x"00",
         15631 => x"00",
         15632 => x"00",
         15633 => x"00",
         15634 => x"00",
         15635 => x"00",
         15636 => x"00",
         15637 => x"00",
         15638 => x"00",
         15639 => x"00",
         15640 => x"00",
         15641 => x"00",
         15642 => x"00",
         15643 => x"00",
         15644 => x"00",
         15645 => x"00",
         15646 => x"00",
         15647 => x"00",
         15648 => x"00",
         15649 => x"20",
         15650 => x"00",
         15651 => x"00",
         15652 => x"00",
         15653 => x"00",
         15654 => x"00",
         15655 => x"00",
         15656 => x"00",
         15657 => x"00",
         15658 => x"25",
         15659 => x"25",
         15660 => x"25",
         15661 => x"25",
         15662 => x"25",
         15663 => x"25",
         15664 => x"25",
         15665 => x"25",
         15666 => x"25",
         15667 => x"25",
         15668 => x"25",
         15669 => x"25",
         15670 => x"25",
         15671 => x"25",
         15672 => x"25",
         15673 => x"25",
         15674 => x"25",
         15675 => x"25",
         15676 => x"25",
         15677 => x"25",
         15678 => x"25",
         15679 => x"25",
         15680 => x"25",
         15681 => x"25",
         15682 => x"03",
         15683 => x"03",
         15684 => x"03",
         15685 => x"00",
         15686 => x"03",
         15687 => x"03",
         15688 => x"22",
         15689 => x"03",
         15690 => x"22",
         15691 => x"22",
         15692 => x"23",
         15693 => x"00",
         15694 => x"00",
         15695 => x"00",
         15696 => x"20",
         15697 => x"25",
         15698 => x"00",
         15699 => x"00",
         15700 => x"00",
         15701 => x"00",
         15702 => x"01",
         15703 => x"01",
         15704 => x"01",
         15705 => x"01",
         15706 => x"01",
         15707 => x"01",
         15708 => x"00",
         15709 => x"01",
         15710 => x"01",
         15711 => x"01",
         15712 => x"01",
         15713 => x"01",
         15714 => x"01",
         15715 => x"01",
         15716 => x"01",
         15717 => x"01",
         15718 => x"01",
         15719 => x"01",
         15720 => x"01",
         15721 => x"01",
         15722 => x"01",
         15723 => x"01",
         15724 => x"01",
         15725 => x"01",
         15726 => x"01",
         15727 => x"01",
         15728 => x"01",
         15729 => x"01",
         15730 => x"01",
         15731 => x"01",
         15732 => x"01",
         15733 => x"01",
         15734 => x"01",
         15735 => x"01",
         15736 => x"01",
         15737 => x"01",
         15738 => x"01",
         15739 => x"01",
         15740 => x"01",
         15741 => x"01",
         15742 => x"01",
         15743 => x"01",
         15744 => x"01",
         15745 => x"01",
         15746 => x"01",
         15747 => x"01",
         15748 => x"01",
         15749 => x"01",
         15750 => x"01",
         15751 => x"00",
         15752 => x"01",
         15753 => x"01",
         15754 => x"02",
         15755 => x"02",
         15756 => x"2c",
         15757 => x"02",
         15758 => x"2c",
         15759 => x"02",
         15760 => x"02",
         15761 => x"01",
         15762 => x"00",
         15763 => x"01",
         15764 => x"01",
         15765 => x"02",
         15766 => x"02",
         15767 => x"02",
         15768 => x"02",
         15769 => x"01",
         15770 => x"02",
         15771 => x"02",
         15772 => x"02",
         15773 => x"01",
         15774 => x"02",
         15775 => x"02",
         15776 => x"02",
         15777 => x"02",
         15778 => x"01",
         15779 => x"02",
         15780 => x"02",
         15781 => x"02",
         15782 => x"02",
         15783 => x"02",
         15784 => x"02",
         15785 => x"01",
         15786 => x"02",
         15787 => x"02",
         15788 => x"02",
         15789 => x"01",
         15790 => x"01",
         15791 => x"02",
         15792 => x"02",
         15793 => x"02",
         15794 => x"01",
         15795 => x"00",
         15796 => x"03",
         15797 => x"03",
         15798 => x"03",
         15799 => x"03",
         15800 => x"03",
         15801 => x"03",
         15802 => x"03",
         15803 => x"03",
         15804 => x"03",
         15805 => x"03",
         15806 => x"03",
         15807 => x"01",
         15808 => x"00",
         15809 => x"03",
         15810 => x"03",
         15811 => x"03",
         15812 => x"03",
         15813 => x"03",
         15814 => x"03",
         15815 => x"07",
         15816 => x"01",
         15817 => x"01",
         15818 => x"01",
         15819 => x"00",
         15820 => x"04",
         15821 => x"05",
         15822 => x"00",
         15823 => x"1d",
         15824 => x"2c",
         15825 => x"01",
         15826 => x"01",
         15827 => x"06",
         15828 => x"06",
         15829 => x"06",
         15830 => x"06",
         15831 => x"06",
         15832 => x"00",
         15833 => x"1f",
         15834 => x"1f",
         15835 => x"1f",
         15836 => x"1f",
         15837 => x"1f",
         15838 => x"1f",
         15839 => x"1f",
         15840 => x"1f",
         15841 => x"1f",
         15842 => x"1f",
         15843 => x"1f",
         15844 => x"1f",
         15845 => x"1f",
         15846 => x"1f",
         15847 => x"1f",
         15848 => x"1f",
         15849 => x"1f",
         15850 => x"1f",
         15851 => x"1f",
         15852 => x"1f",
         15853 => x"06",
         15854 => x"06",
         15855 => x"00",
         15856 => x"1f",
         15857 => x"1f",
         15858 => x"00",
         15859 => x"21",
         15860 => x"21",
         15861 => x"21",
         15862 => x"05",
         15863 => x"04",
         15864 => x"01",
         15865 => x"01",
         15866 => x"01",
         15867 => x"01",
         15868 => x"08",
         15869 => x"03",
         15870 => x"00",
         15871 => x"00",
         15872 => x"01",
         15873 => x"00",
         15874 => x"00",
         15875 => x"00",
         15876 => x"01",
         15877 => x"00",
         15878 => x"00",
         15879 => x"00",
         15880 => x"01",
         15881 => x"00",
         15882 => x"00",
         15883 => x"00",
         15884 => x"01",
         15885 => x"00",
         15886 => x"00",
         15887 => x"00",
         15888 => x"01",
         15889 => x"00",
         15890 => x"00",
         15891 => x"00",
         15892 => x"01",
         15893 => x"00",
         15894 => x"00",
         15895 => x"00",
         15896 => x"01",
         15897 => x"00",
         15898 => x"00",
         15899 => x"00",
         15900 => x"01",
         15901 => x"00",
         15902 => x"00",
         15903 => x"00",
         15904 => x"01",
         15905 => x"00",
         15906 => x"00",
         15907 => x"00",
         15908 => x"01",
         15909 => x"00",
         15910 => x"00",
         15911 => x"00",
         15912 => x"01",
         15913 => x"00",
         15914 => x"00",
         15915 => x"00",
         15916 => x"01",
         15917 => x"00",
         15918 => x"00",
         15919 => x"00",
         15920 => x"01",
         15921 => x"00",
         15922 => x"00",
         15923 => x"00",
         15924 => x"01",
         15925 => x"00",
         15926 => x"00",
         15927 => x"00",
         15928 => x"01",
         15929 => x"00",
         15930 => x"00",
         15931 => x"00",
         15932 => x"01",
         15933 => x"00",
         15934 => x"00",
         15935 => x"00",
         15936 => x"01",
         15937 => x"00",
         15938 => x"00",
         15939 => x"00",
         15940 => x"01",
         15941 => x"00",
         15942 => x"00",
         15943 => x"00",
         15944 => x"01",
         15945 => x"00",
         15946 => x"00",
         15947 => x"00",
         15948 => x"01",
         15949 => x"00",
         15950 => x"00",
         15951 => x"00",
         15952 => x"01",
         15953 => x"00",
         15954 => x"00",
         15955 => x"00",
         15956 => x"01",
         15957 => x"00",
         15958 => x"00",
         15959 => x"00",
         15960 => x"01",
         15961 => x"00",
         15962 => x"00",
         15963 => x"00",
         15964 => x"01",
         15965 => x"00",
         15966 => x"00",
         15967 => x"00",
         15968 => x"01",
         15969 => x"00",
         15970 => x"00",
         15971 => x"00",
         15972 => x"01",
         15973 => x"00",
         15974 => x"00",
         15975 => x"00",
         15976 => x"01",
         15977 => x"00",
         15978 => x"00",
         15979 => x"00",
         15980 => x"01",
         15981 => x"00",
         15982 => x"00",
         15983 => x"00",
         15984 => x"00",
         15985 => x"00",
         15986 => x"00",
         15987 => x"00",
         15988 => x"00",
         15989 => x"00",
         15990 => x"00",
         15991 => x"00",
         15992 => x"01",
         15993 => x"01",
         15994 => x"00",
         15995 => x"00",
         15996 => x"00",
         15997 => x"00",
         15998 => x"05",
         15999 => x"05",
         16000 => x"05",
         16001 => x"00",
         16002 => x"01",
         16003 => x"01",
         16004 => x"01",
         16005 => x"01",
         16006 => x"00",
         16007 => x"00",
         16008 => x"00",
         16009 => x"00",
         16010 => x"00",
         16011 => x"00",
         16012 => x"00",
         16013 => x"00",
         16014 => x"00",
         16015 => x"00",
         16016 => x"00",
         16017 => x"00",
         16018 => x"00",
         16019 => x"00",
         16020 => x"00",
         16021 => x"00",
         16022 => x"00",
         16023 => x"00",
         16024 => x"00",
         16025 => x"00",
         16026 => x"00",
         16027 => x"00",
         16028 => x"00",
         16029 => x"00",
         16030 => x"00",
         16031 => x"01",
         16032 => x"00",
         16033 => x"01",
         16034 => x"00",
         16035 => x"02",
         16036 => x"00",
         16037 => x"1b",
         16038 => x"f0",
         16039 => x"79",
         16040 => x"5d",
         16041 => x"71",
         16042 => x"75",
         16043 => x"69",
         16044 => x"6d",
         16045 => x"61",
         16046 => x"65",
         16047 => x"31",
         16048 => x"35",
         16049 => x"5c",
         16050 => x"30",
         16051 => x"f6",
         16052 => x"f1",
         16053 => x"08",
         16054 => x"f0",
         16055 => x"80",
         16056 => x"84",
         16057 => x"1b",
         16058 => x"f0",
         16059 => x"59",
         16060 => x"5d",
         16061 => x"51",
         16062 => x"55",
         16063 => x"49",
         16064 => x"4d",
         16065 => x"41",
         16066 => x"45",
         16067 => x"31",
         16068 => x"35",
         16069 => x"5c",
         16070 => x"30",
         16071 => x"f6",
         16072 => x"f1",
         16073 => x"08",
         16074 => x"f0",
         16075 => x"80",
         16076 => x"84",
         16077 => x"1b",
         16078 => x"f0",
         16079 => x"59",
         16080 => x"7d",
         16081 => x"51",
         16082 => x"55",
         16083 => x"49",
         16084 => x"4d",
         16085 => x"41",
         16086 => x"45",
         16087 => x"21",
         16088 => x"25",
         16089 => x"7c",
         16090 => x"20",
         16091 => x"f7",
         16092 => x"f9",
         16093 => x"fb",
         16094 => x"f0",
         16095 => x"85",
         16096 => x"89",
         16097 => x"1b",
         16098 => x"f0",
         16099 => x"19",
         16100 => x"1d",
         16101 => x"11",
         16102 => x"15",
         16103 => x"09",
         16104 => x"0d",
         16105 => x"01",
         16106 => x"05",
         16107 => x"f0",
         16108 => x"f0",
         16109 => x"f0",
         16110 => x"f0",
         16111 => x"f0",
         16112 => x"f0",
         16113 => x"f0",
         16114 => x"f0",
         16115 => x"80",
         16116 => x"84",
         16117 => x"bf",
         16118 => x"f0",
         16119 => x"35",
         16120 => x"b7",
         16121 => x"7c",
         16122 => x"39",
         16123 => x"3d",
         16124 => x"1d",
         16125 => x"46",
         16126 => x"74",
         16127 => x"3f",
         16128 => x"7a",
         16129 => x"d3",
         16130 => x"9d",
         16131 => x"c6",
         16132 => x"c3",
         16133 => x"f0",
         16134 => x"f0",
         16135 => x"80",
         16136 => x"84",
         16137 => x"00",
         16138 => x"00",
         16139 => x"00",
         16140 => x"00",
         16141 => x"00",
         16142 => x"00",
         16143 => x"00",
         16144 => x"00",
         16145 => x"00",
         16146 => x"00",
         16147 => x"00",
         16148 => x"00",
         16149 => x"00",
         16150 => x"00",
         16151 => x"00",
         16152 => x"00",
         16153 => x"00",
         16154 => x"00",
         16155 => x"00",
         16156 => x"00",
         16157 => x"00",
         16158 => x"00",
         16159 => x"00",
         16160 => x"00",
         16161 => x"00",
         16162 => x"00",
         16163 => x"00",
         16164 => x"f8",
         16165 => x"00",
         16166 => x"f3",
         16167 => x"00",
         16168 => x"f4",
         16169 => x"00",
         16170 => x"f1",
         16171 => x"00",
         16172 => x"f2",
         16173 => x"00",
         16174 => x"80",
         16175 => x"00",
         16176 => x"81",
         16177 => x"00",
         16178 => x"82",
         16179 => x"00",
         16180 => x"83",
         16181 => x"00",
         16182 => x"84",
         16183 => x"00",
         16184 => x"85",
         16185 => x"00",
         16186 => x"86",
         16187 => x"00",
         16188 => x"87",
         16189 => x"00",
         16190 => x"88",
         16191 => x"00",
         16192 => x"89",
         16193 => x"00",
         16194 => x"f6",
         16195 => x"00",
         16196 => x"7f",
         16197 => x"00",
         16198 => x"f9",
         16199 => x"00",
         16200 => x"e0",
         16201 => x"00",
         16202 => x"e1",
         16203 => x"00",
         16204 => x"71",
         16205 => x"00",
         16206 => x"00",
         16207 => x"00",
         16208 => x"00",
         16209 => x"00",
         16210 => x"00",
         16211 => x"00",
         16212 => x"00",
         16213 => x"00",
         16214 => x"00",
         16215 => x"00",
         16216 => x"00",
         16217 => x"00",
         16218 => x"00",
         16219 => x"00",
         16220 => x"00",
         16221 => x"00",
         16222 => x"00",
         16223 => x"00",
         16224 => x"00",
         16225 => x"00",
         16226 => x"00",
         16227 => x"00",
         16228 => x"00",
         16229 => x"00",
         16230 => x"00",
         16231 => x"00",
         16232 => x"00",
         16233 => x"00",
         16234 => x"00",
         16235 => x"00",
         16236 => x"00",
         16237 => x"00",
         16238 => x"00",
         16239 => x"00",
         16240 => x"00",
         16241 => x"00",
         16242 => x"00",
         16243 => x"00",
         16244 => x"00",
         16245 => x"00",
         16246 => x"00",
         16247 => x"00",
         16248 => x"00",
         16249 => x"00",
         16250 => x"00",
         16251 => x"00",
         16252 => x"00",
         16253 => x"00",
         16254 => x"00",
         16255 => x"00",
         16256 => x"00",
         16257 => x"00",
         16258 => x"00",
         16259 => x"00",
         16260 => x"00",
         16261 => x"00",
         16262 => x"00",
         16263 => x"00",
         16264 => x"00",
         16265 => x"00",
         16266 => x"00",
         16267 => x"00",
         16268 => x"00",
         16269 => x"00",
         16270 => x"00",
         16271 => x"00",
         16272 => x"00",
         16273 => x"00",
         16274 => x"00",
         16275 => x"00",
         16276 => x"00",
         16277 => x"00",
         16278 => x"00",
         16279 => x"00",
         16280 => x"00",
         16281 => x"00",
         16282 => x"00",
         16283 => x"00",
         16284 => x"00",
         16285 => x"00",
         16286 => x"00",
         16287 => x"00",
         16288 => x"00",
         16289 => x"00",
         16290 => x"00",
         16291 => x"00",
         16292 => x"00",
         16293 => x"00",
         16294 => x"00",
         16295 => x"00",
         16296 => x"00",
         16297 => x"00",
         16298 => x"00",
         16299 => x"00",
         16300 => x"00",
         16301 => x"00",
         16302 => x"00",
         16303 => x"00",
         16304 => x"00",
         16305 => x"00",
         16306 => x"00",
         16307 => x"00",
         16308 => x"00",
         16309 => x"00",
         16310 => x"00",
         16311 => x"00",
         16312 => x"00",
         16313 => x"00",
         16314 => x"00",
         16315 => x"00",
         16316 => x"00",
         16317 => x"00",
         16318 => x"00",
         16319 => x"00",
         16320 => x"00",
         16321 => x"00",
         16322 => x"00",
         16323 => x"00",
         16324 => x"00",
         16325 => x"00",
         16326 => x"00",
         16327 => x"00",
         16328 => x"00",
         16329 => x"00",
         16330 => x"00",
         16331 => x"00",
         16332 => x"00",
         16333 => x"00",
         16334 => x"00",
         16335 => x"00",
         16336 => x"00",
         16337 => x"00",
         16338 => x"00",
         16339 => x"00",
         16340 => x"00",
         16341 => x"00",
         16342 => x"00",
         16343 => x"00",
         16344 => x"00",
         16345 => x"00",
         16346 => x"00",
         16347 => x"00",
         16348 => x"00",
         16349 => x"00",
         16350 => x"00",
         16351 => x"00",
         16352 => x"00",
         16353 => x"00",
         16354 => x"00",
         16355 => x"00",
         16356 => x"00",
         16357 => x"00",
         16358 => x"00",
         16359 => x"00",
         16360 => x"00",
         16361 => x"00",
         16362 => x"00",
         16363 => x"00",
         16364 => x"00",
         16365 => x"00",
         16366 => x"00",
         16367 => x"00",
         16368 => x"00",
         16369 => x"00",
         16370 => x"00",
         16371 => x"00",
         16372 => x"00",
         16373 => x"00",
         16374 => x"00",
         16375 => x"00",
         16376 => x"00",
         16377 => x"00",
         16378 => x"00",
         16379 => x"00",
         16380 => x"00",
         16381 => x"00",
         16382 => x"00",
         16383 => x"00",
         16384 => x"00",
         16385 => x"00",
         16386 => x"00",
         16387 => x"00",
         16388 => x"00",
         16389 => x"00",
         16390 => x"00",
         16391 => x"00",
         16392 => x"00",
         16393 => x"00",
         16394 => x"00",
         16395 => x"00",
         16396 => x"00",
         16397 => x"00",
         16398 => x"00",
         16399 => x"00",
         16400 => x"00",
         16401 => x"00",
         16402 => x"00",
         16403 => x"00",
         16404 => x"00",
         16405 => x"00",
         16406 => x"00",
         16407 => x"00",
         16408 => x"00",
         16409 => x"00",
         16410 => x"00",
         16411 => x"00",
         16412 => x"00",
         16413 => x"00",
         16414 => x"00",
         16415 => x"00",
         16416 => x"00",
         16417 => x"00",
         16418 => x"00",
         16419 => x"00",
         16420 => x"00",
         16421 => x"00",
         16422 => x"00",
         16423 => x"00",
         16424 => x"00",
         16425 => x"00",
         16426 => x"00",
         16427 => x"00",
         16428 => x"00",
         16429 => x"00",
         16430 => x"00",
         16431 => x"00",
         16432 => x"00",
         16433 => x"00",
         16434 => x"00",
         16435 => x"00",
         16436 => x"00",
         16437 => x"00",
         16438 => x"00",
         16439 => x"00",
         16440 => x"00",
         16441 => x"00",
         16442 => x"00",
         16443 => x"00",
         16444 => x"00",
         16445 => x"00",
         16446 => x"00",
         16447 => x"00",
         16448 => x"00",
         16449 => x"00",
         16450 => x"00",
         16451 => x"00",
         16452 => x"00",
         16453 => x"00",
         16454 => x"00",
         16455 => x"00",
         16456 => x"00",
         16457 => x"00",
         16458 => x"00",
         16459 => x"00",
         16460 => x"00",
         16461 => x"00",
         16462 => x"00",
         16463 => x"00",
         16464 => x"00",
         16465 => x"00",
         16466 => x"00",
         16467 => x"00",
         16468 => x"00",
         16469 => x"00",
         16470 => x"00",
         16471 => x"00",
         16472 => x"00",
         16473 => x"00",
         16474 => x"00",
         16475 => x"00",
         16476 => x"00",
         16477 => x"00",
         16478 => x"00",
         16479 => x"00",
         16480 => x"00",
         16481 => x"00",
         16482 => x"00",
         16483 => x"00",
         16484 => x"00",
         16485 => x"00",
         16486 => x"00",
         16487 => x"00",
         16488 => x"00",
         16489 => x"00",
         16490 => x"00",
         16491 => x"00",
         16492 => x"00",
         16493 => x"00",
         16494 => x"00",
         16495 => x"00",
         16496 => x"00",
         16497 => x"00",
         16498 => x"00",
         16499 => x"00",
         16500 => x"00",
         16501 => x"00",
         16502 => x"00",
         16503 => x"00",
         16504 => x"00",
         16505 => x"00",
         16506 => x"00",
         16507 => x"00",
         16508 => x"00",
         16509 => x"00",
         16510 => x"00",
         16511 => x"00",
         16512 => x"00",
         16513 => x"00",
         16514 => x"00",
         16515 => x"00",
         16516 => x"00",
         16517 => x"00",
         16518 => x"00",
         16519 => x"00",
         16520 => x"00",
         16521 => x"00",
         16522 => x"00",
         16523 => x"00",
         16524 => x"00",
         16525 => x"00",
         16526 => x"00",
         16527 => x"00",
         16528 => x"00",
         16529 => x"00",
         16530 => x"00",
         16531 => x"00",
         16532 => x"00",
         16533 => x"00",
         16534 => x"00",
         16535 => x"00",
         16536 => x"00",
         16537 => x"00",
         16538 => x"00",
         16539 => x"00",
         16540 => x"00",
         16541 => x"00",
         16542 => x"00",
         16543 => x"00",
         16544 => x"00",
         16545 => x"00",
         16546 => x"00",
         16547 => x"00",
         16548 => x"00",
         16549 => x"00",
         16550 => x"00",
         16551 => x"00",
         16552 => x"00",
         16553 => x"00",
         16554 => x"00",
         16555 => x"00",
         16556 => x"00",
         16557 => x"00",
         16558 => x"00",
         16559 => x"00",
         16560 => x"00",
         16561 => x"00",
         16562 => x"00",
         16563 => x"00",
         16564 => x"00",
         16565 => x"00",
         16566 => x"00",
         16567 => x"00",
         16568 => x"00",
         16569 => x"00",
         16570 => x"00",
         16571 => x"00",
         16572 => x"00",
         16573 => x"00",
         16574 => x"00",
         16575 => x"00",
         16576 => x"00",
         16577 => x"00",
         16578 => x"00",
         16579 => x"00",
         16580 => x"00",
         16581 => x"00",
         16582 => x"00",
         16583 => x"00",
         16584 => x"00",
         16585 => x"00",
         16586 => x"00",
         16587 => x"00",
         16588 => x"00",
         16589 => x"00",
         16590 => x"00",
         16591 => x"00",
         16592 => x"00",
         16593 => x"00",
         16594 => x"00",
         16595 => x"00",
         16596 => x"00",
         16597 => x"00",
         16598 => x"00",
         16599 => x"00",
         16600 => x"00",
         16601 => x"00",
         16602 => x"00",
         16603 => x"00",
         16604 => x"00",
         16605 => x"00",
         16606 => x"00",
         16607 => x"00",
         16608 => x"00",
         16609 => x"00",
         16610 => x"00",
         16611 => x"00",
         16612 => x"00",
         16613 => x"00",
         16614 => x"00",
         16615 => x"00",
         16616 => x"00",
         16617 => x"00",
         16618 => x"00",
         16619 => x"00",
         16620 => x"00",
         16621 => x"00",
         16622 => x"00",
         16623 => x"00",
         16624 => x"00",
         16625 => x"00",
         16626 => x"00",
         16627 => x"00",
         16628 => x"00",
         16629 => x"00",
         16630 => x"00",
         16631 => x"00",
         16632 => x"00",
         16633 => x"00",
         16634 => x"00",
         16635 => x"00",
         16636 => x"00",
         16637 => x"00",
         16638 => x"00",
         16639 => x"00",
         16640 => x"00",
         16641 => x"00",
         16642 => x"00",
         16643 => x"00",
         16644 => x"00",
         16645 => x"00",
         16646 => x"00",
         16647 => x"00",
         16648 => x"00",
         16649 => x"00",
         16650 => x"00",
         16651 => x"00",
         16652 => x"00",
         16653 => x"00",
         16654 => x"00",
         16655 => x"00",
         16656 => x"00",
         16657 => x"00",
         16658 => x"00",
         16659 => x"00",
         16660 => x"00",
         16661 => x"00",
         16662 => x"00",
         16663 => x"00",
         16664 => x"00",
         16665 => x"00",
         16666 => x"00",
         16667 => x"00",
         16668 => x"00",
         16669 => x"00",
         16670 => x"00",
         16671 => x"00",
         16672 => x"00",
         16673 => x"00",
         16674 => x"00",
         16675 => x"00",
         16676 => x"00",
         16677 => x"00",
         16678 => x"00",
         16679 => x"00",
         16680 => x"00",
         16681 => x"00",
         16682 => x"00",
         16683 => x"00",
         16684 => x"00",
         16685 => x"00",
         16686 => x"00",
         16687 => x"00",
         16688 => x"00",
         16689 => x"00",
         16690 => x"00",
         16691 => x"00",
         16692 => x"00",
         16693 => x"00",
         16694 => x"00",
         16695 => x"00",
         16696 => x"00",
         16697 => x"00",
         16698 => x"00",
         16699 => x"00",
         16700 => x"00",
         16701 => x"00",
         16702 => x"00",
         16703 => x"00",
         16704 => x"00",
         16705 => x"00",
         16706 => x"00",
         16707 => x"00",
         16708 => x"00",
         16709 => x"00",
         16710 => x"00",
         16711 => x"00",
         16712 => x"00",
         16713 => x"00",
         16714 => x"00",
         16715 => x"00",
         16716 => x"00",
         16717 => x"00",
         16718 => x"00",
         16719 => x"00",
         16720 => x"00",
         16721 => x"00",
         16722 => x"00",
         16723 => x"00",
         16724 => x"00",
         16725 => x"00",
         16726 => x"00",
         16727 => x"00",
         16728 => x"00",
         16729 => x"00",
         16730 => x"00",
         16731 => x"00",
         16732 => x"00",
         16733 => x"00",
         16734 => x"00",
         16735 => x"00",
         16736 => x"00",
         16737 => x"00",
         16738 => x"00",
         16739 => x"00",
         16740 => x"00",
         16741 => x"00",
         16742 => x"00",
         16743 => x"00",
         16744 => x"00",
         16745 => x"00",
         16746 => x"00",
         16747 => x"00",
         16748 => x"00",
         16749 => x"00",
         16750 => x"00",
         16751 => x"00",
         16752 => x"00",
         16753 => x"00",
         16754 => x"00",
         16755 => x"00",
         16756 => x"00",
         16757 => x"00",
         16758 => x"00",
         16759 => x"00",
         16760 => x"00",
         16761 => x"00",
         16762 => x"00",
         16763 => x"00",
         16764 => x"00",
         16765 => x"00",
         16766 => x"00",
         16767 => x"00",
         16768 => x"00",
         16769 => x"00",
         16770 => x"00",
         16771 => x"00",
         16772 => x"00",
         16773 => x"00",
         16774 => x"00",
         16775 => x"00",
         16776 => x"00",
         16777 => x"00",
         16778 => x"00",
         16779 => x"00",
         16780 => x"00",
         16781 => x"00",
         16782 => x"00",
         16783 => x"00",
         16784 => x"00",
         16785 => x"00",
         16786 => x"00",
         16787 => x"00",
         16788 => x"00",
         16789 => x"00",
         16790 => x"00",
         16791 => x"00",
         16792 => x"00",
         16793 => x"00",
         16794 => x"00",
         16795 => x"00",
         16796 => x"00",
         16797 => x"00",
         16798 => x"00",
         16799 => x"00",
         16800 => x"00",
         16801 => x"00",
         16802 => x"00",
         16803 => x"00",
         16804 => x"00",
         16805 => x"00",
         16806 => x"00",
         16807 => x"00",
         16808 => x"00",
         16809 => x"00",
         16810 => x"00",
         16811 => x"00",
         16812 => x"00",
         16813 => x"00",
         16814 => x"00",
         16815 => x"00",
         16816 => x"00",
         16817 => x"00",
         16818 => x"00",
         16819 => x"00",
         16820 => x"00",
         16821 => x"00",
         16822 => x"00",
         16823 => x"00",
         16824 => x"00",
         16825 => x"00",
         16826 => x"00",
         16827 => x"00",
         16828 => x"00",
         16829 => x"00",
         16830 => x"00",
         16831 => x"00",
         16832 => x"00",
         16833 => x"00",
         16834 => x"00",
         16835 => x"00",
         16836 => x"00",
         16837 => x"00",
         16838 => x"00",
         16839 => x"00",
         16840 => x"00",
         16841 => x"00",
         16842 => x"00",
         16843 => x"00",
         16844 => x"00",
         16845 => x"00",
         16846 => x"00",
         16847 => x"00",
         16848 => x"00",
         16849 => x"00",
         16850 => x"00",
         16851 => x"00",
         16852 => x"00",
         16853 => x"00",
         16854 => x"00",
         16855 => x"00",
         16856 => x"00",
         16857 => x"00",
         16858 => x"00",
         16859 => x"00",
         16860 => x"00",
         16861 => x"00",
         16862 => x"00",
         16863 => x"00",
         16864 => x"00",
         16865 => x"00",
         16866 => x"00",
         16867 => x"00",
         16868 => x"00",
         16869 => x"00",
         16870 => x"00",
         16871 => x"00",
         16872 => x"00",
         16873 => x"00",
         16874 => x"00",
         16875 => x"00",
         16876 => x"00",
         16877 => x"00",
         16878 => x"00",
         16879 => x"00",
         16880 => x"00",
         16881 => x"00",
         16882 => x"00",
         16883 => x"00",
         16884 => x"00",
         16885 => x"00",
         16886 => x"00",
         16887 => x"00",
         16888 => x"00",
         16889 => x"00",
         16890 => x"00",
         16891 => x"00",
         16892 => x"00",
         16893 => x"00",
         16894 => x"00",
         16895 => x"00",
         16896 => x"00",
         16897 => x"00",
         16898 => x"00",
         16899 => x"00",
         16900 => x"00",
         16901 => x"00",
         16902 => x"00",
         16903 => x"00",
         16904 => x"00",
         16905 => x"00",
         16906 => x"00",
         16907 => x"00",
         16908 => x"00",
         16909 => x"00",
         16910 => x"00",
         16911 => x"00",
         16912 => x"00",
         16913 => x"00",
         16914 => x"00",
         16915 => x"00",
         16916 => x"00",
         16917 => x"00",
         16918 => x"00",
         16919 => x"00",
         16920 => x"00",
         16921 => x"00",
         16922 => x"00",
         16923 => x"00",
         16924 => x"00",
         16925 => x"00",
         16926 => x"00",
         16927 => x"00",
         16928 => x"00",
         16929 => x"00",
         16930 => x"00",
         16931 => x"00",
         16932 => x"00",
         16933 => x"00",
         16934 => x"00",
         16935 => x"00",
         16936 => x"00",
         16937 => x"00",
         16938 => x"00",
         16939 => x"00",
         16940 => x"00",
         16941 => x"00",
         16942 => x"00",
         16943 => x"00",
         16944 => x"00",
         16945 => x"00",
         16946 => x"00",
         16947 => x"00",
         16948 => x"00",
         16949 => x"00",
         16950 => x"00",
         16951 => x"00",
         16952 => x"00",
         16953 => x"00",
         16954 => x"00",
         16955 => x"00",
         16956 => x"00",
         16957 => x"00",
         16958 => x"00",
         16959 => x"00",
         16960 => x"00",
         16961 => x"00",
         16962 => x"00",
         16963 => x"00",
         16964 => x"00",
         16965 => x"00",
         16966 => x"00",
         16967 => x"00",
         16968 => x"00",
         16969 => x"00",
         16970 => x"00",
         16971 => x"00",
         16972 => x"00",
         16973 => x"00",
         16974 => x"00",
         16975 => x"00",
         16976 => x"00",
         16977 => x"00",
         16978 => x"00",
         16979 => x"00",
         16980 => x"00",
         16981 => x"00",
         16982 => x"00",
         16983 => x"00",
         16984 => x"00",
         16985 => x"00",
         16986 => x"00",
         16987 => x"00",
         16988 => x"00",
         16989 => x"00",
         16990 => x"00",
         16991 => x"00",
         16992 => x"00",
         16993 => x"00",
         16994 => x"00",
         16995 => x"00",
         16996 => x"00",
         16997 => x"00",
         16998 => x"00",
         16999 => x"00",
         17000 => x"00",
         17001 => x"00",
         17002 => x"00",
         17003 => x"00",
         17004 => x"00",
         17005 => x"00",
         17006 => x"00",
         17007 => x"00",
         17008 => x"00",
         17009 => x"00",
         17010 => x"00",
         17011 => x"00",
         17012 => x"00",
         17013 => x"00",
         17014 => x"00",
         17015 => x"00",
         17016 => x"00",
         17017 => x"00",
         17018 => x"00",
         17019 => x"00",
         17020 => x"00",
         17021 => x"00",
         17022 => x"00",
         17023 => x"00",
         17024 => x"00",
         17025 => x"00",
         17026 => x"00",
         17027 => x"00",
         17028 => x"00",
         17029 => x"00",
         17030 => x"00",
         17031 => x"00",
         17032 => x"00",
         17033 => x"00",
         17034 => x"00",
         17035 => x"00",
         17036 => x"00",
         17037 => x"00",
         17038 => x"00",
         17039 => x"00",
         17040 => x"00",
         17041 => x"00",
         17042 => x"00",
         17043 => x"00",
         17044 => x"00",
         17045 => x"00",
         17046 => x"00",
         17047 => x"00",
         17048 => x"00",
         17049 => x"00",
         17050 => x"00",
         17051 => x"00",
         17052 => x"00",
         17053 => x"00",
         17054 => x"00",
         17055 => x"00",
         17056 => x"00",
         17057 => x"00",
         17058 => x"00",
         17059 => x"00",
         17060 => x"00",
         17061 => x"00",
         17062 => x"00",
         17063 => x"00",
         17064 => x"00",
         17065 => x"00",
         17066 => x"00",
         17067 => x"00",
         17068 => x"00",
         17069 => x"00",
         17070 => x"00",
         17071 => x"00",
         17072 => x"00",
         17073 => x"00",
         17074 => x"00",
         17075 => x"00",
         17076 => x"00",
         17077 => x"00",
         17078 => x"00",
         17079 => x"00",
         17080 => x"00",
         17081 => x"00",
         17082 => x"00",
         17083 => x"00",
         17084 => x"00",
         17085 => x"00",
         17086 => x"00",
         17087 => x"00",
         17088 => x"00",
         17089 => x"00",
         17090 => x"00",
         17091 => x"00",
         17092 => x"00",
         17093 => x"00",
         17094 => x"00",
         17095 => x"00",
         17096 => x"00",
         17097 => x"00",
         17098 => x"00",
         17099 => x"00",
         17100 => x"00",
         17101 => x"00",
         17102 => x"00",
         17103 => x"00",
         17104 => x"00",
         17105 => x"00",
         17106 => x"00",
         17107 => x"00",
         17108 => x"00",
         17109 => x"00",
         17110 => x"00",
         17111 => x"00",
         17112 => x"00",
         17113 => x"00",
         17114 => x"00",
         17115 => x"00",
         17116 => x"00",
         17117 => x"00",
         17118 => x"00",
         17119 => x"00",
         17120 => x"00",
         17121 => x"00",
         17122 => x"00",
         17123 => x"00",
         17124 => x"00",
         17125 => x"00",
         17126 => x"00",
         17127 => x"00",
         17128 => x"00",
         17129 => x"00",
         17130 => x"00",
         17131 => x"00",
         17132 => x"00",
         17133 => x"00",
         17134 => x"00",
         17135 => x"00",
         17136 => x"00",
         17137 => x"00",
         17138 => x"00",
         17139 => x"00",
         17140 => x"00",
         17141 => x"00",
         17142 => x"00",
         17143 => x"00",
         17144 => x"00",
         17145 => x"00",
         17146 => x"00",
         17147 => x"00",
         17148 => x"00",
         17149 => x"00",
         17150 => x"00",
         17151 => x"00",
         17152 => x"00",
         17153 => x"00",
         17154 => x"00",
         17155 => x"00",
         17156 => x"00",
         17157 => x"00",
         17158 => x"00",
         17159 => x"00",
         17160 => x"00",
         17161 => x"00",
         17162 => x"00",
         17163 => x"00",
         17164 => x"00",
         17165 => x"00",
         17166 => x"00",
         17167 => x"00",
         17168 => x"00",
         17169 => x"00",
         17170 => x"00",
         17171 => x"00",
         17172 => x"00",
         17173 => x"00",
         17174 => x"00",
         17175 => x"00",
         17176 => x"00",
         17177 => x"00",
         17178 => x"00",
         17179 => x"00",
         17180 => x"00",
         17181 => x"00",
         17182 => x"00",
         17183 => x"00",
         17184 => x"00",
         17185 => x"00",
         17186 => x"00",
         17187 => x"00",
         17188 => x"00",
         17189 => x"00",
         17190 => x"00",
         17191 => x"00",
         17192 => x"00",
         17193 => x"00",
         17194 => x"00",
         17195 => x"00",
         17196 => x"00",
         17197 => x"00",
         17198 => x"00",
         17199 => x"00",
         17200 => x"00",
         17201 => x"00",
         17202 => x"00",
         17203 => x"00",
         17204 => x"00",
         17205 => x"00",
         17206 => x"00",
         17207 => x"00",
         17208 => x"00",
         17209 => x"00",
         17210 => x"00",
         17211 => x"00",
         17212 => x"00",
         17213 => x"00",
         17214 => x"00",
         17215 => x"00",
         17216 => x"00",
         17217 => x"00",
         17218 => x"00",
         17219 => x"00",
         17220 => x"00",
         17221 => x"00",
         17222 => x"00",
         17223 => x"00",
         17224 => x"00",
         17225 => x"00",
         17226 => x"00",
         17227 => x"00",
         17228 => x"00",
         17229 => x"00",
         17230 => x"00",
         17231 => x"00",
         17232 => x"00",
         17233 => x"00",
         17234 => x"00",
         17235 => x"00",
         17236 => x"00",
         17237 => x"00",
         17238 => x"00",
         17239 => x"00",
         17240 => x"00",
         17241 => x"00",
         17242 => x"00",
         17243 => x"00",
         17244 => x"00",
         17245 => x"00",
         17246 => x"00",
         17247 => x"00",
         17248 => x"00",
         17249 => x"00",
         17250 => x"00",
         17251 => x"00",
         17252 => x"00",
         17253 => x"00",
         17254 => x"00",
         17255 => x"00",
         17256 => x"00",
         17257 => x"00",
         17258 => x"00",
         17259 => x"00",
         17260 => x"00",
         17261 => x"00",
         17262 => x"00",
         17263 => x"00",
         17264 => x"00",
         17265 => x"00",
         17266 => x"00",
         17267 => x"00",
         17268 => x"00",
         17269 => x"00",
         17270 => x"00",
         17271 => x"00",
         17272 => x"00",
         17273 => x"00",
         17274 => x"00",
         17275 => x"00",
         17276 => x"00",
         17277 => x"00",
         17278 => x"00",
         17279 => x"00",
         17280 => x"00",
         17281 => x"00",
         17282 => x"00",
         17283 => x"00",
         17284 => x"00",
         17285 => x"00",
         17286 => x"00",
         17287 => x"00",
         17288 => x"00",
         17289 => x"00",
         17290 => x"00",
         17291 => x"00",
         17292 => x"00",
         17293 => x"00",
         17294 => x"00",
         17295 => x"00",
         17296 => x"00",
         17297 => x"00",
         17298 => x"00",
         17299 => x"00",
         17300 => x"00",
         17301 => x"00",
         17302 => x"00",
         17303 => x"00",
         17304 => x"00",
         17305 => x"00",
         17306 => x"00",
         17307 => x"00",
         17308 => x"00",
         17309 => x"00",
         17310 => x"00",
         17311 => x"00",
         17312 => x"00",
         17313 => x"00",
         17314 => x"00",
         17315 => x"00",
         17316 => x"00",
         17317 => x"00",
         17318 => x"00",
         17319 => x"00",
         17320 => x"00",
         17321 => x"00",
         17322 => x"00",
         17323 => x"00",
         17324 => x"00",
         17325 => x"00",
         17326 => x"00",
         17327 => x"00",
         17328 => x"00",
         17329 => x"00",
         17330 => x"00",
         17331 => x"00",
         17332 => x"00",
         17333 => x"00",
         17334 => x"00",
         17335 => x"00",
         17336 => x"00",
         17337 => x"00",
         17338 => x"00",
         17339 => x"00",
         17340 => x"00",
         17341 => x"00",
         17342 => x"00",
         17343 => x"00",
         17344 => x"00",
         17345 => x"00",
         17346 => x"00",
         17347 => x"00",
         17348 => x"00",
         17349 => x"00",
         17350 => x"00",
         17351 => x"00",
         17352 => x"00",
         17353 => x"00",
         17354 => x"00",
         17355 => x"00",
         17356 => x"00",
         17357 => x"00",
         17358 => x"00",
         17359 => x"00",
         17360 => x"00",
         17361 => x"00",
         17362 => x"00",
         17363 => x"00",
         17364 => x"00",
         17365 => x"00",
         17366 => x"00",
         17367 => x"00",
         17368 => x"00",
         17369 => x"00",
         17370 => x"00",
         17371 => x"00",
         17372 => x"00",
         17373 => x"00",
         17374 => x"00",
         17375 => x"00",
         17376 => x"00",
         17377 => x"00",
         17378 => x"00",
         17379 => x"00",
         17380 => x"00",
         17381 => x"00",
         17382 => x"00",
         17383 => x"00",
         17384 => x"00",
         17385 => x"00",
         17386 => x"00",
         17387 => x"00",
         17388 => x"00",
         17389 => x"00",
         17390 => x"00",
         17391 => x"00",
         17392 => x"00",
         17393 => x"00",
         17394 => x"00",
         17395 => x"00",
         17396 => x"00",
         17397 => x"00",
         17398 => x"00",
         17399 => x"00",
         17400 => x"00",
         17401 => x"00",
         17402 => x"00",
         17403 => x"00",
         17404 => x"00",
         17405 => x"00",
         17406 => x"00",
         17407 => x"00",
         17408 => x"00",
         17409 => x"00",
         17410 => x"00",
         17411 => x"00",
         17412 => x"00",
         17413 => x"00",
         17414 => x"00",
         17415 => x"00",
         17416 => x"00",
         17417 => x"00",
         17418 => x"00",
         17419 => x"00",
         17420 => x"00",
         17421 => x"00",
         17422 => x"00",
         17423 => x"00",
         17424 => x"00",
         17425 => x"00",
         17426 => x"00",
         17427 => x"00",
         17428 => x"00",
         17429 => x"00",
         17430 => x"00",
         17431 => x"00",
         17432 => x"00",
         17433 => x"00",
         17434 => x"00",
         17435 => x"00",
         17436 => x"00",
         17437 => x"00",
         17438 => x"00",
         17439 => x"00",
         17440 => x"00",
         17441 => x"00",
         17442 => x"00",
         17443 => x"00",
         17444 => x"00",
         17445 => x"00",
         17446 => x"00",
         17447 => x"00",
         17448 => x"00",
         17449 => x"00",
         17450 => x"00",
         17451 => x"00",
         17452 => x"00",
         17453 => x"00",
         17454 => x"00",
         17455 => x"00",
         17456 => x"00",
         17457 => x"00",
         17458 => x"00",
         17459 => x"00",
         17460 => x"00",
         17461 => x"00",
         17462 => x"00",
         17463 => x"00",
         17464 => x"00",
         17465 => x"00",
         17466 => x"00",
         17467 => x"00",
         17468 => x"00",
         17469 => x"00",
         17470 => x"00",
         17471 => x"00",
         17472 => x"00",
         17473 => x"00",
         17474 => x"00",
         17475 => x"00",
         17476 => x"00",
         17477 => x"00",
         17478 => x"00",
         17479 => x"00",
         17480 => x"00",
         17481 => x"00",
         17482 => x"00",
         17483 => x"00",
         17484 => x"00",
         17485 => x"00",
         17486 => x"00",
         17487 => x"00",
         17488 => x"00",
         17489 => x"00",
         17490 => x"00",
         17491 => x"00",
         17492 => x"00",
         17493 => x"00",
         17494 => x"00",
         17495 => x"00",
         17496 => x"00",
         17497 => x"00",
         17498 => x"00",
         17499 => x"00",
         17500 => x"00",
         17501 => x"00",
         17502 => x"00",
         17503 => x"00",
         17504 => x"00",
         17505 => x"00",
         17506 => x"00",
         17507 => x"00",
         17508 => x"00",
         17509 => x"00",
         17510 => x"00",
         17511 => x"00",
         17512 => x"00",
         17513 => x"00",
         17514 => x"00",
         17515 => x"00",
         17516 => x"00",
         17517 => x"00",
         17518 => x"00",
         17519 => x"00",
         17520 => x"00",
         17521 => x"00",
         17522 => x"00",
         17523 => x"00",
         17524 => x"00",
         17525 => x"00",
         17526 => x"00",
         17527 => x"00",
         17528 => x"00",
         17529 => x"00",
         17530 => x"00",
         17531 => x"00",
         17532 => x"00",
         17533 => x"00",
         17534 => x"00",
         17535 => x"00",
         17536 => x"00",
         17537 => x"00",
         17538 => x"00",
         17539 => x"00",
         17540 => x"00",
         17541 => x"00",
         17542 => x"00",
         17543 => x"00",
         17544 => x"00",
         17545 => x"00",
         17546 => x"00",
         17547 => x"00",
         17548 => x"00",
         17549 => x"00",
         17550 => x"00",
         17551 => x"00",
         17552 => x"00",
         17553 => x"00",
         17554 => x"00",
         17555 => x"00",
         17556 => x"00",
         17557 => x"00",
         17558 => x"00",
         17559 => x"00",
         17560 => x"00",
         17561 => x"00",
         17562 => x"00",
         17563 => x"00",
         17564 => x"00",
         17565 => x"00",
         17566 => x"00",
         17567 => x"00",
         17568 => x"00",
         17569 => x"00",
         17570 => x"00",
         17571 => x"00",
         17572 => x"00",
         17573 => x"00",
         17574 => x"00",
         17575 => x"00",
         17576 => x"00",
         17577 => x"00",
         17578 => x"00",
         17579 => x"00",
         17580 => x"00",
         17581 => x"00",
         17582 => x"00",
         17583 => x"00",
         17584 => x"00",
         17585 => x"00",
         17586 => x"00",
         17587 => x"00",
         17588 => x"00",
         17589 => x"00",
         17590 => x"00",
         17591 => x"00",
         17592 => x"00",
         17593 => x"00",
         17594 => x"00",
         17595 => x"00",
         17596 => x"00",
         17597 => x"00",
         17598 => x"00",
         17599 => x"00",
         17600 => x"00",
         17601 => x"00",
         17602 => x"00",
         17603 => x"00",
         17604 => x"00",
         17605 => x"00",
         17606 => x"00",
         17607 => x"00",
         17608 => x"00",
         17609 => x"00",
         17610 => x"00",
         17611 => x"00",
         17612 => x"00",
         17613 => x"00",
         17614 => x"00",
         17615 => x"00",
         17616 => x"00",
         17617 => x"00",
         17618 => x"00",
         17619 => x"00",
         17620 => x"00",
         17621 => x"00",
         17622 => x"00",
         17623 => x"00",
         17624 => x"00",
         17625 => x"00",
         17626 => x"00",
         17627 => x"00",
         17628 => x"00",
         17629 => x"00",
         17630 => x"00",
         17631 => x"00",
         17632 => x"00",
         17633 => x"00",
         17634 => x"00",
         17635 => x"00",
         17636 => x"00",
         17637 => x"00",
         17638 => x"00",
         17639 => x"00",
         17640 => x"00",
         17641 => x"00",
         17642 => x"00",
         17643 => x"00",
         17644 => x"00",
         17645 => x"00",
         17646 => x"00",
         17647 => x"00",
         17648 => x"00",
         17649 => x"00",
         17650 => x"00",
         17651 => x"00",
         17652 => x"00",
         17653 => x"00",
         17654 => x"00",
         17655 => x"00",
         17656 => x"00",
         17657 => x"00",
         17658 => x"00",
         17659 => x"00",
         17660 => x"00",
         17661 => x"00",
         17662 => x"00",
         17663 => x"00",
         17664 => x"00",
         17665 => x"00",
         17666 => x"00",
         17667 => x"00",
         17668 => x"00",
         17669 => x"00",
         17670 => x"00",
         17671 => x"00",
         17672 => x"00",
         17673 => x"00",
         17674 => x"00",
         17675 => x"00",
         17676 => x"00",
         17677 => x"00",
         17678 => x"00",
         17679 => x"00",
         17680 => x"00",
         17681 => x"00",
         17682 => x"00",
         17683 => x"00",
         17684 => x"00",
         17685 => x"00",
         17686 => x"00",
         17687 => x"00",
         17688 => x"00",
         17689 => x"00",
         17690 => x"00",
         17691 => x"00",
         17692 => x"00",
         17693 => x"00",
         17694 => x"00",
         17695 => x"00",
         17696 => x"00",
         17697 => x"00",
         17698 => x"00",
         17699 => x"00",
         17700 => x"00",
         17701 => x"00",
         17702 => x"00",
         17703 => x"00",
         17704 => x"00",
         17705 => x"00",
         17706 => x"00",
         17707 => x"00",
         17708 => x"00",
         17709 => x"00",
         17710 => x"00",
         17711 => x"00",
         17712 => x"00",
         17713 => x"00",
         17714 => x"00",
         17715 => x"00",
         17716 => x"00",
         17717 => x"00",
         17718 => x"00",
         17719 => x"00",
         17720 => x"00",
         17721 => x"00",
         17722 => x"00",
         17723 => x"00",
         17724 => x"00",
         17725 => x"00",
         17726 => x"00",
         17727 => x"00",
         17728 => x"00",
         17729 => x"00",
         17730 => x"00",
         17731 => x"00",
         17732 => x"00",
         17733 => x"00",
         17734 => x"00",
         17735 => x"00",
         17736 => x"00",
         17737 => x"00",
         17738 => x"00",
         17739 => x"00",
         17740 => x"00",
         17741 => x"00",
         17742 => x"00",
         17743 => x"00",
         17744 => x"00",
         17745 => x"00",
         17746 => x"00",
         17747 => x"00",
         17748 => x"00",
         17749 => x"00",
         17750 => x"00",
         17751 => x"00",
         17752 => x"00",
         17753 => x"00",
         17754 => x"00",
         17755 => x"00",
         17756 => x"00",
         17757 => x"00",
         17758 => x"00",
         17759 => x"00",
         17760 => x"00",
         17761 => x"00",
         17762 => x"00",
         17763 => x"00",
         17764 => x"00",
         17765 => x"00",
         17766 => x"00",
         17767 => x"00",
         17768 => x"00",
         17769 => x"00",
         17770 => x"00",
         17771 => x"00",
         17772 => x"00",
         17773 => x"00",
         17774 => x"00",
         17775 => x"00",
         17776 => x"00",
         17777 => x"00",
         17778 => x"00",
         17779 => x"00",
         17780 => x"00",
         17781 => x"00",
         17782 => x"00",
         17783 => x"00",
         17784 => x"00",
         17785 => x"00",
         17786 => x"00",
         17787 => x"00",
         17788 => x"00",
         17789 => x"00",
         17790 => x"00",
         17791 => x"00",
         17792 => x"00",
         17793 => x"00",
         17794 => x"00",
         17795 => x"00",
         17796 => x"00",
         17797 => x"00",
         17798 => x"00",
         17799 => x"00",
         17800 => x"00",
         17801 => x"00",
         17802 => x"00",
         17803 => x"00",
         17804 => x"00",
         17805 => x"00",
         17806 => x"00",
         17807 => x"00",
         17808 => x"00",
         17809 => x"00",
         17810 => x"00",
         17811 => x"00",
         17812 => x"00",
         17813 => x"00",
         17814 => x"00",
         17815 => x"00",
         17816 => x"00",
         17817 => x"00",
         17818 => x"00",
         17819 => x"00",
         17820 => x"00",
         17821 => x"00",
         17822 => x"00",
         17823 => x"00",
         17824 => x"00",
         17825 => x"00",
         17826 => x"00",
         17827 => x"00",
         17828 => x"00",
         17829 => x"00",
         17830 => x"00",
         17831 => x"00",
         17832 => x"00",
         17833 => x"00",
         17834 => x"00",
         17835 => x"00",
         17836 => x"00",
         17837 => x"00",
         17838 => x"00",
         17839 => x"00",
         17840 => x"00",
         17841 => x"00",
         17842 => x"00",
         17843 => x"00",
         17844 => x"00",
         17845 => x"00",
         17846 => x"00",
         17847 => x"00",
         17848 => x"00",
         17849 => x"00",
         17850 => x"00",
         17851 => x"00",
         17852 => x"00",
         17853 => x"00",
         17854 => x"00",
         17855 => x"00",
         17856 => x"00",
         17857 => x"00",
         17858 => x"00",
         17859 => x"00",
         17860 => x"00",
         17861 => x"00",
         17862 => x"00",
         17863 => x"00",
         17864 => x"00",
         17865 => x"00",
         17866 => x"00",
         17867 => x"00",
         17868 => x"00",
         17869 => x"00",
         17870 => x"00",
         17871 => x"00",
         17872 => x"00",
         17873 => x"00",
         17874 => x"00",
         17875 => x"00",
         17876 => x"00",
         17877 => x"00",
         17878 => x"00",
         17879 => x"00",
         17880 => x"00",
         17881 => x"00",
         17882 => x"00",
         17883 => x"00",
         17884 => x"00",
         17885 => x"00",
         17886 => x"00",
         17887 => x"00",
         17888 => x"00",
         17889 => x"00",
         17890 => x"00",
         17891 => x"00",
         17892 => x"00",
         17893 => x"00",
         17894 => x"00",
         17895 => x"00",
         17896 => x"00",
         17897 => x"00",
         17898 => x"00",
         17899 => x"00",
         17900 => x"00",
         17901 => x"00",
         17902 => x"00",
         17903 => x"00",
         17904 => x"00",
         17905 => x"00",
         17906 => x"00",
         17907 => x"00",
         17908 => x"00",
         17909 => x"00",
         17910 => x"00",
         17911 => x"00",
         17912 => x"00",
         17913 => x"00",
         17914 => x"00",
         17915 => x"00",
         17916 => x"00",
         17917 => x"00",
         17918 => x"00",
         17919 => x"00",
         17920 => x"00",
         17921 => x"00",
         17922 => x"00",
         17923 => x"00",
         17924 => x"00",
         17925 => x"00",
         17926 => x"00",
         17927 => x"00",
         17928 => x"00",
         17929 => x"00",
         17930 => x"00",
         17931 => x"00",
         17932 => x"00",
         17933 => x"00",
         17934 => x"00",
         17935 => x"00",
         17936 => x"00",
         17937 => x"00",
         17938 => x"00",
         17939 => x"00",
         17940 => x"00",
         17941 => x"00",
         17942 => x"00",
         17943 => x"00",
         17944 => x"00",
         17945 => x"00",
         17946 => x"00",
         17947 => x"00",
         17948 => x"00",
         17949 => x"00",
         17950 => x"00",
         17951 => x"00",
         17952 => x"00",
         17953 => x"00",
         17954 => x"00",
         17955 => x"00",
         17956 => x"00",
         17957 => x"00",
         17958 => x"00",
         17959 => x"00",
         17960 => x"00",
         17961 => x"00",
         17962 => x"00",
         17963 => x"00",
         17964 => x"00",
         17965 => x"00",
         17966 => x"00",
         17967 => x"00",
         17968 => x"00",
         17969 => x"00",
         17970 => x"00",
         17971 => x"00",
         17972 => x"00",
         17973 => x"00",
         17974 => x"00",
         17975 => x"00",
         17976 => x"00",
         17977 => x"00",
         17978 => x"00",
         17979 => x"00",
         17980 => x"00",
         17981 => x"00",
         17982 => x"00",
         17983 => x"00",
         17984 => x"00",
         17985 => x"00",
         17986 => x"00",
         17987 => x"00",
         17988 => x"00",
         17989 => x"00",
         17990 => x"00",
         17991 => x"00",
         17992 => x"00",
         17993 => x"00",
         17994 => x"00",
         17995 => x"00",
         17996 => x"00",
         17997 => x"00",
         17998 => x"00",
         17999 => x"00",
         18000 => x"00",
         18001 => x"00",
         18002 => x"00",
         18003 => x"00",
         18004 => x"00",
         18005 => x"00",
         18006 => x"00",
         18007 => x"00",
         18008 => x"00",
         18009 => x"00",
         18010 => x"00",
         18011 => x"00",
         18012 => x"00",
         18013 => x"00",
         18014 => x"00",
         18015 => x"00",
         18016 => x"00",
         18017 => x"00",
         18018 => x"00",
         18019 => x"00",
         18020 => x"00",
         18021 => x"00",
         18022 => x"00",
         18023 => x"00",
         18024 => x"00",
         18025 => x"00",
         18026 => x"00",
         18027 => x"00",
         18028 => x"00",
         18029 => x"00",
         18030 => x"00",
         18031 => x"00",
         18032 => x"00",
         18033 => x"00",
         18034 => x"00",
         18035 => x"00",
         18036 => x"00",
         18037 => x"00",
         18038 => x"00",
         18039 => x"00",
         18040 => x"00",
         18041 => x"00",
         18042 => x"00",
         18043 => x"00",
         18044 => x"00",
         18045 => x"00",
         18046 => x"00",
         18047 => x"00",
         18048 => x"00",
         18049 => x"00",
         18050 => x"00",
         18051 => x"00",
         18052 => x"00",
         18053 => x"00",
         18054 => x"00",
         18055 => x"00",
         18056 => x"00",
         18057 => x"00",
         18058 => x"00",
         18059 => x"00",
         18060 => x"00",
         18061 => x"00",
         18062 => x"00",
         18063 => x"00",
         18064 => x"00",
         18065 => x"00",
         18066 => x"00",
         18067 => x"00",
         18068 => x"00",
         18069 => x"00",
         18070 => x"00",
         18071 => x"00",
         18072 => x"00",
         18073 => x"00",
         18074 => x"00",
         18075 => x"00",
         18076 => x"00",
         18077 => x"00",
         18078 => x"00",
         18079 => x"00",
         18080 => x"00",
         18081 => x"00",
         18082 => x"00",
         18083 => x"00",
         18084 => x"00",
         18085 => x"00",
         18086 => x"00",
         18087 => x"00",
         18088 => x"00",
         18089 => x"00",
         18090 => x"00",
         18091 => x"00",
         18092 => x"00",
         18093 => x"00",
         18094 => x"00",
         18095 => x"00",
         18096 => x"00",
         18097 => x"00",
         18098 => x"00",
         18099 => x"00",
         18100 => x"00",
         18101 => x"00",
         18102 => x"00",
         18103 => x"00",
         18104 => x"00",
         18105 => x"00",
         18106 => x"00",
         18107 => x"00",
         18108 => x"00",
         18109 => x"00",
         18110 => x"00",
         18111 => x"00",
         18112 => x"00",
         18113 => x"00",
         18114 => x"00",
         18115 => x"00",
         18116 => x"00",
         18117 => x"00",
         18118 => x"00",
         18119 => x"00",
         18120 => x"00",
         18121 => x"00",
         18122 => x"00",
         18123 => x"00",
         18124 => x"00",
         18125 => x"00",
         18126 => x"00",
         18127 => x"00",
         18128 => x"00",
         18129 => x"00",
         18130 => x"00",
         18131 => x"00",
         18132 => x"00",
         18133 => x"00",
         18134 => x"00",
         18135 => x"00",
         18136 => x"00",
         18137 => x"00",
         18138 => x"00",
         18139 => x"00",
         18140 => x"00",
         18141 => x"00",
         18142 => x"00",
         18143 => x"00",
         18144 => x"00",
         18145 => x"00",
         18146 => x"00",
         18147 => x"00",
         18148 => x"00",
         18149 => x"00",
         18150 => x"00",
         18151 => x"00",
         18152 => x"00",
         18153 => x"00",
         18154 => x"00",
         18155 => x"00",
         18156 => x"00",
         18157 => x"00",
         18158 => x"00",
         18159 => x"00",
         18160 => x"00",
         18161 => x"00",
         18162 => x"00",
         18163 => x"00",
         18164 => x"00",
         18165 => x"00",
         18166 => x"00",
         18167 => x"00",
         18168 => x"00",
         18169 => x"00",
         18170 => x"00",
         18171 => x"00",
         18172 => x"00",
         18173 => x"00",
         18174 => x"00",
         18175 => x"00",
         18176 => x"00",
         18177 => x"00",
         18178 => x"00",
         18179 => x"00",
         18180 => x"00",
         18181 => x"00",
         18182 => x"00",
         18183 => x"00",
         18184 => x"00",
         18185 => x"00",
         18186 => x"00",
         18187 => x"00",
         18188 => x"00",
         18189 => x"00",
         18190 => x"00",
         18191 => x"00",
         18192 => x"00",
         18193 => x"00",
         18194 => x"00",
         18195 => x"00",
         18196 => x"00",
         18197 => x"00",
         18198 => x"00",
         18199 => x"00",
         18200 => x"00",
         18201 => x"00",
         18202 => x"00",
         18203 => x"00",
         18204 => x"00",
         18205 => x"00",
         18206 => x"50",
         18207 => x"00",
         18208 => x"cc",
         18209 => x"ce",
         18210 => x"f8",
         18211 => x"fc",
         18212 => x"e1",
         18213 => x"c4",
         18214 => x"e3",
         18215 => x"eb",
         18216 => x"00",
         18217 => x"64",
         18218 => x"68",
         18219 => x"2f",
         18220 => x"20",
         18221 => x"24",
         18222 => x"28",
         18223 => x"51",
         18224 => x"55",
         18225 => x"04",
         18226 => x"08",
         18227 => x"0c",
         18228 => x"10",
         18229 => x"14",
         18230 => x"18",
         18231 => x"59",
         18232 => x"c7",
         18233 => x"84",
         18234 => x"88",
         18235 => x"8c",
         18236 => x"90",
         18237 => x"94",
         18238 => x"98",
         18239 => x"80",
         18240 => x"00",
         18241 => x"00",
         18242 => x"00",
         18243 => x"00",
         18244 => x"00",
         18245 => x"00",
         18246 => x"00",
         18247 => x"00",
         18248 => x"00",
         18249 => x"00",
         18250 => x"00",
         18251 => x"00",
         18252 => x"00",
         18253 => x"00",
         18254 => x"00",
         18255 => x"00",
         18256 => x"00",
         18257 => x"00",
         18258 => x"00",
         18259 => x"00",
         18260 => x"00",
         18261 => x"00",
         18262 => x"00",
         18263 => x"00",
         18264 => x"00",
         18265 => x"00",
         18266 => x"00",
         18267 => x"00",
         18268 => x"00",
         18269 => x"00",
         18270 => x"00",
         18271 => x"00",
         18272 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
