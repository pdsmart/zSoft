-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87fa",
             1 => x"f80d0b0b",
             2 => x"0b93e904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"cd040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b93b0",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b83bd",
           162 => x"e4738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93b50400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0bac",
           171 => x"cc2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0bab",
           179 => x"ab2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"96040b0b",
           269 => x"0b8ca604",
           270 => x"0b0b0b8c",
           271 => x"b6040b0b",
           272 => x"0b8cc604",
           273 => x"0b0b0b8c",
           274 => x"d6040b0b",
           275 => x"0b8ce604",
           276 => x"0b0b0b8c",
           277 => x"f6040b0b",
           278 => x"0b8d8604",
           279 => x"0b0b0b8d",
           280 => x"96040b0b",
           281 => x"0b8da604",
           282 => x"0b0b0b8d",
           283 => x"b6040b0b",
           284 => x"0b8dc604",
           285 => x"0b0b0b8d",
           286 => x"d7040b0b",
           287 => x"0b8de804",
           288 => x"0b0b0b8d",
           289 => x"f9040b0b",
           290 => x"0b8e8a04",
           291 => x"0b0b0b8e",
           292 => x"9b040b0b",
           293 => x"0b8eac04",
           294 => x"0b0b0b8e",
           295 => x"bd040b0b",
           296 => x"0b8ece04",
           297 => x"0b0b0b8e",
           298 => x"df040b0b",
           299 => x"0b8ef004",
           300 => x"0b0b0b8f",
           301 => x"81040b0b",
           302 => x"0b8f9204",
           303 => x"0b0b0b8f",
           304 => x"a3040b0b",
           305 => x"0b8fb404",
           306 => x"0b0b0b8f",
           307 => x"c5040b0b",
           308 => x"0b8fd604",
           309 => x"0b0b0b8f",
           310 => x"e7040b0b",
           311 => x"0b8ff804",
           312 => x"0b0b0b90",
           313 => x"89040b0b",
           314 => x"0b909a04",
           315 => x"0b0b0b90",
           316 => x"ab040b0b",
           317 => x"0b90bc04",
           318 => x"0b0b0b90",
           319 => x"cd040b0b",
           320 => x"0b90de04",
           321 => x"0b0b0b90",
           322 => x"ef040b0b",
           323 => x"0b918004",
           324 => x"0b0b0b91",
           325 => x"91040b0b",
           326 => x"0b91a204",
           327 => x"0b0b0b91",
           328 => x"b3040b0b",
           329 => x"0b91c404",
           330 => x"0b0b0b91",
           331 => x"d5040b0b",
           332 => x"0b91e604",
           333 => x"0b0b0b91",
           334 => x"f7040b0b",
           335 => x"0b928804",
           336 => x"0b0b0b92",
           337 => x"99040b0b",
           338 => x"0b92aa04",
           339 => x"0b0b0b92",
           340 => x"bb040b0b",
           341 => x"0b92cb04",
           342 => x"0b0b0b92",
           343 => x"dc040b0b",
           344 => x"0b92ed04",
           345 => x"0b0b0b92",
           346 => x"fe04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0484b8f0",
           386 => x"0c80d5ec",
           387 => x"2d84b8f0",
           388 => x"0880c080",
           389 => x"900484b8",
           390 => x"f00ca2ee",
           391 => x"2d84b8f0",
           392 => x"0880c080",
           393 => x"900484b8",
           394 => x"f00ca0f3",
           395 => x"2d84b8f0",
           396 => x"0880c080",
           397 => x"900484b8",
           398 => x"f00ca0e0",
           399 => x"2d84b8f0",
           400 => x"0880c080",
           401 => x"900484b8",
           402 => x"f00c94a3",
           403 => x"2d84b8f0",
           404 => x"0880c080",
           405 => x"900484b8",
           406 => x"f00ca1f6",
           407 => x"2d84b8f0",
           408 => x"0880c080",
           409 => x"900484b8",
           410 => x"f00caf86",
           411 => x"2d84b8f0",
           412 => x"0880c080",
           413 => x"900484b8",
           414 => x"f00cad82",
           415 => x"2d84b8f0",
           416 => x"0880c080",
           417 => x"900484b8",
           418 => x"f00c9488",
           419 => x"2d84b8f0",
           420 => x"0880c080",
           421 => x"900484b8",
           422 => x"f00c95a8",
           423 => x"2d84b8f0",
           424 => x"0880c080",
           425 => x"900484b8",
           426 => x"f00c95d1",
           427 => x"2d84b8f0",
           428 => x"0880c080",
           429 => x"900484b8",
           430 => x"f00cb18a",
           431 => x"2d84b8f0",
           432 => x"0880c080",
           433 => x"900484b8",
           434 => x"f00c80d4",
           435 => x"d12d84b8",
           436 => x"f00880c0",
           437 => x"80900484",
           438 => x"b8f00c80",
           439 => x"d5b62d84",
           440 => x"b8f00880",
           441 => x"c0809004",
           442 => x"84b8f00c",
           443 => x"80d28d2d",
           444 => x"84b8f008",
           445 => x"80c08090",
           446 => x"0484b8f0",
           447 => x"0c80d3c0",
           448 => x"2d84b8f0",
           449 => x"0880c080",
           450 => x"900484b8",
           451 => x"f00c82c9",
           452 => x"9d2d84b8",
           453 => x"f00880c0",
           454 => x"80900484",
           455 => x"b8f00c82",
           456 => x"e2ef2d84",
           457 => x"b8f00880",
           458 => x"c0809004",
           459 => x"84b8f00c",
           460 => x"82d28d2d",
           461 => x"84b8f008",
           462 => x"80c08090",
           463 => x"0484b8f0",
           464 => x"0c82d7af",
           465 => x"2d84b8f0",
           466 => x"0880c080",
           467 => x"900484b8",
           468 => x"f00c82ed",
           469 => x"8c2d84b8",
           470 => x"f00880c0",
           471 => x"80900484",
           472 => x"b8f00c82",
           473 => x"fa942d84",
           474 => x"b8f00880",
           475 => x"c0809004",
           476 => x"84b8f00c",
           477 => x"82def62d",
           478 => x"84b8f008",
           479 => x"80c08090",
           480 => x"0484b8f0",
           481 => x"0c82f1ad",
           482 => x"2d84b8f0",
           483 => x"0880c080",
           484 => x"900484b8",
           485 => x"f00c82f2",
           486 => x"fa2d84b8",
           487 => x"f00880c0",
           488 => x"80900484",
           489 => x"b8f00c82",
           490 => x"f3cf2d84",
           491 => x"b8f00880",
           492 => x"c0809004",
           493 => x"84b8f00c",
           494 => x"8384912d",
           495 => x"84b8f008",
           496 => x"80c08090",
           497 => x"0484b8f0",
           498 => x"0c82fed6",
           499 => x"2d84b8f0",
           500 => x"0880c080",
           501 => x"900484b8",
           502 => x"f00c838a",
           503 => x"f52d84b8",
           504 => x"f00880c0",
           505 => x"80900484",
           506 => x"b8f00c82",
           507 => x"f5ac2d84",
           508 => x"b8f00880",
           509 => x"c0809004",
           510 => x"84b8f00c",
           511 => x"8393ec2d",
           512 => x"84b8f008",
           513 => x"80c08090",
           514 => x"0484b8f0",
           515 => x"0c8394f7",
           516 => x"2d84b8f0",
           517 => x"0880c080",
           518 => x"900484b8",
           519 => x"f00c82e5",
           520 => x"bf2d84b8",
           521 => x"f00880c0",
           522 => x"80900484",
           523 => x"b8f00c82",
           524 => x"e3d62d84",
           525 => x"b8f00880",
           526 => x"c0809004",
           527 => x"84b8f00c",
           528 => x"82e6fd2d",
           529 => x"84b8f008",
           530 => x"80c08090",
           531 => x"0484b8f0",
           532 => x"0c82f696",
           533 => x"2d84b8f0",
           534 => x"0880c080",
           535 => x"900484b8",
           536 => x"f00c8396",
           537 => x"892d84b8",
           538 => x"f00880c0",
           539 => x"80900484",
           540 => x"b8f00c83",
           541 => x"99e62d84",
           542 => x"b8f00880",
           543 => x"c0809004",
           544 => x"84b8f00c",
           545 => x"83a0d82d",
           546 => x"84b8f008",
           547 => x"80c08090",
           548 => x"0484b8f0",
           549 => x"0c82c6ee",
           550 => x"2d84b8f0",
           551 => x"0880c080",
           552 => x"900484b8",
           553 => x"f00c83a4",
           554 => x"812d84b8",
           555 => x"f00880c0",
           556 => x"80900484",
           557 => x"b8f00c83",
           558 => x"b9822d84",
           559 => x"b8f00880",
           560 => x"c0809004",
           561 => x"84b8f00c",
           562 => x"83b7b42d",
           563 => x"84b8f008",
           564 => x"80c08090",
           565 => x"0484b8f0",
           566 => x"0c81f3d2",
           567 => x"2d84b8f0",
           568 => x"0880c080",
           569 => x"900484b8",
           570 => x"f00c81f4",
           571 => x"d12d84b8",
           572 => x"f00880c0",
           573 => x"80900484",
           574 => x"b8f00c81",
           575 => x"f5d02d84",
           576 => x"b8f00880",
           577 => x"c0809004",
           578 => x"84b8f00c",
           579 => x"80d08f2d",
           580 => x"84b8f008",
           581 => x"80c08090",
           582 => x"0484b8f0",
           583 => x"0c80d1df",
           584 => x"2d84b8f0",
           585 => x"0880c080",
           586 => x"900484b8",
           587 => x"f00c80d7",
           588 => x"8a2d84b8",
           589 => x"f00880c0",
           590 => x"80900484",
           591 => x"b8f00cb1",
           592 => x"9a2d84b8",
           593 => x"f00880c0",
           594 => x"80900484",
           595 => x"b8f00c81",
           596 => x"daf02d84",
           597 => x"b8f00880",
           598 => x"c0809004",
           599 => x"84b8f00c",
           600 => x"81dcab2d",
           601 => x"84b8f008",
           602 => x"80c08090",
           603 => x"0484b8f0",
           604 => x"0c81f1ac",
           605 => x"2d84b8f0",
           606 => x"0880c080",
           607 => x"900484b8",
           608 => x"f00c81d5",
           609 => x"802d84b8",
           610 => x"f00880c0",
           611 => x"8090043c",
           612 => x"04101010",
           613 => x"10101010",
           614 => x"10101010",
           615 => x"10101010",
           616 => x"10101010",
           617 => x"10101010",
           618 => x"10101010",
           619 => x"10101010",
           620 => x"53510400",
           621 => x"007381ff",
           622 => x"06738306",
           623 => x"09810583",
           624 => x"05101010",
           625 => x"2b0772fc",
           626 => x"060c5151",
           627 => x"04727280",
           628 => x"728106ff",
           629 => x"05097206",
           630 => x"05711052",
           631 => x"720a100a",
           632 => x"5372ed38",
           633 => x"51515351",
           634 => x"0484b8e4",
           635 => x"7084d4d0",
           636 => x"278e3880",
           637 => x"71708405",
           638 => x"530c0b0b",
           639 => x"0b93ec04",
           640 => x"8c815180",
           641 => x"ceba0400",
           642 => x"fc3d0d87",
           643 => x"3d707084",
           644 => x"05520856",
           645 => x"53745284",
           646 => x"d4c80851",
           647 => x"81c53f86",
           648 => x"3d0d04fa",
           649 => x"3d0d787a",
           650 => x"7c851133",
           651 => x"81328106",
           652 => x"80732507",
           653 => x"56585557",
           654 => x"80527272",
           655 => x"2e098106",
           656 => x"80d338ff",
           657 => x"1477748a",
           658 => x"32703070",
           659 => x"72079f2a",
           660 => x"51555556",
           661 => x"54807425",
           662 => x"b7387180",
           663 => x"2eb23875",
           664 => x"518efa3f",
           665 => x"84b8e408",
           666 => x"5384b8e4",
           667 => x"08ff2eae",
           668 => x"3884b8e4",
           669 => x"08757081",
           670 => x"055734ff",
           671 => x"14738a32",
           672 => x"70307072",
           673 => x"079f2a51",
           674 => x"54545473",
           675 => x"8024cb38",
           676 => x"80753476",
           677 => x"527184b8",
           678 => x"e40c883d",
           679 => x"0d04800b",
           680 => x"84b8e40c",
           681 => x"883d0d04",
           682 => x"f53d0d7d",
           683 => x"54860284",
           684 => x"05990534",
           685 => x"7356fe0a",
           686 => x"588e3d88",
           687 => x"05537e52",
           688 => x"8d3de405",
           689 => x"519d3f73",
           690 => x"19548074",
           691 => x"348d3d0d",
           692 => x"04fd3d0d",
           693 => x"863d8805",
           694 => x"53765275",
           695 => x"51853f85",
           696 => x"3d0d04f1",
           697 => x"3d0d6163",
           698 => x"65425d5d",
           699 => x"80708c1f",
           700 => x"0c851e33",
           701 => x"70812a81",
           702 => x"32810655",
           703 => x"555bff54",
           704 => x"727b2e09",
           705 => x"810680d2",
           706 => x"387b3357",
           707 => x"767b2e80",
           708 => x"c538811c",
           709 => x"7b810654",
           710 => x"5c72802e",
           711 => x"818138d0",
           712 => x"175f7e89",
           713 => x"2681a338",
           714 => x"76b03270",
           715 => x"30708025",
           716 => x"51545578",
           717 => x"ae387280",
           718 => x"2ea9387a",
           719 => x"832a7081",
           720 => x"32810640",
           721 => x"547e802e",
           722 => x"9e387a82",
           723 => x"80075b7b",
           724 => x"335776ff",
           725 => x"bd388c1d",
           726 => x"08547384",
           727 => x"b8e40c91",
           728 => x"3d0d047a",
           729 => x"832a5478",
           730 => x"10101079",
           731 => x"10057098",
           732 => x"2b70982c",
           733 => x"19708180",
           734 => x"0a298b0a",
           735 => x"0570982c",
           736 => x"525a5b56",
           737 => x"5f807924",
           738 => x"81863873",
           739 => x"81065372",
           740 => x"ffbd3878",
           741 => x"7c335858",
           742 => x"76fef738",
           743 => x"ffb83976",
           744 => x"a52e0981",
           745 => x"06933881",
           746 => x"73745a5a",
           747 => x"5b8a7c33",
           748 => x"585a76fe",
           749 => x"dd38ff9e",
           750 => x"397c5276",
           751 => x"518baf3f",
           752 => x"7b335776",
           753 => x"fecc38ff",
           754 => x"8d397a83",
           755 => x"2a708106",
           756 => x"5455788a",
           757 => x"38817074",
           758 => x"0640547e",
           759 => x"9538e017",
           760 => x"537280d8",
           761 => x"26973872",
           762 => x"101083c9",
           763 => x"f4055473",
           764 => x"080473e0",
           765 => x"18545980",
           766 => x"d87327eb",
           767 => x"387c5276",
           768 => x"518aeb3f",
           769 => x"807c3358",
           770 => x"5b76fe86",
           771 => x"38fec739",
           772 => x"80ff59fe",
           773 => x"f639885a",
           774 => x"7f608405",
           775 => x"71087d83",
           776 => x"ffcf065e",
           777 => x"58415484",
           778 => x"b8f45e79",
           779 => x"52755193",
           780 => x"9a3f84b8",
           781 => x"e40881ff",
           782 => x"0684b8e4",
           783 => x"0818df05",
           784 => x"56537289",
           785 => x"26883884",
           786 => x"b8e408b0",
           787 => x"0555747e",
           788 => x"70810540",
           789 => x"34795275",
           790 => x"5190ca3f",
           791 => x"84b8e408",
           792 => x"5684b8e4",
           793 => x"08c5387d",
           794 => x"84b8f431",
           795 => x"982b7bb2",
           796 => x"0640567e",
           797 => x"802e8f38",
           798 => x"77848080",
           799 => x"29fc8080",
           800 => x"0570902c",
           801 => x"59557a86",
           802 => x"2a708106",
           803 => x"555f7380",
           804 => x"2e9e3877",
           805 => x"84808029",
           806 => x"f8808005",
           807 => x"5379902e",
           808 => x"8b387784",
           809 => x"808029fc",
           810 => x"80800553",
           811 => x"72902c58",
           812 => x"7a832a70",
           813 => x"81065455",
           814 => x"72802e9e",
           815 => x"3875982c",
           816 => x"7081ff06",
           817 => x"54547873",
           818 => x"2486cc38",
           819 => x"7a83fff7",
           820 => x"0670832a",
           821 => x"71862a41",
           822 => x"565b7481",
           823 => x"06547380",
           824 => x"2e85f038",
           825 => x"77793190",
           826 => x"2b70902c",
           827 => x"7c838006",
           828 => x"56595373",
           829 => x"802e8596",
           830 => x"387a812a",
           831 => x"81065473",
           832 => x"85eb387a",
           833 => x"842a8106",
           834 => x"54738698",
           835 => x"387a852a",
           836 => x"81065473",
           837 => x"8697387e",
           838 => x"81065473",
           839 => x"858f387a",
           840 => x"882a8106",
           841 => x"5f7e802e",
           842 => x"b2387778",
           843 => x"84808029",
           844 => x"fc808005",
           845 => x"70902c5a",
           846 => x"40548074",
           847 => x"259d387c",
           848 => x"52b05188",
           849 => x"a93f7778",
           850 => x"84808029",
           851 => x"fc808005",
           852 => x"70902c5a",
           853 => x"40547380",
           854 => x"24e53874",
           855 => x"81065372",
           856 => x"802eb238",
           857 => x"78798180",
           858 => x"0a2981ff",
           859 => x"0a057098",
           860 => x"2c5b5555",
           861 => x"8075259d",
           862 => x"387c52b0",
           863 => x"5187ef3f",
           864 => x"78798180",
           865 => x"0a2981ff",
           866 => x"0a057098",
           867 => x"2c5b5555",
           868 => x"748024e5",
           869 => x"387a872a",
           870 => x"7081065c",
           871 => x"557a802e",
           872 => x"81b93876",
           873 => x"80e32e84",
           874 => x"d8387680",
           875 => x"f32e81ca",
           876 => x"387680d3",
           877 => x"2e81e238",
           878 => x"7d84b8f4",
           879 => x"2e96387c",
           880 => x"52ff1e70",
           881 => x"33525e87",
           882 => x"a53f7d84",
           883 => x"b8f42e09",
           884 => x"8106ec38",
           885 => x"7481065b",
           886 => x"7a802efc",
           887 => x"a7387778",
           888 => x"84808029",
           889 => x"fc808005",
           890 => x"70902c5a",
           891 => x"40558075",
           892 => x"25fc9138",
           893 => x"7c52a051",
           894 => x"86f43fe2",
           895 => x"397a9007",
           896 => x"5b7aa007",
           897 => x"7c33585b",
           898 => x"76fa8738",
           899 => x"fac8397a",
           900 => x"80c0075b",
           901 => x"80f85790",
           902 => x"60618405",
           903 => x"71087e83",
           904 => x"ffcf065f",
           905 => x"5942555a",
           906 => x"fbfd397f",
           907 => x"60840577",
           908 => x"fe800a06",
           909 => x"83133370",
           910 => x"982b7207",
           911 => x"7c848080",
           912 => x"29fc8080",
           913 => x"0570902c",
           914 => x"5e525a56",
           915 => x"57415f7a",
           916 => x"872a7081",
           917 => x"065c557a",
           918 => x"fec93877",
           919 => x"78848080",
           920 => x"29fc8080",
           921 => x"0570902c",
           922 => x"5a545f80",
           923 => x"7f25feb3",
           924 => x"387c52a0",
           925 => x"5185f73f",
           926 => x"e239ff1a",
           927 => x"7083ffff",
           928 => x"065b5779",
           929 => x"83ffff2e",
           930 => x"feca387c",
           931 => x"52757081",
           932 => x"05573351",
           933 => x"85d83fe2",
           934 => x"39ff1a70",
           935 => x"83ffff06",
           936 => x"5b547983",
           937 => x"ffff2efe",
           938 => x"ab387c52",
           939 => x"75708105",
           940 => x"57335185",
           941 => x"b93fe239",
           942 => x"75fc0a06",
           943 => x"81fc0a07",
           944 => x"78848080",
           945 => x"29fc8080",
           946 => x"0570902c",
           947 => x"5a585680",
           948 => x"e37b872a",
           949 => x"7081065d",
           950 => x"56577afd",
           951 => x"c638fefb",
           952 => x"397f6084",
           953 => x"05710870",
           954 => x"53404156",
           955 => x"807e2482",
           956 => x"df387a83",
           957 => x"ffbf065b",
           958 => x"84b8f45e",
           959 => x"faad397a",
           960 => x"84077c33",
           961 => x"585b76f8",
           962 => x"8938f8ca",
           963 => x"397a8807",
           964 => x"5b807c33",
           965 => x"585976f7",
           966 => x"f938f8ba",
           967 => x"397f6084",
           968 => x"05710877",
           969 => x"81065658",
           970 => x"415f7282",
           971 => x"8a387551",
           972 => x"87f63f84",
           973 => x"b8e40883",
           974 => x"ffff0678",
           975 => x"7131902b",
           976 => x"545a7290",
           977 => x"2c58fe87",
           978 => x"397a80c0",
           979 => x"077c3358",
           980 => x"5b76f7be",
           981 => x"38f7ff39",
           982 => x"7f608405",
           983 => x"71087781",
           984 => x"065d5841",
           985 => x"547981cf",
           986 => x"38755187",
           987 => x"bb3f84b8",
           988 => x"e40883ff",
           989 => x"ff067871",
           990 => x"31902b54",
           991 => x"5ac4397a",
           992 => x"8180077c",
           993 => x"33585b76",
           994 => x"f78838f7",
           995 => x"c9397778",
           996 => x"84808029",
           997 => x"fc808005",
           998 => x"70902c5a",
           999 => x"54548074",
          1000 => x"25fad638",
          1001 => x"7c52a051",
          1002 => x"83c43fe2",
          1003 => x"397c52b0",
          1004 => x"5183bb3f",
          1005 => x"79902e09",
          1006 => x"8106fae3",
          1007 => x"387c5276",
          1008 => x"5183ab3f",
          1009 => x"7a882a81",
          1010 => x"065f7e80",
          1011 => x"2efb8c38",
          1012 => x"fad83975",
          1013 => x"982c7871",
          1014 => x"31902b70",
          1015 => x"902c7d83",
          1016 => x"8006575a",
          1017 => x"515373fa",
          1018 => x"9038ffa2",
          1019 => x"397c52ad",
          1020 => x"5182fb3f",
          1021 => x"7e810654",
          1022 => x"73802efa",
          1023 => x"a238ffad",
          1024 => x"397c5275",
          1025 => x"982a5182",
          1026 => x"e53f7481",
          1027 => x"065b7a80",
          1028 => x"2ef7f138",
          1029 => x"fbc83978",
          1030 => x"7431982b",
          1031 => x"70982c5a",
          1032 => x"53f9b739",
          1033 => x"7c52ab51",
          1034 => x"82c43fc8",
          1035 => x"397c52a0",
          1036 => x"5182bb3f",
          1037 => x"ffbe3978",
          1038 => x"52755188",
          1039 => x"8b3f84b8",
          1040 => x"e40883ff",
          1041 => x"ff067871",
          1042 => x"31902b54",
          1043 => x"5afdf339",
          1044 => x"7a82077e",
          1045 => x"307183ff",
          1046 => x"bf065257",
          1047 => x"5bfd9939",
          1048 => x"fe3d0d84",
          1049 => x"d4c40853",
          1050 => x"75527451",
          1051 => x"f3b53f84",
          1052 => x"3d0d04fa",
          1053 => x"3d0d7855",
          1054 => x"800b84d4",
          1055 => x"c8088511",
          1056 => x"3370812a",
          1057 => x"81327081",
          1058 => x"06515658",
          1059 => x"5557ff56",
          1060 => x"72772e09",
          1061 => x"810680d5",
          1062 => x"38747081",
          1063 => x"05563353",
          1064 => x"72772eb0",
          1065 => x"3884d4c8",
          1066 => x"08527251",
          1067 => x"90140853",
          1068 => x"722d84b8",
          1069 => x"e408802e",
          1070 => x"8338ff57",
          1071 => x"74708105",
          1072 => x"56335372",
          1073 => x"802e8838",
          1074 => x"84d4c808",
          1075 => x"54d73984",
          1076 => x"d4c80854",
          1077 => x"84d4c808",
          1078 => x"528a5190",
          1079 => x"14085574",
          1080 => x"2d84b8e4",
          1081 => x"08802e83",
          1082 => x"38ff5776",
          1083 => x"567584b8",
          1084 => x"e40c883d",
          1085 => x"0d04fa3d",
          1086 => x"0d787a56",
          1087 => x"54800b85",
          1088 => x"16337081",
          1089 => x"2a813270",
          1090 => x"81065155",
          1091 => x"5757ff56",
          1092 => x"72772e09",
          1093 => x"81069238",
          1094 => x"73708105",
          1095 => x"55335372",
          1096 => x"772e0981",
          1097 => x"06983876",
          1098 => x"567584b8",
          1099 => x"e40c883d",
          1100 => x"0d047370",
          1101 => x"81055533",
          1102 => x"5372802e",
          1103 => x"ea387452",
          1104 => x"72519015",
          1105 => x"0853722d",
          1106 => x"84b8e408",
          1107 => x"802ee338",
          1108 => x"ff747081",
          1109 => x"05563354",
          1110 => x"5772e338",
          1111 => x"ca39ff3d",
          1112 => x"0d84d4c8",
          1113 => x"08527351",
          1114 => x"853f833d",
          1115 => x"0d04fa3d",
          1116 => x"0d787a85",
          1117 => x"11337081",
          1118 => x"2a813281",
          1119 => x"06565656",
          1120 => x"57ff5672",
          1121 => x"ae387382",
          1122 => x"2a810654",
          1123 => x"73802eac",
          1124 => x"388c1508",
          1125 => x"53728816",
          1126 => x"08259138",
          1127 => x"74085676",
          1128 => x"76347408",
          1129 => x"8105750c",
          1130 => x"8c150853",
          1131 => x"81138c16",
          1132 => x"0c765675",
          1133 => x"84b8e40c",
          1134 => x"883d0d04",
          1135 => x"74527681",
          1136 => x"ff065190",
          1137 => x"15085473",
          1138 => x"2dff5684",
          1139 => x"b8e408e3",
          1140 => x"388c1508",
          1141 => x"81058c16",
          1142 => x"0c7656d7",
          1143 => x"39fb3d0d",
          1144 => x"77851133",
          1145 => x"7081ff06",
          1146 => x"70813281",
          1147 => x"06555556",
          1148 => x"56ff5471",
          1149 => x"b3387286",
          1150 => x"2a810652",
          1151 => x"71b33872",
          1152 => x"822a8106",
          1153 => x"5271802e",
          1154 => x"80c33875",
          1155 => x"08703353",
          1156 => x"5371802e",
          1157 => x"80f03881",
          1158 => x"13760c8c",
          1159 => x"16088105",
          1160 => x"8c170c71",
          1161 => x"81ff0654",
          1162 => x"7384b8e4",
          1163 => x"0c873d0d",
          1164 => x"0474ffbf",
          1165 => x"06537285",
          1166 => x"17348c16",
          1167 => x"0881058c",
          1168 => x"170c8416",
          1169 => x"3384b8e4",
          1170 => x"0c873d0d",
          1171 => x"04755194",
          1172 => x"16085574",
          1173 => x"2d84b8e4",
          1174 => x"085284b8",
          1175 => x"e4088025",
          1176 => x"ffb93885",
          1177 => x"16337090",
          1178 => x"07545284",
          1179 => x"b8e408ff",
          1180 => x"2e853871",
          1181 => x"a0075372",
          1182 => x"851734ff",
          1183 => x"547384b8",
          1184 => x"e40c873d",
          1185 => x"0d0474a0",
          1186 => x"07537285",
          1187 => x"1734ff54",
          1188 => x"ec39fd3d",
          1189 => x"0d757771",
          1190 => x"54545471",
          1191 => x"70810553",
          1192 => x"335170f7",
          1193 => x"38ff1252",
          1194 => x"72708105",
          1195 => x"54335170",
          1196 => x"72708105",
          1197 => x"543470f0",
          1198 => x"387384b8",
          1199 => x"e40c853d",
          1200 => x"0d04fc3d",
          1201 => x"0d767971",
          1202 => x"7a555552",
          1203 => x"5470802e",
          1204 => x"9d387372",
          1205 => x"27a13870",
          1206 => x"802e9338",
          1207 => x"71708105",
          1208 => x"53337370",
          1209 => x"81055534",
          1210 => x"ff115170",
          1211 => x"ef387384",
          1212 => x"b8e40c86",
          1213 => x"3d0d0470",
          1214 => x"12557375",
          1215 => x"27d93870",
          1216 => x"14755353",
          1217 => x"ff13ff13",
          1218 => x"53537133",
          1219 => x"7334ff11",
          1220 => x"5170802e",
          1221 => x"d938ff13",
          1222 => x"ff135353",
          1223 => x"71337334",
          1224 => x"ff115170",
          1225 => x"df38c739",
          1226 => x"fe3d0d74",
          1227 => x"70535371",
          1228 => x"70810553",
          1229 => x"335170f7",
          1230 => x"38ff1270",
          1231 => x"743184b8",
          1232 => x"e40c5184",
          1233 => x"3d0d04fd",
          1234 => x"3d0d7577",
          1235 => x"71545454",
          1236 => x"72708105",
          1237 => x"54335170",
          1238 => x"72708105",
          1239 => x"543470f0",
          1240 => x"387384b8",
          1241 => x"e40c853d",
          1242 => x"0d04fd3d",
          1243 => x"0d757871",
          1244 => x"79555552",
          1245 => x"5470802e",
          1246 => x"93387170",
          1247 => x"81055333",
          1248 => x"73708105",
          1249 => x"5534ff11",
          1250 => x"5170ef38",
          1251 => x"7384b8e4",
          1252 => x"0c853d0d",
          1253 => x"04fc3d0d",
          1254 => x"76787a55",
          1255 => x"56547280",
          1256 => x"2ea13873",
          1257 => x"33757081",
          1258 => x"05573352",
          1259 => x"5271712e",
          1260 => x"0981069a",
          1261 => x"38811454",
          1262 => x"71802eb7",
          1263 => x"38ff1353",
          1264 => x"72e13880",
          1265 => x"517084b8",
          1266 => x"e40c863d",
          1267 => x"0d047280",
          1268 => x"2ef13873",
          1269 => x"3353ff51",
          1270 => x"72802ee9",
          1271 => x"38ff1533",
          1272 => x"52815171",
          1273 => x"802ede38",
          1274 => x"72723184",
          1275 => x"b8e40c86",
          1276 => x"3d0d0471",
          1277 => x"84b8e40c",
          1278 => x"863d0d04",
          1279 => x"fb3d0d77",
          1280 => x"79537052",
          1281 => x"5680c13f",
          1282 => x"84b8e408",
          1283 => x"84b8e408",
          1284 => x"81055255",
          1285 => x"81b2d93f",
          1286 => x"84b8e408",
          1287 => x"5484b8e4",
          1288 => x"08802e9b",
          1289 => x"3884b8e4",
          1290 => x"08155480",
          1291 => x"74347453",
          1292 => x"755284b8",
          1293 => x"e40851fe",
          1294 => x"b13f84b8",
          1295 => x"e4085473",
          1296 => x"84b8e40c",
          1297 => x"873d0d04",
          1298 => x"fd3d0d75",
          1299 => x"77717154",
          1300 => x"55535471",
          1301 => x"802e9f38",
          1302 => x"72708105",
          1303 => x"54335170",
          1304 => x"802e8c38",
          1305 => x"ff125271",
          1306 => x"ff2e0981",
          1307 => x"06ea38ff",
          1308 => x"13707531",
          1309 => x"52527084",
          1310 => x"b8e40c85",
          1311 => x"3d0d04fd",
          1312 => x"3d0d7577",
          1313 => x"79725553",
          1314 => x"54547080",
          1315 => x"2e8e3872",
          1316 => x"72708105",
          1317 => x"5434ff11",
          1318 => x"5170f438",
          1319 => x"7384b8e4",
          1320 => x"0c853d0d",
          1321 => x"04fa3d0d",
          1322 => x"787a5854",
          1323 => x"a0527680",
          1324 => x"2e8b3876",
          1325 => x"5180f53f",
          1326 => x"84b8e408",
          1327 => x"52e01253",
          1328 => x"73802e8d",
          1329 => x"38735180",
          1330 => x"e33f7184",
          1331 => x"b8e40831",
          1332 => x"53805272",
          1333 => x"9f2680cb",
          1334 => x"38735272",
          1335 => x"9f2e80c3",
          1336 => x"38811374",
          1337 => x"712aa072",
          1338 => x"3176712b",
          1339 => x"57545455",
          1340 => x"80567476",
          1341 => x"2ea83872",
          1342 => x"10749f2a",
          1343 => x"07741077",
          1344 => x"07787231",
          1345 => x"ff119f2c",
          1346 => x"7081067b",
          1347 => x"72067571",
          1348 => x"31ff1c5c",
          1349 => x"56525255",
          1350 => x"58555374",
          1351 => x"da387310",
          1352 => x"76075271",
          1353 => x"84b8e40c",
          1354 => x"883d0d04",
          1355 => x"fc3d0d76",
          1356 => x"70fc8080",
          1357 => x"06703070",
          1358 => x"72078025",
          1359 => x"70842b90",
          1360 => x"71317571",
          1361 => x"2a7083fe",
          1362 => x"80067030",
          1363 => x"70802583",
          1364 => x"2b887131",
          1365 => x"74712a70",
          1366 => x"81f00670",
          1367 => x"30708025",
          1368 => x"822b8471",
          1369 => x"3174712a",
          1370 => x"5553751b",
          1371 => x"05738c06",
          1372 => x"70307080",
          1373 => x"25108271",
          1374 => x"3177712a",
          1375 => x"70812a81",
          1376 => x"32708106",
          1377 => x"70308274",
          1378 => x"31067519",
          1379 => x"0584b8e4",
          1380 => x"0c515254",
          1381 => x"55515456",
          1382 => x"5a535555",
          1383 => x"55515656",
          1384 => x"56565158",
          1385 => x"56545286",
          1386 => x"3d0d04fd",
          1387 => x"3d0d7577",
          1388 => x"70547153",
          1389 => x"54548194",
          1390 => x"3f84b8e4",
          1391 => x"08732974",
          1392 => x"713184b8",
          1393 => x"e40c5385",
          1394 => x"3d0d04fa",
          1395 => x"3d0d787a",
          1396 => x"5854a053",
          1397 => x"76802e8b",
          1398 => x"387651fe",
          1399 => x"cf3f84b8",
          1400 => x"e40853e0",
          1401 => x"13527380",
          1402 => x"2e8d3873",
          1403 => x"51febd3f",
          1404 => x"7284b8e4",
          1405 => x"08315273",
          1406 => x"53719f26",
          1407 => x"80c53880",
          1408 => x"53719f2e",
          1409 => x"be388112",
          1410 => x"74712aa0",
          1411 => x"72317671",
          1412 => x"2b575454",
          1413 => x"55805674",
          1414 => x"762ea838",
          1415 => x"7210749f",
          1416 => x"2a077410",
          1417 => x"77077872",
          1418 => x"31ff119f",
          1419 => x"2c708106",
          1420 => x"7b720675",
          1421 => x"7131ff1c",
          1422 => x"5c565252",
          1423 => x"55585553",
          1424 => x"74da3872",
          1425 => x"84b8e40c",
          1426 => x"883d0d04",
          1427 => x"fa3d0d78",
          1428 => x"9f2c7a9f",
          1429 => x"2c7a9f2c",
          1430 => x"7b327c9f",
          1431 => x"2c7d3273",
          1432 => x"73327174",
          1433 => x"31577275",
          1434 => x"31565956",
          1435 => x"595556fc",
          1436 => x"b43f84b8",
          1437 => x"e4087532",
          1438 => x"753184b8",
          1439 => x"e40c883d",
          1440 => x"0d04f73d",
          1441 => x"0d7b7d5b",
          1442 => x"5780707b",
          1443 => x"0c770870",
          1444 => x"33565659",
          1445 => x"73a02e09",
          1446 => x"81068f38",
          1447 => x"81157078",
          1448 => x"0c703355",
          1449 => x"5573a02e",
          1450 => x"f33873ad",
          1451 => x"2e80f538",
          1452 => x"73b02e81",
          1453 => x"8338d014",
          1454 => x"58805677",
          1455 => x"892680db",
          1456 => x"388a5880",
          1457 => x"56a07427",
          1458 => x"80c43880",
          1459 => x"e0742789",
          1460 => x"38e01470",
          1461 => x"81ff0655",
          1462 => x"53d01470",
          1463 => x"81ff0651",
          1464 => x"53907327",
          1465 => x"8f38f913",
          1466 => x"7081ff06",
          1467 => x"54548973",
          1468 => x"27818938",
          1469 => x"72782781",
          1470 => x"83387776",
          1471 => x"29138116",
          1472 => x"70790c70",
          1473 => x"33565656",
          1474 => x"73a026ff",
          1475 => x"be387880",
          1476 => x"2e843875",
          1477 => x"3056757a",
          1478 => x"0c815675",
          1479 => x"84b8e40c",
          1480 => x"8b3d0d04",
          1481 => x"81701670",
          1482 => x"790c7033",
          1483 => x"56565973",
          1484 => x"b02e0981",
          1485 => x"06feff38",
          1486 => x"81157078",
          1487 => x"0c703355",
          1488 => x"557380e2",
          1489 => x"2ea63890",
          1490 => x"587380f8",
          1491 => x"2ea03881",
          1492 => x"56a07427",
          1493 => x"c638d014",
          1494 => x"53805688",
          1495 => x"58897327",
          1496 => x"fee13875",
          1497 => x"84b8e40c",
          1498 => x"8b3d0d04",
          1499 => x"82588115",
          1500 => x"70780c70",
          1501 => x"33555580",
          1502 => x"56feca39",
          1503 => x"800b84b8",
          1504 => x"e40c8b3d",
          1505 => x"0d04f73d",
          1506 => x"0d7b7d5b",
          1507 => x"5780707b",
          1508 => x"0c770870",
          1509 => x"33565659",
          1510 => x"73a02e09",
          1511 => x"81068f38",
          1512 => x"81157078",
          1513 => x"0c703355",
          1514 => x"5573a02e",
          1515 => x"f33873ad",
          1516 => x"2e80f538",
          1517 => x"73b02e81",
          1518 => x"8338d014",
          1519 => x"58805677",
          1520 => x"892680db",
          1521 => x"388a5880",
          1522 => x"56a07427",
          1523 => x"80c43880",
          1524 => x"e0742789",
          1525 => x"38e01470",
          1526 => x"81ff0655",
          1527 => x"53d01470",
          1528 => x"81ff0651",
          1529 => x"53907327",
          1530 => x"8f38f913",
          1531 => x"7081ff06",
          1532 => x"54548973",
          1533 => x"27818938",
          1534 => x"72782781",
          1535 => x"83387776",
          1536 => x"29138116",
          1537 => x"70790c70",
          1538 => x"33565656",
          1539 => x"73a026ff",
          1540 => x"be387880",
          1541 => x"2e843875",
          1542 => x"3056757a",
          1543 => x"0c815675",
          1544 => x"84b8e40c",
          1545 => x"8b3d0d04",
          1546 => x"81701670",
          1547 => x"790c7033",
          1548 => x"56565973",
          1549 => x"b02e0981",
          1550 => x"06feff38",
          1551 => x"81157078",
          1552 => x"0c703355",
          1553 => x"557380e2",
          1554 => x"2ea63890",
          1555 => x"587380f8",
          1556 => x"2ea03881",
          1557 => x"56a07427",
          1558 => x"c638d014",
          1559 => x"53805688",
          1560 => x"58897327",
          1561 => x"fee13875",
          1562 => x"84b8e40c",
          1563 => x"8b3d0d04",
          1564 => x"82588115",
          1565 => x"70780c70",
          1566 => x"33555580",
          1567 => x"56feca39",
          1568 => x"800b84b8",
          1569 => x"e40c8b3d",
          1570 => x"0d0480d6",
          1571 => x"d13f84b8",
          1572 => x"e40881ff",
          1573 => x"0684b8e4",
          1574 => x"0c04ff3d",
          1575 => x"0d735271",
          1576 => x"93268c38",
          1577 => x"71101083",
          1578 => x"bdf40552",
          1579 => x"71080483",
          1580 => x"ce8c51ef",
          1581 => x"be3f833d",
          1582 => x"0d0483ce",
          1583 => x"9c51efb3",
          1584 => x"3f833d0d",
          1585 => x"0483ceb4",
          1586 => x"51efa83f",
          1587 => x"833d0d04",
          1588 => x"83cecc51",
          1589 => x"ef9d3f83",
          1590 => x"3d0d0483",
          1591 => x"cee451ef",
          1592 => x"923f833d",
          1593 => x"0d0483ce",
          1594 => x"f451ef87",
          1595 => x"3f833d0d",
          1596 => x"0483cf94",
          1597 => x"51eefc3f",
          1598 => x"833d0d04",
          1599 => x"83cfa451",
          1600 => x"eef13f83",
          1601 => x"3d0d0483",
          1602 => x"cfcc51ee",
          1603 => x"e63f833d",
          1604 => x"0d0483cf",
          1605 => x"e051eedb",
          1606 => x"3f833d0d",
          1607 => x"0483cffc",
          1608 => x"51eed03f",
          1609 => x"833d0d04",
          1610 => x"83d09451",
          1611 => x"eec53f83",
          1612 => x"3d0d0483",
          1613 => x"d0ac51ee",
          1614 => x"ba3f833d",
          1615 => x"0d0483d0",
          1616 => x"c451eeaf",
          1617 => x"3f833d0d",
          1618 => x"0483d0d4",
          1619 => x"51eea43f",
          1620 => x"833d0d04",
          1621 => x"83d0e851",
          1622 => x"ee993f83",
          1623 => x"3d0d0483",
          1624 => x"d0f851ee",
          1625 => x"8e3f833d",
          1626 => x"0d0483d1",
          1627 => x"8851ee83",
          1628 => x"3f833d0d",
          1629 => x"0483d198",
          1630 => x"51edf83f",
          1631 => x"833d0d04",
          1632 => x"83d1a851",
          1633 => x"eded3f83",
          1634 => x"3d0d0483",
          1635 => x"d1b451ed",
          1636 => x"e23f833d",
          1637 => x"0d04ec3d",
          1638 => x"0d660284",
          1639 => x"0580e305",
          1640 => x"335b5880",
          1641 => x"68793070",
          1642 => x"7b077325",
          1643 => x"51575759",
          1644 => x"78577587",
          1645 => x"ff268338",
          1646 => x"81577477",
          1647 => x"077081ff",
          1648 => x"06515593",
          1649 => x"577480e2",
          1650 => x"38815377",
          1651 => x"528c3d70",
          1652 => x"52588295",
          1653 => x"c83f84b8",
          1654 => x"e4085784",
          1655 => x"b8e40880",
          1656 => x"2e80d038",
          1657 => x"775182af",
          1658 => x"863f7630",
          1659 => x"70780780",
          1660 => x"257b3070",
          1661 => x"9f2a7206",
          1662 => x"53575758",
          1663 => x"77802eaa",
          1664 => x"3887c098",
          1665 => x"88085574",
          1666 => x"87e72680",
          1667 => x"e0387452",
          1668 => x"7887e829",
          1669 => x"51f58e3f",
          1670 => x"84b8e408",
          1671 => x"5483d1e4",
          1672 => x"53785283",
          1673 => x"d1c051df",
          1674 => x"df3f7684",
          1675 => x"b8e40c96",
          1676 => x"3d0d0484",
          1677 => x"b8e40887",
          1678 => x"c098880c",
          1679 => x"84b8e408",
          1680 => x"59963dd4",
          1681 => x"05548480",
          1682 => x"53755277",
          1683 => x"51829dbd",
          1684 => x"3f84b8e4",
          1685 => x"085784b8",
          1686 => x"e408ff88",
          1687 => x"387a5574",
          1688 => x"802eff80",
          1689 => x"38741975",
          1690 => x"175759d5",
          1691 => x"3987e852",
          1692 => x"7451f4b1",
          1693 => x"3f84b8e4",
          1694 => x"08527851",
          1695 => x"f4a73f84",
          1696 => x"b8e40854",
          1697 => x"83d1e453",
          1698 => x"785283d1",
          1699 => x"c051def8",
          1700 => x"3fff9739",
          1701 => x"f83d0d7c",
          1702 => x"028405b7",
          1703 => x"05335859",
          1704 => x"ff588053",
          1705 => x"7b527a51",
          1706 => x"fdec3f84",
          1707 => x"b8e4088b",
          1708 => x"3876802e",
          1709 => x"91387681",
          1710 => x"2e8a3877",
          1711 => x"84b8e40c",
          1712 => x"8a3d0d04",
          1713 => x"780484d4",
          1714 => x"c4566155",
          1715 => x"605484b8",
          1716 => x"e4537f52",
          1717 => x"7e51782d",
          1718 => x"84b8e408",
          1719 => x"84b8e40c",
          1720 => x"8a3d0d04",
          1721 => x"f33d0d7f",
          1722 => x"6163028c",
          1723 => x"0580cf05",
          1724 => x"33737315",
          1725 => x"68415f5c",
          1726 => x"5c5f5d5e",
          1727 => x"78802e83",
          1728 => x"82387a52",
          1729 => x"83d1ec51",
          1730 => x"ddfe3f83",
          1731 => x"d1f451dd",
          1732 => x"f73f8054",
          1733 => x"737927b2",
          1734 => x"387c902e",
          1735 => x"81ed387c",
          1736 => x"a02e82a8",
          1737 => x"38731853",
          1738 => x"727a2781",
          1739 => x"a7387233",
          1740 => x"5283d1f8",
          1741 => x"51ddd13f",
          1742 => x"811484d4",
          1743 => x"c8085354",
          1744 => x"a051ecaa",
          1745 => x"3f787426",
          1746 => x"dc3883d2",
          1747 => x"8051ddb8",
          1748 => x"3f805675",
          1749 => x"792780c0",
          1750 => x"38751870",
          1751 => x"33555380",
          1752 => x"55727a27",
          1753 => x"83388155",
          1754 => x"80539f74",
          1755 => x"27833881",
          1756 => x"53747306",
          1757 => x"7081ff06",
          1758 => x"56577480",
          1759 => x"2e883880",
          1760 => x"fe742781",
          1761 => x"ee3884d4",
          1762 => x"c80852a0",
          1763 => x"51ebdf3f",
          1764 => x"81165678",
          1765 => x"7626c238",
          1766 => x"83d28451",
          1767 => x"e9d53f78",
          1768 => x"18791c5c",
          1769 => x"5880519d",
          1770 => x"a83f84b8",
          1771 => x"e408982b",
          1772 => x"70982c58",
          1773 => x"5476a02e",
          1774 => x"81ee3876",
          1775 => x"9b2e82c3",
          1776 => x"387b1e57",
          1777 => x"767826fe",
          1778 => x"b938ff0b",
          1779 => x"84b8e40c",
          1780 => x"8f3d0d04",
          1781 => x"83d28851",
          1782 => x"dcae3f81",
          1783 => x"1484d4c8",
          1784 => x"085354a0",
          1785 => x"51eb873f",
          1786 => x"787426fe",
          1787 => x"b838feda",
          1788 => x"3983d298",
          1789 => x"51dc913f",
          1790 => x"821484d4",
          1791 => x"c8085354",
          1792 => x"a051eaea",
          1793 => x"3f737927",
          1794 => x"fec03873",
          1795 => x"1853727a",
          1796 => x"27df3872",
          1797 => x"225283d2",
          1798 => x"8c51dbec",
          1799 => x"3f821484",
          1800 => x"d4c80853",
          1801 => x"54a051ea",
          1802 => x"c53f7874",
          1803 => x"26dd38fe",
          1804 => x"993983d2",
          1805 => x"9451dbd0",
          1806 => x"3f841484",
          1807 => x"d4c80853",
          1808 => x"54a051ea",
          1809 => x"a93f7379",
          1810 => x"27fdff38",
          1811 => x"73185372",
          1812 => x"7a27df38",
          1813 => x"72085283",
          1814 => x"d1ec51db",
          1815 => x"ab3f8414",
          1816 => x"84d4c808",
          1817 => x"5354a051",
          1818 => x"ea843f78",
          1819 => x"7426dd38",
          1820 => x"fdd83984",
          1821 => x"d4c80852",
          1822 => x"7351e9f2",
          1823 => x"3f811656",
          1824 => x"fe913980",
          1825 => x"ced83f84",
          1826 => x"b8e40881",
          1827 => x"ff065388",
          1828 => x"5972a82e",
          1829 => x"fcec38a0",
          1830 => x"597280d0",
          1831 => x"2e098106",
          1832 => x"fce03890",
          1833 => x"59fcdb39",
          1834 => x"80519ba5",
          1835 => x"3f84b8e4",
          1836 => x"08982b70",
          1837 => x"982c70a0",
          1838 => x"32703072",
          1839 => x"9b327030",
          1840 => x"70720773",
          1841 => x"75070651",
          1842 => x"55585957",
          1843 => x"58537280",
          1844 => x"25fde838",
          1845 => x"80519af9",
          1846 => x"3f84b8e4",
          1847 => x"08982b70",
          1848 => x"982c70a0",
          1849 => x"32703072",
          1850 => x"9b327030",
          1851 => x"70720773",
          1852 => x"75070651",
          1853 => x"55585957",
          1854 => x"58538073",
          1855 => x"24ffa938",
          1856 => x"fdb93980",
          1857 => x"0b84b8e4",
          1858 => x"0c8f3d0d",
          1859 => x"04fe3d0d",
          1860 => x"87c09680",
          1861 => x"0853aac7",
          1862 => x"3f81519c",
          1863 => x"ed3f83d2",
          1864 => x"dc519cfe",
          1865 => x"3f80519c",
          1866 => x"e13f7281",
          1867 => x"2a708106",
          1868 => x"51527182",
          1869 => x"b7387282",
          1870 => x"2a708106",
          1871 => x"51527182",
          1872 => x"89387283",
          1873 => x"2a708106",
          1874 => x"51527181",
          1875 => x"db387284",
          1876 => x"2a708106",
          1877 => x"51527181",
          1878 => x"ad387285",
          1879 => x"2a708106",
          1880 => x"51527180",
          1881 => x"ff387286",
          1882 => x"2a708106",
          1883 => x"51527180",
          1884 => x"d2387287",
          1885 => x"2a708106",
          1886 => x"515271a9",
          1887 => x"3872882a",
          1888 => x"81065372",
          1889 => x"8838a9df",
          1890 => x"3f843d0d",
          1891 => x"0481519b",
          1892 => x"f93f83d2",
          1893 => x"f4519c8a",
          1894 => x"3f80519b",
          1895 => x"ed3fa9c7",
          1896 => x"3f843d0d",
          1897 => x"0481519b",
          1898 => x"e13f83d3",
          1899 => x"88519bf2",
          1900 => x"3f80519b",
          1901 => x"d53f7288",
          1902 => x"2a810653",
          1903 => x"72802ec6",
          1904 => x"38cb3981",
          1905 => x"519bc33f",
          1906 => x"83d39c51",
          1907 => x"9bd43f80",
          1908 => x"519bb73f",
          1909 => x"72872a70",
          1910 => x"81065152",
          1911 => x"71802eff",
          1912 => x"9c38c239",
          1913 => x"81519ba2",
          1914 => x"3f83d3b0",
          1915 => x"519bb33f",
          1916 => x"80519b96",
          1917 => x"3f72862a",
          1918 => x"70810651",
          1919 => x"5271802e",
          1920 => x"fef038ff",
          1921 => x"be398151",
          1922 => x"9b803f83",
          1923 => x"d3c4519b",
          1924 => x"913f8051",
          1925 => x"9af43f72",
          1926 => x"852a7081",
          1927 => x"06515271",
          1928 => x"802efec2",
          1929 => x"38ffbd39",
          1930 => x"81519ade",
          1931 => x"3f83d3d8",
          1932 => x"519aef3f",
          1933 => x"80519ad2",
          1934 => x"3f72842a",
          1935 => x"70810651",
          1936 => x"5271802e",
          1937 => x"fe9438ff",
          1938 => x"bd398151",
          1939 => x"9abc3f83",
          1940 => x"d3ec519a",
          1941 => x"cd3f8051",
          1942 => x"9ab03f72",
          1943 => x"832a7081",
          1944 => x"06515271",
          1945 => x"802efde6",
          1946 => x"38ffbd39",
          1947 => x"81519a9a",
          1948 => x"3f83d3fc",
          1949 => x"519aab3f",
          1950 => x"80519a8e",
          1951 => x"3f72822a",
          1952 => x"70810651",
          1953 => x"5271802e",
          1954 => x"fdb838ff",
          1955 => x"bd39ca3d",
          1956 => x"0d807041",
          1957 => x"41ff6184",
          1958 => x"cff00c42",
          1959 => x"81526051",
          1960 => x"81b5fb3f",
          1961 => x"84b8e408",
          1962 => x"81ff069b",
          1963 => x"3d405978",
          1964 => x"612e84b1",
          1965 => x"3883d4d0",
          1966 => x"51e3b83f",
          1967 => x"983d4383",
          1968 => x"d58851d6",
          1969 => x"c33f7e48",
          1970 => x"80f85380",
          1971 => x"527e51eb",
          1972 => x"ae3f0b0b",
          1973 => x"83edd833",
          1974 => x"7081ff06",
          1975 => x"5b597980",
          1976 => x"2e82f138",
          1977 => x"79812e83",
          1978 => x"88387881",
          1979 => x"ff065e7d",
          1980 => x"822e83c1",
          1981 => x"3867705a",
          1982 => x"5a79802e",
          1983 => x"83dc3879",
          1984 => x"335c7ba0",
          1985 => x"2e098106",
          1986 => x"8c38811a",
          1987 => x"70335d5a",
          1988 => x"7ba02ef6",
          1989 => x"38805c7b",
          1990 => x"9b26be38",
          1991 => x"7b902983",
          1992 => x"eddc0570",
          1993 => x"08525be7",
          1994 => x"ff3f84b8",
          1995 => x"e40884b8",
          1996 => x"e408547a",
          1997 => x"537b0852",
          1998 => x"5de8da3f",
          1999 => x"84b8e408",
          2000 => x"8b38841b",
          2001 => x"335e7d81",
          2002 => x"2e838038",
          2003 => x"811c7081",
          2004 => x"ff065d5b",
          2005 => x"9b7c27c4",
          2006 => x"389a3d33",
          2007 => x"5c7b802e",
          2008 => x"fedd3880",
          2009 => x"f8527e51",
          2010 => x"e9923f84",
          2011 => x"b8e4085e",
          2012 => x"84b8e408",
          2013 => x"802e8dc9",
          2014 => x"3884b8e4",
          2015 => x"0848b83d",
          2016 => x"ff800551",
          2017 => x"91893f84",
          2018 => x"b8e40860",
          2019 => x"62065c5c",
          2020 => x"7a802e81",
          2021 => x"843884b8",
          2022 => x"e40851e7",
          2023 => x"8b3f84b8",
          2024 => x"e4088f26",
          2025 => x"80f33881",
          2026 => x"0ba53d5e",
          2027 => x"5b7a822e",
          2028 => x"8d85387a",
          2029 => x"82248ce2",
          2030 => x"387a812e",
          2031 => x"82e4387b",
          2032 => x"54805383",
          2033 => x"d58c527c",
          2034 => x"51d5dd3f",
          2035 => x"83f1a058",
          2036 => x"84b99457",
          2037 => x"7d566755",
          2038 => x"80549080",
          2039 => x"0a539080",
          2040 => x"0a527c51",
          2041 => x"f5ae3f84",
          2042 => x"b8e40884",
          2043 => x"b8e40809",
          2044 => x"70307072",
          2045 => x"07802551",
          2046 => x"5b5b4280",
          2047 => x"5a7a8326",
          2048 => x"8338815a",
          2049 => x"787a0659",
          2050 => x"78802e8d",
          2051 => x"38811b70",
          2052 => x"81ff065c",
          2053 => x"5a7aff95",
          2054 => x"387f8132",
          2055 => x"61813207",
          2056 => x"5d7c81ee",
          2057 => x"3861ff2e",
          2058 => x"81e8387d",
          2059 => x"518194d0",
          2060 => x"3f83d588",
          2061 => x"51d3d13f",
          2062 => x"7e4880f8",
          2063 => x"5380527e",
          2064 => x"51e8bc3f",
          2065 => x"0b0b83ed",
          2066 => x"d8337081",
          2067 => x"ff065b59",
          2068 => x"79fd9138",
          2069 => x"815383d4",
          2070 => x"b45284cf",
          2071 => x"f4518288",
          2072 => x"bc3f84b8",
          2073 => x"e40880c5",
          2074 => x"38810b0b",
          2075 => x"0b83edd8",
          2076 => x"3484cff4",
          2077 => x"5380f852",
          2078 => x"7e5182f6",
          2079 => x"b73f84b8",
          2080 => x"e408802e",
          2081 => x"a03884b8",
          2082 => x"e40851df",
          2083 => x"e63f0b0b",
          2084 => x"83edd833",
          2085 => x"7081ff06",
          2086 => x"5f597d82",
          2087 => x"2e098106",
          2088 => x"fcd33891",
          2089 => x"3984cff4",
          2090 => x"5182a1c3",
          2091 => x"3f820b0b",
          2092 => x"0b83edd8",
          2093 => x"3483d4c4",
          2094 => x"5380f852",
          2095 => x"7e51a7c3",
          2096 => x"3f67705a",
          2097 => x"5a79fcb7",
          2098 => x"3890397c",
          2099 => x"1a630c85",
          2100 => x"1b335978",
          2101 => x"818926fd",
          2102 => x"80387810",
          2103 => x"1083bec4",
          2104 => x"055a7908",
          2105 => x"04835383",
          2106 => x"d594527e",
          2107 => x"51e4fb3f",
          2108 => x"60537e52",
          2109 => x"84ba9051",
          2110 => x"8284f33f",
          2111 => x"84b8e408",
          2112 => x"612e0981",
          2113 => x"06fbae38",
          2114 => x"81709a3d",
          2115 => x"454141fb",
          2116 => x"ae3983d5",
          2117 => x"9851dedb",
          2118 => x"3f7d5181",
          2119 => x"92e23ffe",
          2120 => x"903983d5",
          2121 => x"a8567b55",
          2122 => x"83d5ac54",
          2123 => x"805383d5",
          2124 => x"b0527c51",
          2125 => x"d2f23ffd",
          2126 => x"9339818c",
          2127 => x"9a3ffaff",
          2128 => x"399add3f",
          2129 => x"faf93981",
          2130 => x"528351bf",
          2131 => x"933ffaef",
          2132 => x"39818dc5",
          2133 => x"3ffae839",
          2134 => x"83d5c051",
          2135 => x"de953f80",
          2136 => x"59780483",
          2137 => x"d5d451de",
          2138 => x"8a3fd0fd",
          2139 => x"3ffad039",
          2140 => x"b83dff84",
          2141 => x"1153ff80",
          2142 => x"0551ec8a",
          2143 => x"3f84b8e4",
          2144 => x"08802efa",
          2145 => x"ba386852",
          2146 => x"83d5f051",
          2147 => x"d0fa3f68",
          2148 => x"5a792d84",
          2149 => x"b8e40880",
          2150 => x"2efaa438",
          2151 => x"84b8e408",
          2152 => x"5283d68c",
          2153 => x"51d0e13f",
          2154 => x"fa9539b8",
          2155 => x"3dff8411",
          2156 => x"53ff8005",
          2157 => x"51ebcf3f",
          2158 => x"84b8e408",
          2159 => x"802ef9ff",
          2160 => x"38685283",
          2161 => x"d6a851d0",
          2162 => x"bf3f6859",
          2163 => x"7804b83d",
          2164 => x"fef41153",
          2165 => x"ff800551",
          2166 => x"e9a83f84",
          2167 => x"b8e40880",
          2168 => x"2ef9dc38",
          2169 => x"b83dfef0",
          2170 => x"1153ff80",
          2171 => x"0551e992",
          2172 => x"3f84b8e4",
          2173 => x"0886d038",
          2174 => x"64597808",
          2175 => x"53785283",
          2176 => x"d6c451d0",
          2177 => x"833f84d4",
          2178 => x"c4085380",
          2179 => x"f8527e51",
          2180 => x"d0913f7e",
          2181 => x"487e3359",
          2182 => x"78ae2ef9",
          2183 => x"a238789f",
          2184 => x"2687d338",
          2185 => x"64840570",
          2186 => x"4659cf39",
          2187 => x"b83dfef4",
          2188 => x"1153ff80",
          2189 => x"0551e8ca",
          2190 => x"3f84b8e4",
          2191 => x"08802ef8",
          2192 => x"fe38b83d",
          2193 => x"fef01153",
          2194 => x"ff800551",
          2195 => x"e8b43f84",
          2196 => x"b8e40886",
          2197 => x"b0386459",
          2198 => x"78225378",
          2199 => x"5283d6d4",
          2200 => x"51cfa53f",
          2201 => x"84d4c408",
          2202 => x"5380f852",
          2203 => x"7e51cfb3",
          2204 => x"3f7e487e",
          2205 => x"335978ae",
          2206 => x"2ef8c438",
          2207 => x"789f2687",
          2208 => x"ca386482",
          2209 => x"05704659",
          2210 => x"cf39b83d",
          2211 => x"ff841153",
          2212 => x"ff800551",
          2213 => x"e9f03f84",
          2214 => x"b8e40880",
          2215 => x"2ef8a038",
          2216 => x"b83dfefc",
          2217 => x"1153ff80",
          2218 => x"0551e9da",
          2219 => x"3f84b8e4",
          2220 => x"08802ef8",
          2221 => x"8a38b83d",
          2222 => x"fef81153",
          2223 => x"ff800551",
          2224 => x"e9c43f84",
          2225 => x"b8e40880",
          2226 => x"2ef7f438",
          2227 => x"83d6e051",
          2228 => x"ceb63f68",
          2229 => x"675d5978",
          2230 => x"7c27838d",
          2231 => x"38657033",
          2232 => x"7a335f5c",
          2233 => x"5a7a7d2e",
          2234 => x"95387a55",
          2235 => x"79547833",
          2236 => x"53785283",
          2237 => x"d6f051ce",
          2238 => x"8f3f6666",
          2239 => x"5b5c8119",
          2240 => x"811b4759",
          2241 => x"d239b83d",
          2242 => x"ff841153",
          2243 => x"ff800551",
          2244 => x"e8f43f84",
          2245 => x"b8e40880",
          2246 => x"2ef7a438",
          2247 => x"b83dfefc",
          2248 => x"1153ff80",
          2249 => x"0551e8de",
          2250 => x"3f84b8e4",
          2251 => x"08802ef7",
          2252 => x"8e38b83d",
          2253 => x"fef81153",
          2254 => x"ff800551",
          2255 => x"e8c83f84",
          2256 => x"b8e40880",
          2257 => x"2ef6f838",
          2258 => x"83d78c51",
          2259 => x"cdba3f68",
          2260 => x"5a796727",
          2261 => x"82933865",
          2262 => x"5c797081",
          2263 => x"055b337c",
          2264 => x"34658105",
          2265 => x"46eb39b8",
          2266 => x"3dff8411",
          2267 => x"53ff8005",
          2268 => x"51e8933f",
          2269 => x"84b8e408",
          2270 => x"802ef6c3",
          2271 => x"38b83dfe",
          2272 => x"fc1153ff",
          2273 => x"800551e7",
          2274 => x"fd3f84b8",
          2275 => x"e408b138",
          2276 => x"68703354",
          2277 => x"5283d798",
          2278 => x"51cced3f",
          2279 => x"84d4c408",
          2280 => x"5380f852",
          2281 => x"7e51ccfb",
          2282 => x"3f7e487e",
          2283 => x"335978ae",
          2284 => x"2ef68c38",
          2285 => x"789f2684",
          2286 => x"97386881",
          2287 => x"0549d139",
          2288 => x"68590280",
          2289 => x"db053379",
          2290 => x"34688105",
          2291 => x"49b83dfe",
          2292 => x"fc1153ff",
          2293 => x"800551e7",
          2294 => x"ad3f84b8",
          2295 => x"e408802e",
          2296 => x"f5dd3868",
          2297 => x"590280db",
          2298 => x"05337934",
          2299 => x"68810549",
          2300 => x"b83dfefc",
          2301 => x"1153ff80",
          2302 => x"0551e78a",
          2303 => x"3f84b8e4",
          2304 => x"08ffbd38",
          2305 => x"f5b939b8",
          2306 => x"3dff8411",
          2307 => x"53ff8005",
          2308 => x"51e6f33f",
          2309 => x"84b8e408",
          2310 => x"802ef5a3",
          2311 => x"38b83dfe",
          2312 => x"fc1153ff",
          2313 => x"800551e6",
          2314 => x"dd3f84b8",
          2315 => x"e408802e",
          2316 => x"f58d38b8",
          2317 => x"3dfef811",
          2318 => x"53ff8005",
          2319 => x"51e6c73f",
          2320 => x"84b8e408",
          2321 => x"863884b8",
          2322 => x"e4084683",
          2323 => x"d7a451cb",
          2324 => x"b73f6867",
          2325 => x"5b59787a",
          2326 => x"278f3865",
          2327 => x"5b7a7970",
          2328 => x"84055b0c",
          2329 => x"797926f5",
          2330 => x"388a51d9",
          2331 => x"f13ff4cf",
          2332 => x"39b83dff",
          2333 => x"80055187",
          2334 => x"963f84b8",
          2335 => x"e408b93d",
          2336 => x"ff800552",
          2337 => x"5988d83f",
          2338 => x"815384b8",
          2339 => x"e4085278",
          2340 => x"51ea833f",
          2341 => x"84b8e408",
          2342 => x"802ef4a3",
          2343 => x"3884b8e4",
          2344 => x"0851e7f6",
          2345 => x"3ff49839",
          2346 => x"b83dff84",
          2347 => x"1153ff80",
          2348 => x"0551e5d2",
          2349 => x"3f84b8e4",
          2350 => x"08913883",
          2351 => x"f1e8335a",
          2352 => x"79802e83",
          2353 => x"c03883f1",
          2354 => x"a00849b8",
          2355 => x"3dfefc11",
          2356 => x"53ff8005",
          2357 => x"51e5af3f",
          2358 => x"84b8e408",
          2359 => x"913883f1",
          2360 => x"e8335a79",
          2361 => x"802e838a",
          2362 => x"3883f1a4",
          2363 => x"0847b83d",
          2364 => x"fef81153",
          2365 => x"ff800551",
          2366 => x"e58c3f84",
          2367 => x"b8e40880",
          2368 => x"2ea53880",
          2369 => x"665c5c7a",
          2370 => x"882e8338",
          2371 => x"815c7a90",
          2372 => x"32703070",
          2373 => x"72079f2a",
          2374 => x"7e065c5f",
          2375 => x"5d79802e",
          2376 => x"88387aa0",
          2377 => x"2e833888",
          2378 => x"4683d7b4",
          2379 => x"51d6c43f",
          2380 => x"80556854",
          2381 => x"65536652",
          2382 => x"6851eba8",
          2383 => x"3f83d7c0",
          2384 => x"51d6b03f",
          2385 => x"f2f93964",
          2386 => x"64710c59",
          2387 => x"64840545",
          2388 => x"b83dfef0",
          2389 => x"1153ff80",
          2390 => x"0551e2a6",
          2391 => x"3f84b8e4",
          2392 => x"08802ef2",
          2393 => x"da386464",
          2394 => x"710c5964",
          2395 => x"840545b8",
          2396 => x"3dfef011",
          2397 => x"53ff8005",
          2398 => x"51e2873f",
          2399 => x"84b8e408",
          2400 => x"c638f2bb",
          2401 => x"39645e02",
          2402 => x"80ce0522",
          2403 => x"7e708205",
          2404 => x"40237d45",
          2405 => x"b83dfef0",
          2406 => x"1153ff80",
          2407 => x"0551e1e2",
          2408 => x"3f84b8e4",
          2409 => x"08802ef2",
          2410 => x"9638645e",
          2411 => x"0280ce05",
          2412 => x"227e7082",
          2413 => x"0540237d",
          2414 => x"45b83dfe",
          2415 => x"f01153ff",
          2416 => x"800551e1",
          2417 => x"bd3f84b8",
          2418 => x"e408ffb9",
          2419 => x"38f1f039",
          2420 => x"b83dfefc",
          2421 => x"1153ff80",
          2422 => x"0551e3aa",
          2423 => x"3f84b8e4",
          2424 => x"08802e81",
          2425 => x"dc38685c",
          2426 => x"0280db05",
          2427 => x"337c3468",
          2428 => x"810549fb",
          2429 => x"9b39b83d",
          2430 => x"fef01153",
          2431 => x"ff800551",
          2432 => x"e1803f84",
          2433 => x"b8e40880",
          2434 => x"2e819838",
          2435 => x"6464710c",
          2436 => x"5d648405",
          2437 => x"704659f7",
          2438 => x"e1397a83",
          2439 => x"2e098106",
          2440 => x"f39d387b",
          2441 => x"5583d5ac",
          2442 => x"54805383",
          2443 => x"d7cc527c",
          2444 => x"51c8f53f",
          2445 => x"f396397b",
          2446 => x"527c51da",
          2447 => x"8a3ff38c",
          2448 => x"3983d7d8",
          2449 => x"51d4ac3f",
          2450 => x"f0f539b8",
          2451 => x"3dfef011",
          2452 => x"53ff8005",
          2453 => x"51e0ab3f",
          2454 => x"84b8e408",
          2455 => x"802eb838",
          2456 => x"64590280",
          2457 => x"ce052279",
          2458 => x"7082055b",
          2459 => x"237845f7",
          2460 => x"e73983f1",
          2461 => x"e9335c7b",
          2462 => x"802e80cf",
          2463 => x"3883f1ac",
          2464 => x"0847fcea",
          2465 => x"3983f1e9",
          2466 => x"335c7b80",
          2467 => x"2ea13883",
          2468 => x"f1a80849",
          2469 => x"fcb53983",
          2470 => x"d88451d3",
          2471 => x"d63f6459",
          2472 => x"f7b63983",
          2473 => x"d88451d3",
          2474 => x"ca3f6459",
          2475 => x"f6cc3983",
          2476 => x"f1ea3359",
          2477 => x"78802ea5",
          2478 => x"3883f1b0",
          2479 => x"0849fc8b",
          2480 => x"3983d884",
          2481 => x"51d3ac3f",
          2482 => x"f9c63983",
          2483 => x"f1ea3359",
          2484 => x"78802e9b",
          2485 => x"3883f1b4",
          2486 => x"0847fc92",
          2487 => x"3983f1eb",
          2488 => x"335e7d80",
          2489 => x"2e9b3883",
          2490 => x"f1b80849",
          2491 => x"fbdd3983",
          2492 => x"f1eb335e",
          2493 => x"7d802e9b",
          2494 => x"3883f1bc",
          2495 => x"0847fbee",
          2496 => x"3983f1e6",
          2497 => x"335d7c80",
          2498 => x"2e9b3883",
          2499 => x"f1c00849",
          2500 => x"fbb93983",
          2501 => x"f1e6335d",
          2502 => x"7c802e94",
          2503 => x"3883f1c4",
          2504 => x"0847fbca",
          2505 => x"3983f1d0",
          2506 => x"08fc8005",
          2507 => x"49fb9c39",
          2508 => x"83f1d008",
          2509 => x"880547fb",
          2510 => x"b539f33d",
          2511 => x"0d800b84",
          2512 => x"b9943487",
          2513 => x"c0948c70",
          2514 => x"08565787",
          2515 => x"84805274",
          2516 => x"51dad23f",
          2517 => x"84b8e408",
          2518 => x"902b7708",
          2519 => x"57558784",
          2520 => x"80527551",
          2521 => x"dabf3f74",
          2522 => x"84b8e408",
          2523 => x"07770c87",
          2524 => x"c0949c70",
          2525 => x"08565787",
          2526 => x"84805274",
          2527 => x"51daa63f",
          2528 => x"84b8e408",
          2529 => x"902b7708",
          2530 => x"57558784",
          2531 => x"80527551",
          2532 => x"da933f74",
          2533 => x"84b8e408",
          2534 => x"07770c8c",
          2535 => x"80830b87",
          2536 => x"c094840c",
          2537 => x"8c80830b",
          2538 => x"87c09494",
          2539 => x"0c81bce1",
          2540 => x"5c81c7e0",
          2541 => x"5d830284",
          2542 => x"05a10534",
          2543 => x"805e84d4",
          2544 => x"c40b893d",
          2545 => x"7088130c",
          2546 => x"70720c84",
          2547 => x"d4c80c56",
          2548 => x"b6f43f89",
          2549 => x"833f9587",
          2550 => x"3fba8d51",
          2551 => x"94fc3f83",
          2552 => x"d2a05283",
          2553 => x"d2a451c4",
          2554 => x"9f3f83f1",
          2555 => x"d4702252",
          2556 => x"5594873f",
          2557 => x"83d2ac54",
          2558 => x"83d2b853",
          2559 => x"81153352",
          2560 => x"83d2c051",
          2561 => x"c4823f8d",
          2562 => x"973fed82",
          2563 => x"3f8004fb",
          2564 => x"3d0d7770",
          2565 => x"08565680",
          2566 => x"75525374",
          2567 => x"732e8183",
          2568 => x"38743370",
          2569 => x"81ff0652",
          2570 => x"5270a02e",
          2571 => x"09810691",
          2572 => x"38811570",
          2573 => x"337081ff",
          2574 => x"06535355",
          2575 => x"70a02ef1",
          2576 => x"387181ff",
          2577 => x"065473a2",
          2578 => x"2e818238",
          2579 => x"74527281",
          2580 => x"2e80e738",
          2581 => x"80723370",
          2582 => x"81ff0653",
          2583 => x"545470a0",
          2584 => x"2e833881",
          2585 => x"5470802e",
          2586 => x"8b387380",
          2587 => x"2e863881",
          2588 => x"1252e139",
          2589 => x"807381ff",
          2590 => x"06525470",
          2591 => x"a02e0981",
          2592 => x"06833881",
          2593 => x"5470a232",
          2594 => x"70307080",
          2595 => x"25760752",
          2596 => x"52537280",
          2597 => x"2e883880",
          2598 => x"72708105",
          2599 => x"54347176",
          2600 => x"0c745170",
          2601 => x"84b8e40c",
          2602 => x"873d0d04",
          2603 => x"70802ec4",
          2604 => x"3873802e",
          2605 => x"ffbe3881",
          2606 => x"12528072",
          2607 => x"337081ff",
          2608 => x"06535454",
          2609 => x"70a22ee4",
          2610 => x"388154e0",
          2611 => x"39811555",
          2612 => x"81755353",
          2613 => x"72812e09",
          2614 => x"8106fef8",
          2615 => x"38dc39fc",
          2616 => x"3d0d7653",
          2617 => x"72088b38",
          2618 => x"800b84b8",
          2619 => x"e40c863d",
          2620 => x"0d04863d",
          2621 => x"fc055272",
          2622 => x"51db873f",
          2623 => x"84b8e408",
          2624 => x"802ee538",
          2625 => x"7484b8e4",
          2626 => x"0c863d0d",
          2627 => x"04fc3d0d",
          2628 => x"76821133",
          2629 => x"ff055253",
          2630 => x"8152708b",
          2631 => x"26819838",
          2632 => x"831333ff",
          2633 => x"05548252",
          2634 => x"739e2681",
          2635 => x"8a388413",
          2636 => x"33518352",
          2637 => x"70972680",
          2638 => x"fe388513",
          2639 => x"33548452",
          2640 => x"73bb2680",
          2641 => x"f2388613",
          2642 => x"33558552",
          2643 => x"74bb2680",
          2644 => x"e6388813",
          2645 => x"22558652",
          2646 => x"7487e726",
          2647 => x"80d9388a",
          2648 => x"13225487",
          2649 => x"527387e7",
          2650 => x"2680cc38",
          2651 => x"810b87c0",
          2652 => x"989c0c72",
          2653 => x"2287c098",
          2654 => x"bc0c8213",
          2655 => x"3387c098",
          2656 => x"b80c8313",
          2657 => x"3387c098",
          2658 => x"b40c8413",
          2659 => x"3387c098",
          2660 => x"b00c8513",
          2661 => x"3387c098",
          2662 => x"ac0c8613",
          2663 => x"3387c098",
          2664 => x"a80c7487",
          2665 => x"c098a40c",
          2666 => x"7387c098",
          2667 => x"a00c800b",
          2668 => x"87c0989c",
          2669 => x"0c805271",
          2670 => x"84b8e40c",
          2671 => x"863d0d04",
          2672 => x"f33d0d7f",
          2673 => x"5b87c098",
          2674 => x"9c5d817d",
          2675 => x"0c87c098",
          2676 => x"bc085e7d",
          2677 => x"7b2387c0",
          2678 => x"98b8085c",
          2679 => x"7b821c34",
          2680 => x"87c098b4",
          2681 => x"085a7983",
          2682 => x"1c3487c0",
          2683 => x"98b0085c",
          2684 => x"7b841c34",
          2685 => x"87c098ac",
          2686 => x"085a7985",
          2687 => x"1c3487c0",
          2688 => x"98a8085c",
          2689 => x"7b861c34",
          2690 => x"87c098a4",
          2691 => x"085c7b88",
          2692 => x"1c2387c0",
          2693 => x"98a0085a",
          2694 => x"798a1c23",
          2695 => x"807d0c79",
          2696 => x"83ffff06",
          2697 => x"597b83ff",
          2698 => x"ff065886",
          2699 => x"1b335785",
          2700 => x"1b335684",
          2701 => x"1b335583",
          2702 => x"1b335482",
          2703 => x"1b33537d",
          2704 => x"83ffff06",
          2705 => x"5283d888",
          2706 => x"51ffbfbc",
          2707 => x"3f8f3d0d",
          2708 => x"04fe3d0d",
          2709 => x"02930533",
          2710 => x"5372812e",
          2711 => x"a8387251",
          2712 => x"80e8b03f",
          2713 => x"84b8e408",
          2714 => x"982b7098",
          2715 => x"2c515271",
          2716 => x"ff2e0981",
          2717 => x"06863872",
          2718 => x"832ee338",
          2719 => x"7184b8e4",
          2720 => x"0c843d0d",
          2721 => x"04725180",
          2722 => x"e8893f84",
          2723 => x"b8e40898",
          2724 => x"2b70982c",
          2725 => x"515271ff",
          2726 => x"2e098106",
          2727 => x"df387251",
          2728 => x"80e7f03f",
          2729 => x"84b8e408",
          2730 => x"982b7098",
          2731 => x"2c515271",
          2732 => x"ff2ed238",
          2733 => x"c739fd3d",
          2734 => x"0d807054",
          2735 => x"5271882b",
          2736 => x"54815180",
          2737 => x"e7cd3f84",
          2738 => x"b8e40898",
          2739 => x"2b70982c",
          2740 => x"515271ff",
          2741 => x"2eeb3873",
          2742 => x"72078114",
          2743 => x"54528373",
          2744 => x"25db3871",
          2745 => x"84b8e40c",
          2746 => x"853d0d04",
          2747 => x"fc3d0d02",
          2748 => x"9b053383",
          2749 => x"f19c3370",
          2750 => x"81ff0653",
          2751 => x"55557080",
          2752 => x"2e80f438",
          2753 => x"87c09494",
          2754 => x"0870962a",
          2755 => x"70810653",
          2756 => x"54527080",
          2757 => x"2e8c3871",
          2758 => x"912a7081",
          2759 => x"06515170",
          2760 => x"e3387281",
          2761 => x"32810653",
          2762 => x"72802e8a",
          2763 => x"3871932a",
          2764 => x"81065271",
          2765 => x"cf387381",
          2766 => x"ff065187",
          2767 => x"c0948052",
          2768 => x"70802e86",
          2769 => x"3887c094",
          2770 => x"90527472",
          2771 => x"0c7484b8",
          2772 => x"e40c863d",
          2773 => x"0d047191",
          2774 => x"2a708106",
          2775 => x"51517097",
          2776 => x"38728132",
          2777 => x"81065372",
          2778 => x"802ecb38",
          2779 => x"71932a81",
          2780 => x"06527180",
          2781 => x"2ec03887",
          2782 => x"c0948408",
          2783 => x"70962a70",
          2784 => x"81065354",
          2785 => x"5270cf38",
          2786 => x"d839ff3d",
          2787 => x"0d028f05",
          2788 => x"33703070",
          2789 => x"9f2a5152",
          2790 => x"527083f1",
          2791 => x"9c34833d",
          2792 => x"0d04fa3d",
          2793 => x"0d785580",
          2794 => x"75337056",
          2795 => x"52577077",
          2796 => x"2e80e738",
          2797 => x"811583f1",
          2798 => x"9c337081",
          2799 => x"ff065457",
          2800 => x"5571802e",
          2801 => x"80ff3887",
          2802 => x"c0949408",
          2803 => x"70962a70",
          2804 => x"81065354",
          2805 => x"5270802e",
          2806 => x"8c387191",
          2807 => x"2a708106",
          2808 => x"515170e3",
          2809 => x"38728132",
          2810 => x"81065372",
          2811 => x"802e8a38",
          2812 => x"71932a81",
          2813 => x"065271cf",
          2814 => x"387581ff",
          2815 => x"065187c0",
          2816 => x"94805270",
          2817 => x"802e8638",
          2818 => x"87c09490",
          2819 => x"5273720c",
          2820 => x"81177533",
          2821 => x"555773ff",
          2822 => x"9b387684",
          2823 => x"b8e40c88",
          2824 => x"3d0d0471",
          2825 => x"912a7081",
          2826 => x"06515170",
          2827 => x"98387281",
          2828 => x"32810653",
          2829 => x"72802ec1",
          2830 => x"3871932a",
          2831 => x"81065271",
          2832 => x"802effb5",
          2833 => x"3887c094",
          2834 => x"84087096",
          2835 => x"2a708106",
          2836 => x"53545270",
          2837 => x"ce38d739",
          2838 => x"ff3d0d87",
          2839 => x"c09e8008",
          2840 => x"709c2a8a",
          2841 => x"06525270",
          2842 => x"802e84ab",
          2843 => x"3887c09e",
          2844 => x"a40883f1",
          2845 => x"a00c87c0",
          2846 => x"9ea80883",
          2847 => x"f1a40c87",
          2848 => x"c09e9408",
          2849 => x"83f1a80c",
          2850 => x"87c09e98",
          2851 => x"0883f1ac",
          2852 => x"0c87c09e",
          2853 => x"9c0883f1",
          2854 => x"b00c87c0",
          2855 => x"9ea00883",
          2856 => x"f1b40c87",
          2857 => x"c09eac08",
          2858 => x"83f1b80c",
          2859 => x"87c09eb0",
          2860 => x"0883f1bc",
          2861 => x"0c87c09e",
          2862 => x"b40883f1",
          2863 => x"c00c87c0",
          2864 => x"9eb80883",
          2865 => x"f1c40c87",
          2866 => x"c09ebc08",
          2867 => x"83f1c80c",
          2868 => x"87c09ec0",
          2869 => x"0883f1cc",
          2870 => x"0c87c09e",
          2871 => x"c40883f1",
          2872 => x"d00c87c0",
          2873 => x"9e800852",
          2874 => x"7183f1d4",
          2875 => x"2387c09e",
          2876 => x"840883f1",
          2877 => x"d80c87c0",
          2878 => x"9e880883",
          2879 => x"f1dc0c87",
          2880 => x"c09e8c08",
          2881 => x"83f1e00c",
          2882 => x"810b83f1",
          2883 => x"e434800b",
          2884 => x"87c09e90",
          2885 => x"08708480",
          2886 => x"0a065152",
          2887 => x"527082fb",
          2888 => x"387183f1",
          2889 => x"e534800b",
          2890 => x"87c09e90",
          2891 => x"08708880",
          2892 => x"0a065152",
          2893 => x"5270802e",
          2894 => x"83388152",
          2895 => x"7183f1e6",
          2896 => x"34800b87",
          2897 => x"c09e9008",
          2898 => x"7090800a",
          2899 => x"06515252",
          2900 => x"70802e83",
          2901 => x"38815271",
          2902 => x"83f1e734",
          2903 => x"800b87c0",
          2904 => x"9e900870",
          2905 => x"88808006",
          2906 => x"51525270",
          2907 => x"802e8338",
          2908 => x"81527183",
          2909 => x"f1e83480",
          2910 => x"0b87c09e",
          2911 => x"900870a0",
          2912 => x"80800651",
          2913 => x"52527080",
          2914 => x"2e833881",
          2915 => x"527183f1",
          2916 => x"e934800b",
          2917 => x"87c09e90",
          2918 => x"08709080",
          2919 => x"80065152",
          2920 => x"5270802e",
          2921 => x"83388152",
          2922 => x"7183f1ea",
          2923 => x"34800b87",
          2924 => x"c09e9008",
          2925 => x"70848080",
          2926 => x"06515252",
          2927 => x"70802e83",
          2928 => x"38815271",
          2929 => x"83f1eb34",
          2930 => x"800b87c0",
          2931 => x"9e900870",
          2932 => x"82808006",
          2933 => x"51525270",
          2934 => x"802e8338",
          2935 => x"81527183",
          2936 => x"f1ec3480",
          2937 => x"0b87c09e",
          2938 => x"90087081",
          2939 => x"80800651",
          2940 => x"52527080",
          2941 => x"2e833881",
          2942 => x"527183f1",
          2943 => x"ed34800b",
          2944 => x"87c09e90",
          2945 => x"087080c0",
          2946 => x"80065152",
          2947 => x"5270802e",
          2948 => x"83388152",
          2949 => x"7183f1ee",
          2950 => x"34800b87",
          2951 => x"c09e9008",
          2952 => x"70a08006",
          2953 => x"51525270",
          2954 => x"802e8338",
          2955 => x"81527183",
          2956 => x"f1ef3487",
          2957 => x"c09e9008",
          2958 => x"98800670",
          2959 => x"8a2a5351",
          2960 => x"7183f1f0",
          2961 => x"34800b87",
          2962 => x"c09e9008",
          2963 => x"70848006",
          2964 => x"51525270",
          2965 => x"802e8338",
          2966 => x"81527183",
          2967 => x"f1f13487",
          2968 => x"c09e9008",
          2969 => x"83f00670",
          2970 => x"842a5351",
          2971 => x"7183f1f2",
          2972 => x"34800b87",
          2973 => x"c09e9008",
          2974 => x"70880651",
          2975 => x"52527080",
          2976 => x"2e833881",
          2977 => x"527183f1",
          2978 => x"f33487c0",
          2979 => x"9e900887",
          2980 => x"06517083",
          2981 => x"f1f43483",
          2982 => x"3d0d0481",
          2983 => x"52fd8239",
          2984 => x"fb3d0d83",
          2985 => x"d8a051ff",
          2986 => x"b6de3f83",
          2987 => x"f1e43354",
          2988 => x"7386aa38",
          2989 => x"83d8b451",
          2990 => x"c3b93f83",
          2991 => x"f1e63355",
          2992 => x"7485fa38",
          2993 => x"83f1eb33",
          2994 => x"547385d1",
          2995 => x"3883f1e8",
          2996 => x"33567585",
          2997 => x"a83883f1",
          2998 => x"e9335574",
          2999 => x"84ff3883",
          3000 => x"f1ea3354",
          3001 => x"7384d638",
          3002 => x"83f1ef33",
          3003 => x"567584b3",
          3004 => x"3883f1f3",
          3005 => x"33547384",
          3006 => x"903883f1",
          3007 => x"f1335574",
          3008 => x"83ed3883",
          3009 => x"f1e53356",
          3010 => x"7583cf38",
          3011 => x"83f1e733",
          3012 => x"547383b1",
          3013 => x"3883f1ec",
          3014 => x"33557483",
          3015 => x"933883f1",
          3016 => x"ed335675",
          3017 => x"82f43883",
          3018 => x"f1ee3354",
          3019 => x"7381ec38",
          3020 => x"83d8cc51",
          3021 => x"c2bd3f83",
          3022 => x"f1c80852",
          3023 => x"83d8d851",
          3024 => x"ffb5c53f",
          3025 => x"83f1cc08",
          3026 => x"5283d980",
          3027 => x"51ffb5b8",
          3028 => x"3f83f1d0",
          3029 => x"085283d9",
          3030 => x"a851ffb5",
          3031 => x"ab3f83d9",
          3032 => x"d051c28f",
          3033 => x"3f83f1d4",
          3034 => x"225283d9",
          3035 => x"d851ffb5",
          3036 => x"973f83f1",
          3037 => x"d80856bd",
          3038 => x"84c05275",
          3039 => x"51caa63f",
          3040 => x"84b8e408",
          3041 => x"bd84c029",
          3042 => x"76713154",
          3043 => x"5484b8e4",
          3044 => x"085283da",
          3045 => x"8051ffb4",
          3046 => x"ef3f83f1",
          3047 => x"eb335574",
          3048 => x"80c33883",
          3049 => x"f1e63355",
          3050 => x"748a388a",
          3051 => x"51c3af3f",
          3052 => x"873d0d04",
          3053 => x"83f1e008",
          3054 => x"56bd84c0",
          3055 => x"527551c9",
          3056 => x"e43f84b8",
          3057 => x"e408bd84",
          3058 => x"c0297671",
          3059 => x"31545484",
          3060 => x"b8e40852",
          3061 => x"83daac51",
          3062 => x"ffb4ad3f",
          3063 => x"8a51c2fe",
          3064 => x"3f873d0d",
          3065 => x"0483f1dc",
          3066 => x"0856bd84",
          3067 => x"c0527551",
          3068 => x"c9b33f84",
          3069 => x"b8e408bd",
          3070 => x"84c02976",
          3071 => x"71315454",
          3072 => x"84b8e408",
          3073 => x"5283dad8",
          3074 => x"51ffb3fc",
          3075 => x"3f83f1e6",
          3076 => x"33557480",
          3077 => x"2eff9438",
          3078 => x"ff9a3983",
          3079 => x"db8451c0",
          3080 => x"d23f83d8",
          3081 => x"cc51c0cb",
          3082 => x"3f83f1c8",
          3083 => x"085283d8",
          3084 => x"d851ffb3",
          3085 => x"d33f83f1",
          3086 => x"cc085283",
          3087 => x"d98051ff",
          3088 => x"b3c63f83",
          3089 => x"f1d00852",
          3090 => x"83d9a851",
          3091 => x"ffb3b93f",
          3092 => x"83d9d051",
          3093 => x"c09d3f83",
          3094 => x"f1d42252",
          3095 => x"83d9d851",
          3096 => x"ffb3a53f",
          3097 => x"83f1d808",
          3098 => x"56bd84c0",
          3099 => x"527551c8",
          3100 => x"b43f84b8",
          3101 => x"e408bd84",
          3102 => x"c0297671",
          3103 => x"31545484",
          3104 => x"b8e40852",
          3105 => x"83da8051",
          3106 => x"ffb2fd3f",
          3107 => x"83f1eb33",
          3108 => x"5574802e",
          3109 => x"fe8d38fe",
          3110 => x"cc3983db",
          3111 => x"8c51ffbf",
          3112 => x"d23f83f1",
          3113 => x"ee335473",
          3114 => x"802efd84",
          3115 => x"38feec39",
          3116 => x"83db9451",
          3117 => x"ffbfbc3f",
          3118 => x"83f1ed33",
          3119 => x"5675802e",
          3120 => x"fce538d6",
          3121 => x"3983dba0",
          3122 => x"51ffbfa7",
          3123 => x"3f83f1ec",
          3124 => x"33557480",
          3125 => x"2efcc738",
          3126 => x"d73983db",
          3127 => x"ac51ffbf",
          3128 => x"923f83f1",
          3129 => x"e7335473",
          3130 => x"802efca9",
          3131 => x"38d73983",
          3132 => x"f1f23352",
          3133 => x"83dbc051",
          3134 => x"ffb28d3f",
          3135 => x"83f1e533",
          3136 => x"5675802e",
          3137 => x"fc8638d2",
          3138 => x"3983f1f4",
          3139 => x"335283db",
          3140 => x"e051ffb1",
          3141 => x"f33f83f1",
          3142 => x"f1335574",
          3143 => x"802efbe3",
          3144 => x"38cd3983",
          3145 => x"f1f03352",
          3146 => x"83dc8051",
          3147 => x"ffb1d93f",
          3148 => x"83f1f333",
          3149 => x"5473802e",
          3150 => x"fbc038cd",
          3151 => x"3983f1b0",
          3152 => x"0883f1b4",
          3153 => x"08115452",
          3154 => x"83dca051",
          3155 => x"ffb1b93f",
          3156 => x"83f1ef33",
          3157 => x"5675802e",
          3158 => x"fb9738c7",
          3159 => x"3983f1a8",
          3160 => x"0883f1ac",
          3161 => x"08115452",
          3162 => x"83dcbc51",
          3163 => x"ffb1993f",
          3164 => x"83f1ea33",
          3165 => x"5473802e",
          3166 => x"faee38c1",
          3167 => x"3983f1a0",
          3168 => x"0883f1a4",
          3169 => x"08115452",
          3170 => x"83dcd851",
          3171 => x"ffb0f93f",
          3172 => x"83f1e933",
          3173 => x"5574802e",
          3174 => x"fac538c1",
          3175 => x"3983f1b8",
          3176 => x"0883f1bc",
          3177 => x"08115452",
          3178 => x"83dcf451",
          3179 => x"ffb0d93f",
          3180 => x"83f1e833",
          3181 => x"5675802e",
          3182 => x"fa9c38c1",
          3183 => x"3983f1c0",
          3184 => x"0883f1c4",
          3185 => x"08115452",
          3186 => x"83dd9051",
          3187 => x"ffb0b93f",
          3188 => x"83f1eb33",
          3189 => x"5473802e",
          3190 => x"f9f338c1",
          3191 => x"3983ddac",
          3192 => x"51ffb0a4",
          3193 => x"3f83d8b4",
          3194 => x"51ffbd87",
          3195 => x"3f83f1e6",
          3196 => x"33557480",
          3197 => x"2ef9cd38",
          3198 => x"c439ff3d",
          3199 => x"0d028e05",
          3200 => x"33527185",
          3201 => x"268c3871",
          3202 => x"101083c2",
          3203 => x"ec055271",
          3204 => x"080483dd",
          3205 => x"c051ffaf",
          3206 => x"ef3f833d",
          3207 => x"0d0483dd",
          3208 => x"c851ffaf",
          3209 => x"e33f833d",
          3210 => x"0d0483dd",
          3211 => x"d051ffaf",
          3212 => x"d73f833d",
          3213 => x"0d0483dd",
          3214 => x"d851ffaf",
          3215 => x"cb3f833d",
          3216 => x"0d0483dd",
          3217 => x"e051ffaf",
          3218 => x"bf3f833d",
          3219 => x"0d0483dd",
          3220 => x"e851ffaf",
          3221 => x"b33f833d",
          3222 => x"0d047188",
          3223 => x"800c0480",
          3224 => x"0b87c096",
          3225 => x"840c0483",
          3226 => x"f1f80887",
          3227 => x"c096840c",
          3228 => x"04d93d0d",
          3229 => x"aa3d08ad",
          3230 => x"3d085a5a",
          3231 => x"81705758",
          3232 => x"805283f2",
          3233 => x"d0085182",
          3234 => x"88823f84",
          3235 => x"b8e40880",
          3236 => x"ed388b3d",
          3237 => x"57ff0b83",
          3238 => x"f2d00854",
          3239 => x"5580f852",
          3240 => x"765182d2",
          3241 => x"8f3f84b8",
          3242 => x"e408802e",
          3243 => x"a4387651",
          3244 => x"c0f63f84",
          3245 => x"b8e40881",
          3246 => x"17575580",
          3247 => x"0b84b8e4",
          3248 => x"08258e38",
          3249 => x"84b8e408",
          3250 => x"ff057018",
          3251 => x"55558074",
          3252 => x"34740970",
          3253 => x"30707207",
          3254 => x"9f2a5155",
          3255 => x"5578762e",
          3256 => x"853873ff",
          3257 => x"b03883f2",
          3258 => x"d0088c11",
          3259 => x"08535182",
          3260 => x"879a3f84",
          3261 => x"b8e4088f",
          3262 => x"3878762e",
          3263 => x"9a387784",
          3264 => x"b8e40ca9",
          3265 => x"3d0d0483",
          3266 => x"e19851ff",
          3267 => x"adfa3f78",
          3268 => x"762e0981",
          3269 => x"06e83876",
          3270 => x"527951c0",
          3271 => x"aa3f7951",
          3272 => x"c0863fab",
          3273 => x"3d085684",
          3274 => x"b8e40876",
          3275 => x"34765283",
          3276 => x"e1c451ff",
          3277 => x"add23f80",
          3278 => x"0b84b8e4",
          3279 => x"0ca93d0d",
          3280 => x"04d83d0d",
          3281 => x"ab3d08ad",
          3282 => x"3d087172",
          3283 => x"5d723357",
          3284 => x"575a5773",
          3285 => x"a02e8191",
          3286 => x"38800b8d",
          3287 => x"3d595675",
          3288 => x"10101083",
          3289 => x"f2d80570",
          3290 => x"085254ff",
          3291 => x"bfba3f84",
          3292 => x"b8e40853",
          3293 => x"79527308",
          3294 => x"51c09a3f",
          3295 => x"84b8e408",
          3296 => x"90388414",
          3297 => x"33547381",
          3298 => x"2e818838",
          3299 => x"73822e99",
          3300 => x"38811670",
          3301 => x"81ff0657",
          3302 => x"54827627",
          3303 => x"c2388054",
          3304 => x"7384b8e4",
          3305 => x"0caa3d0d",
          3306 => x"04811a5a",
          3307 => x"aa3dff84",
          3308 => x"1153ff80",
          3309 => x"0551c7ce",
          3310 => x"3f84b8e4",
          3311 => x"08802ed1",
          3312 => x"38ff1b53",
          3313 => x"78527651",
          3314 => x"fda73f84",
          3315 => x"b8e40881",
          3316 => x"ff065473",
          3317 => x"802ec938",
          3318 => x"81167081",
          3319 => x"ff065754",
          3320 => x"827627fe",
          3321 => x"fa38ffb6",
          3322 => x"39783377",
          3323 => x"05567676",
          3324 => x"27fee638",
          3325 => x"8115705b",
          3326 => x"70335555",
          3327 => x"73a02e09",
          3328 => x"8106fed5",
          3329 => x"38757526",
          3330 => x"eb38800b",
          3331 => x"8d3d5956",
          3332 => x"fecd3973",
          3333 => x"84b8e408",
          3334 => x"5383f2d0",
          3335 => x"08525682",
          3336 => x"84ea3f84",
          3337 => x"b8e40880",
          3338 => x"d03883f2",
          3339 => x"d0085380",
          3340 => x"f8527751",
          3341 => x"82cefd3f",
          3342 => x"84b8e408",
          3343 => x"802eba38",
          3344 => x"7751ffbd",
          3345 => x"e33f84b8",
          3346 => x"e4085580",
          3347 => x"0b84b8e4",
          3348 => x"08259d38",
          3349 => x"84b8e408",
          3350 => x"ff057019",
          3351 => x"58558077",
          3352 => x"34775375",
          3353 => x"52811683",
          3354 => x"e18c5256",
          3355 => x"ffab993f",
          3356 => x"74ff2e09",
          3357 => x"8106ffb2",
          3358 => x"38810b84",
          3359 => x"b8e40caa",
          3360 => x"3d0d04ce",
          3361 => x"3d0db53d",
          3362 => x"08b73d08",
          3363 => x"b93d085a",
          3364 => x"415c800b",
          3365 => x"b43d3483",
          3366 => x"f2d43383",
          3367 => x"f2d00856",
          3368 => x"5d749e38",
          3369 => x"7483f2cc",
          3370 => x"33565674",
          3371 => x"802e82cb",
          3372 => x"3877802e",
          3373 => x"918d3881",
          3374 => x"7077065a",
          3375 => x"577890a0",
          3376 => x"3877802e",
          3377 => x"90fd3893",
          3378 => x"3db43d5f",
          3379 => x"5f8051eb",
          3380 => x"803f84b8",
          3381 => x"e408982b",
          3382 => x"70982c5b",
          3383 => x"5679ff2e",
          3384 => x"ec387981",
          3385 => x"ff0684d0",
          3386 => x"a0337098",
          3387 => x"2b70982c",
          3388 => x"84d09c33",
          3389 => x"70982b70",
          3390 => x"972c7198",
          3391 => x"2c057010",
          3392 => x"1083ddec",
          3393 => x"05700815",
          3394 => x"70335253",
          3395 => x"5c5d4652",
          3396 => x"5b585c59",
          3397 => x"81577479",
          3398 => x"2e80cd38",
          3399 => x"78752781",
          3400 => x"87387581",
          3401 => x"800a2981",
          3402 => x"ff0a0570",
          3403 => x"982c5755",
          3404 => x"80762481",
          3405 => x"cb387510",
          3406 => x"1670822b",
          3407 => x"5657800b",
          3408 => x"83ddf016",
          3409 => x"33425777",
          3410 => x"61259138",
          3411 => x"83ddec15",
          3412 => x"08187033",
          3413 => x"56417875",
          3414 => x"2e819538",
          3415 => x"76802ec2",
          3416 => x"387584d0",
          3417 => x"9c348157",
          3418 => x"76802e81",
          3419 => x"9938811b",
          3420 => x"70982b70",
          3421 => x"982c84d0",
          3422 => x"9c337098",
          3423 => x"2b70972c",
          3424 => x"71982c05",
          3425 => x"70822b83",
          3426 => x"ddf01133",
          3427 => x"5f535f5d",
          3428 => x"585d5757",
          3429 => x"7a782e81",
          3430 => x"90387684",
          3431 => x"d0a034fe",
          3432 => x"ac398157",
          3433 => x"76ffba38",
          3434 => x"7581800a",
          3435 => x"2981800a",
          3436 => x"0570982c",
          3437 => x"7081ff06",
          3438 => x"59574176",
          3439 => x"952680c0",
          3440 => x"38751016",
          3441 => x"70822b51",
          3442 => x"55800b83",
          3443 => x"ddf01633",
          3444 => x"42577761",
          3445 => x"25ce3883",
          3446 => x"ddec1508",
          3447 => x"18703342",
          3448 => x"5578612e",
          3449 => x"ffbc3876",
          3450 => x"802effbc",
          3451 => x"38fef239",
          3452 => x"81577680",
          3453 => x"2efeab38",
          3454 => x"fee73981",
          3455 => x"56fdb239",
          3456 => x"805776fe",
          3457 => x"e9387684",
          3458 => x"d0a03476",
          3459 => x"84d09c34",
          3460 => x"797e3476",
          3461 => x"7f0c6255",
          3462 => x"749526fd",
          3463 => x"b0387410",
          3464 => x"1083c384",
          3465 => x"05577608",
          3466 => x"0483ddf4",
          3467 => x"15087f0c",
          3468 => x"800b84d0",
          3469 => x"a034800b",
          3470 => x"84d09c34",
          3471 => x"d93984d0",
          3472 => x"a8335675",
          3473 => x"802efd85",
          3474 => x"3884d4c8",
          3475 => x"08528851",
          3476 => x"ffb69b3f",
          3477 => x"84d0a833",
          3478 => x"ff055776",
          3479 => x"84d0a834",
          3480 => x"fceb3984",
          3481 => x"d0a83370",
          3482 => x"81ff0684",
          3483 => x"d0a4335b",
          3484 => x"57557579",
          3485 => x"27fcd638",
          3486 => x"84d4c808",
          3487 => x"52811558",
          3488 => x"7784d0a8",
          3489 => x"347b1670",
          3490 => x"335255ff",
          3491 => x"b5e03ffc",
          3492 => x"bc397c93",
          3493 => x"2e8bda38",
          3494 => x"7c101083",
          3495 => x"f2800570",
          3496 => x"08575975",
          3497 => x"8f833875",
          3498 => x"84d0a434",
          3499 => x"757c3484",
          3500 => x"d0a43384",
          3501 => x"d0a83356",
          3502 => x"5674802e",
          3503 => x"b63884d4",
          3504 => x"c8085288",
          3505 => x"51ffb5a6",
          3506 => x"3f84d4c8",
          3507 => x"0852a051",
          3508 => x"ffb59b3f",
          3509 => x"84d4c808",
          3510 => x"528851ff",
          3511 => x"b5903f84",
          3512 => x"d0a833ff",
          3513 => x"055b7a84",
          3514 => x"d0a8347a",
          3515 => x"81ff0655",
          3516 => x"74cc387b",
          3517 => x"51ffa690",
          3518 => x"3f7584d0",
          3519 => x"a834fbcd",
          3520 => x"397c8a38",
          3521 => x"83f2c808",
          3522 => x"56758d9e",
          3523 => x"387c1010",
          3524 => x"83f1fc05",
          3525 => x"fc110857",
          3526 => x"55758ef9",
          3527 => x"38740856",
          3528 => x"75802efb",
          3529 => x"a8387551",
          3530 => x"ffb7fd3f",
          3531 => x"84b8e408",
          3532 => x"84d0a434",
          3533 => x"84b8e408",
          3534 => x"81ff0681",
          3535 => x"05537552",
          3536 => x"7b51ffb8",
          3537 => x"a53f84d0",
          3538 => x"a43384d0",
          3539 => x"a8335656",
          3540 => x"74802eff",
          3541 => x"9e3884d4",
          3542 => x"c8085288",
          3543 => x"51ffb48e",
          3544 => x"3f84d4c8",
          3545 => x"0852a051",
          3546 => x"ffb4833f",
          3547 => x"84d4c808",
          3548 => x"528851ff",
          3549 => x"b3f83f84",
          3550 => x"d0a833ff",
          3551 => x"05557484",
          3552 => x"d0a83474",
          3553 => x"81ff0655",
          3554 => x"c73984d0",
          3555 => x"a8337081",
          3556 => x"ff0684d0",
          3557 => x"a4335b57",
          3558 => x"55757927",
          3559 => x"faaf3884",
          3560 => x"d4c80852",
          3561 => x"81155776",
          3562 => x"84d0a834",
          3563 => x"7b167033",
          3564 => x"5255ffb3",
          3565 => x"b93f84d0",
          3566 => x"a8337081",
          3567 => x"ff0684d0",
          3568 => x"a4335a57",
          3569 => x"55757827",
          3570 => x"fa833884",
          3571 => x"d4c80852",
          3572 => x"81155776",
          3573 => x"84d0a834",
          3574 => x"7b167033",
          3575 => x"5255ffb3",
          3576 => x"8d3f84d0",
          3577 => x"a8337081",
          3578 => x"ff0684d0",
          3579 => x"a4335a57",
          3580 => x"55777626",
          3581 => x"ffa938f9",
          3582 => x"d43984d0",
          3583 => x"a83384d0",
          3584 => x"a4335656",
          3585 => x"74762ef9",
          3586 => x"c438ff15",
          3587 => x"5b7a84d0",
          3588 => x"a4347598",
          3589 => x"2b70982c",
          3590 => x"7c81ff06",
          3591 => x"43575a60",
          3592 => x"762480ef",
          3593 => x"3884d4c8",
          3594 => x"0852a051",
          3595 => x"ffb2bf3f",
          3596 => x"84d0a833",
          3597 => x"70982b70",
          3598 => x"982c84d0",
          3599 => x"a4335a57",
          3600 => x"57417477",
          3601 => x"24f98638",
          3602 => x"84d4c808",
          3603 => x"528851ff",
          3604 => x"b29c3f74",
          3605 => x"81800a29",
          3606 => x"81800a05",
          3607 => x"70982c84",
          3608 => x"d0a4335d",
          3609 => x"565a747b",
          3610 => x"24f8e238",
          3611 => x"84d4c808",
          3612 => x"528851ff",
          3613 => x"b1f83f74",
          3614 => x"81800a29",
          3615 => x"81800a05",
          3616 => x"70982c84",
          3617 => x"d0a4335d",
          3618 => x"565a7a75",
          3619 => x"25ffb938",
          3620 => x"f8bb397b",
          3621 => x"16588118",
          3622 => x"33783484",
          3623 => x"d4c80852",
          3624 => x"773351ff",
          3625 => x"b1c83f75",
          3626 => x"81800a29",
          3627 => x"81800a05",
          3628 => x"70982c84",
          3629 => x"d0a4335b",
          3630 => x"57557579",
          3631 => x"25fee638",
          3632 => x"7b165881",
          3633 => x"18337834",
          3634 => x"84d4c808",
          3635 => x"52773351",
          3636 => x"ffb19b3f",
          3637 => x"7581800a",
          3638 => x"2981800a",
          3639 => x"0570982c",
          3640 => x"84d0a433",
          3641 => x"5b575578",
          3642 => x"7624ffa7",
          3643 => x"38feb639",
          3644 => x"84d0a833",
          3645 => x"5574802e",
          3646 => x"f7d33884",
          3647 => x"d4c80852",
          3648 => x"8851ffb0",
          3649 => x"e93f84d0",
          3650 => x"a833ff05",
          3651 => x"577684d0",
          3652 => x"a8347681",
          3653 => x"ff0655dd",
          3654 => x"3984d0a4",
          3655 => x"337c055f",
          3656 => x"807f3484",
          3657 => x"d4c80852",
          3658 => x"8a51ffb0",
          3659 => x"c13f84d0",
          3660 => x"a4527b51",
          3661 => x"f48b3f84",
          3662 => x"b8e40881",
          3663 => x"ff065877",
          3664 => x"89cf3884",
          3665 => x"d0a43357",
          3666 => x"76802e80",
          3667 => x"d83883f2",
          3668 => x"d4337010",
          3669 => x"1083f1fc",
          3670 => x"05700857",
          3671 => x"5e56748b",
          3672 => x"a0387582",
          3673 => x"2b87fc06",
          3674 => x"83f1fc05",
          3675 => x"81187053",
          3676 => x"575b80e7",
          3677 => x"fb3f84b8",
          3678 => x"e4087b0c",
          3679 => x"83f2d433",
          3680 => x"70101083",
          3681 => x"f1fc0570",
          3682 => x"08574141",
          3683 => x"748bad38",
          3684 => x"83f2d008",
          3685 => x"5675802e",
          3686 => x"8c3883f2",
          3687 => x"cc335877",
          3688 => x"802e8bbc",
          3689 => x"38800b84",
          3690 => x"d0a83480",
          3691 => x"0b84d0a4",
          3692 => x"347b84b8",
          3693 => x"e40cb43d",
          3694 => x"0d0484d0",
          3695 => x"a8335574",
          3696 => x"802eb638",
          3697 => x"84d4c808",
          3698 => x"528851ff",
          3699 => x"afa03f84",
          3700 => x"d4c80852",
          3701 => x"a051ffaf",
          3702 => x"953f84d4",
          3703 => x"c8085288",
          3704 => x"51ffaf8a",
          3705 => x"3f84d0a8",
          3706 => x"33ff0556",
          3707 => x"7584d0a8",
          3708 => x"347581ff",
          3709 => x"065574cc",
          3710 => x"3883d1e0",
          3711 => x"51ffa088",
          3712 => x"3f800b84",
          3713 => x"d0a83480",
          3714 => x"0b84d0a4",
          3715 => x"34f5be39",
          3716 => x"837c3480",
          3717 => x"0b811d34",
          3718 => x"84d0a833",
          3719 => x"5574802e",
          3720 => x"b63884d4",
          3721 => x"c8085288",
          3722 => x"51ffaec2",
          3723 => x"3f84d4c8",
          3724 => x"0852a051",
          3725 => x"ffaeb73f",
          3726 => x"84d4c808",
          3727 => x"528851ff",
          3728 => x"aeac3f84",
          3729 => x"d0a833ff",
          3730 => x"055d7c84",
          3731 => x"d0a8347c",
          3732 => x"81ff0655",
          3733 => x"74cc3883",
          3734 => x"d1e051ff",
          3735 => x"9faa3f80",
          3736 => x"0b84d0a8",
          3737 => x"34800b84",
          3738 => x"d0a4347b",
          3739 => x"84b8e40c",
          3740 => x"b43d0d04",
          3741 => x"84d0a833",
          3742 => x"7081ff06",
          3743 => x"5c567a80",
          3744 => x"2ef4ca38",
          3745 => x"84d0a433",
          3746 => x"ff055978",
          3747 => x"84d0a434",
          3748 => x"ff165877",
          3749 => x"84d0a834",
          3750 => x"84d4c808",
          3751 => x"528851ff",
          3752 => x"adcc3f84",
          3753 => x"d0a83370",
          3754 => x"982b7098",
          3755 => x"2c84d0a4",
          3756 => x"335a525b",
          3757 => x"56767624",
          3758 => x"80ef3884",
          3759 => x"d4c80852",
          3760 => x"a051ffad",
          3761 => x"a93f84d0",
          3762 => x"a8337098",
          3763 => x"2b70982c",
          3764 => x"84d0a433",
          3765 => x"5d575956",
          3766 => x"747a24f3",
          3767 => x"f03884d4",
          3768 => x"c8085288",
          3769 => x"51ffad86",
          3770 => x"3f748180",
          3771 => x"0a298180",
          3772 => x"0a057098",
          3773 => x"2c84d0a4",
          3774 => x"335b5155",
          3775 => x"747924f3",
          3776 => x"cc3884d4",
          3777 => x"c8085288",
          3778 => x"51fface2",
          3779 => x"3f748180",
          3780 => x"0a298180",
          3781 => x"0a057098",
          3782 => x"2c84d0a4",
          3783 => x"335b5155",
          3784 => x"787525ff",
          3785 => x"b938f3a5",
          3786 => x"397b1657",
          3787 => x"81173377",
          3788 => x"3484d4c8",
          3789 => x"08527633",
          3790 => x"51ffacb2",
          3791 => x"3f758180",
          3792 => x"0a298180",
          3793 => x"0a057098",
          3794 => x"2c84d0a4",
          3795 => x"3343575b",
          3796 => x"756125fe",
          3797 => x"e6387b16",
          3798 => x"57811733",
          3799 => x"773484d4",
          3800 => x"c8085276",
          3801 => x"3351ffac",
          3802 => x"853f7581",
          3803 => x"800a2981",
          3804 => x"800a0570",
          3805 => x"982c84d0",
          3806 => x"a4334357",
          3807 => x"5b607624",
          3808 => x"ffa738fe",
          3809 => x"b63984d0",
          3810 => x"a8337081",
          3811 => x"ff065858",
          3812 => x"76602ef2",
          3813 => x"b83884d0",
          3814 => x"a4335576",
          3815 => x"7527ae38",
          3816 => x"74982b70",
          3817 => x"982c5741",
          3818 => x"767624a1",
          3819 => x"387b165b",
          3820 => x"7a33811c",
          3821 => x"34758180",
          3822 => x"0a2981ff",
          3823 => x"0a057098",
          3824 => x"2c84d0a8",
          3825 => x"33525758",
          3826 => x"757825e1",
          3827 => x"38811855",
          3828 => x"7484d0a8",
          3829 => x"347781ff",
          3830 => x"067c055a",
          3831 => x"b33d337a",
          3832 => x"3484d0a4",
          3833 => x"33577660",
          3834 => x"258b3881",
          3835 => x"17567584",
          3836 => x"d0a43475",
          3837 => x"5784d0a8",
          3838 => x"33708180",
          3839 => x"0a2981ff",
          3840 => x"0a057098",
          3841 => x"2c7981ff",
          3842 => x"0644585c",
          3843 => x"58607624",
          3844 => x"81ef3877",
          3845 => x"982b7098",
          3846 => x"2c7881ff",
          3847 => x"065c5759",
          3848 => x"757a25f1",
          3849 => x"a83884d4",
          3850 => x"c8085288",
          3851 => x"51ffaabe",
          3852 => x"3f758180",
          3853 => x"0a298180",
          3854 => x"0a057098",
          3855 => x"2c84d0a4",
          3856 => x"33575741",
          3857 => x"757525f1",
          3858 => x"843884d4",
          3859 => x"c8085288",
          3860 => x"51ffaa9a",
          3861 => x"3f758180",
          3862 => x"0a298180",
          3863 => x"0a057098",
          3864 => x"2c84d0a4",
          3865 => x"33575741",
          3866 => x"747624ff",
          3867 => x"b938f0dd",
          3868 => x"3983f1fc",
          3869 => x"08567580",
          3870 => x"2ef49d38",
          3871 => x"7551ffad",
          3872 => x"a73f84b8",
          3873 => x"e40884d0",
          3874 => x"a43484b8",
          3875 => x"e40881ff",
          3876 => x"06810553",
          3877 => x"75527b51",
          3878 => x"ffadcf3f",
          3879 => x"84d0a433",
          3880 => x"84d0a833",
          3881 => x"56567480",
          3882 => x"2ef4c838",
          3883 => x"84d4c808",
          3884 => x"528851ff",
          3885 => x"a9b83f84",
          3886 => x"d4c80852",
          3887 => x"a051ffa9",
          3888 => x"ad3f84d4",
          3889 => x"c8085288",
          3890 => x"51ffa9a2",
          3891 => x"3f84d0a8",
          3892 => x"33ff055b",
          3893 => x"7a84d0a8",
          3894 => x"347a81ff",
          3895 => x"0655c739",
          3896 => x"a85180e1",
          3897 => x"8b3f84b8",
          3898 => x"e40883f2",
          3899 => x"d00c84b8",
          3900 => x"e40885a5",
          3901 => x"387683f2",
          3902 => x"cc3477ef",
          3903 => x"ca3880c3",
          3904 => x"3984d4c8",
          3905 => x"08527b16",
          3906 => x"70335258",
          3907 => x"ffa8df3f",
          3908 => x"7581800a",
          3909 => x"2981800a",
          3910 => x"0570982c",
          3911 => x"84d0a433",
          3912 => x"52575776",
          3913 => x"7624da38",
          3914 => x"84d0a833",
          3915 => x"70982b70",
          3916 => x"982c7981",
          3917 => x"ff065d58",
          3918 => x"5a58757a",
          3919 => x"25ef8e38",
          3920 => x"fde43983",
          3921 => x"f2d00880",
          3922 => x"2eeefc38",
          3923 => x"83f1fc57",
          3924 => x"93567608",
          3925 => x"5574bb38",
          3926 => x"ff168418",
          3927 => x"58567580",
          3928 => x"25f03880",
          3929 => x"0b83f2d4",
          3930 => x"3483f2d0",
          3931 => x"08557480",
          3932 => x"2eeed438",
          3933 => x"745181e7",
          3934 => x"f63f83f2",
          3935 => x"d0085180",
          3936 => x"d9fe3f80",
          3937 => x"0b83f2d0",
          3938 => x"0c933db4",
          3939 => x"3d5f5fee",
          3940 => x"bc397451",
          3941 => x"80d9e93f",
          3942 => x"80770cff",
          3943 => x"16841858",
          3944 => x"56758025",
          3945 => x"ffac38ff",
          3946 => x"ba397551",
          3947 => x"ffaaf93f",
          3948 => x"84b8e408",
          3949 => x"84d0a434",
          3950 => x"84b8e408",
          3951 => x"81ff0681",
          3952 => x"05537552",
          3953 => x"7b51ffab",
          3954 => x"a13f930b",
          3955 => x"84d0a433",
          3956 => x"84d0a833",
          3957 => x"57575d74",
          3958 => x"802ef297",
          3959 => x"3884d4c8",
          3960 => x"08528851",
          3961 => x"ffa7873f",
          3962 => x"84d4c808",
          3963 => x"52a051ff",
          3964 => x"a6fc3f84",
          3965 => x"d4c80852",
          3966 => x"8851ffa6",
          3967 => x"f13f84d0",
          3968 => x"a833ff05",
          3969 => x"5a7984d0",
          3970 => x"a8347981",
          3971 => x"ff0655c7",
          3972 => x"39807c34",
          3973 => x"800b84d0",
          3974 => x"a834800b",
          3975 => x"84d0a434",
          3976 => x"7b84b8e4",
          3977 => x"0cb43d0d",
          3978 => x"047551ff",
          3979 => x"a9fa3f84",
          3980 => x"b8e40884",
          3981 => x"d0a43484",
          3982 => x"b8e40881",
          3983 => x"ff068105",
          3984 => x"5375527b",
          3985 => x"51ffaaa2",
          3986 => x"3f811d70",
          3987 => x"81ff0684",
          3988 => x"d0a43384",
          3989 => x"d0a83358",
          3990 => x"525e5674",
          3991 => x"802ef193",
          3992 => x"3884d4c8",
          3993 => x"08528851",
          3994 => x"ffa6833f",
          3995 => x"84d4c808",
          3996 => x"52a051ff",
          3997 => x"a5f83f84",
          3998 => x"d4c80852",
          3999 => x"8851ffa5",
          4000 => x"ed3f84d0",
          4001 => x"a833ff05",
          4002 => x"577684d0",
          4003 => x"a8347681",
          4004 => x"ff0655c7",
          4005 => x"397551ff",
          4006 => x"a98e3f84",
          4007 => x"b8e40884",
          4008 => x"d0a43484",
          4009 => x"b8e40881",
          4010 => x"ff068105",
          4011 => x"5375527b",
          4012 => x"51ffa9b6",
          4013 => x"3fff1d70",
          4014 => x"81ff0684",
          4015 => x"d0a43384",
          4016 => x"d0a83358",
          4017 => x"585e5874",
          4018 => x"802ef0a7",
          4019 => x"3884d4c8",
          4020 => x"08528851",
          4021 => x"ffa5973f",
          4022 => x"84d4c808",
          4023 => x"52a051ff",
          4024 => x"a58c3f84",
          4025 => x"d4c80852",
          4026 => x"8851ffa5",
          4027 => x"813f84d0",
          4028 => x"a833ff05",
          4029 => x"416084d0",
          4030 => x"a8346081",
          4031 => x"ff0655c7",
          4032 => x"39745180",
          4033 => x"d6fa3f83",
          4034 => x"f2d43370",
          4035 => x"822b87fc",
          4036 => x"0683f1fc",
          4037 => x"05811970",
          4038 => x"54525c56",
          4039 => x"80dcd13f",
          4040 => x"84b8e408",
          4041 => x"7b0c83f2",
          4042 => x"d4337010",
          4043 => x"1083f1fc",
          4044 => x"05700857",
          4045 => x"41417480",
          4046 => x"2ef4d538",
          4047 => x"75537b52",
          4048 => x"7451ffa8",
          4049 => x"a53f83f2",
          4050 => x"d4338105",
          4051 => x"7081ff06",
          4052 => x"5a569379",
          4053 => x"2782f238",
          4054 => x"7783f2d4",
          4055 => x"34f4b139",
          4056 => x"b43dfef8",
          4057 => x"05547653",
          4058 => x"7b527551",
          4059 => x"81d8c03f",
          4060 => x"83f2d008",
          4061 => x"528a5182",
          4062 => x"ba883f83",
          4063 => x"f2d00851",
          4064 => x"81dff33f",
          4065 => x"800b84d0",
          4066 => x"a834800b",
          4067 => x"84d0a434",
          4068 => x"7b84b8e4",
          4069 => x"0cb43d0d",
          4070 => x"04935377",
          4071 => x"5284b8e4",
          4072 => x"085181c9",
          4073 => x"f83f84b8",
          4074 => x"e40882a5",
          4075 => x"3884b8e4",
          4076 => x"08963d5c",
          4077 => x"5d83f2d0",
          4078 => x"085380f8",
          4079 => x"527a5182",
          4080 => x"b7f23f84",
          4081 => x"b8e4085a",
          4082 => x"84b8e408",
          4083 => x"7b2e0981",
          4084 => x"06e9ee38",
          4085 => x"84b8e408",
          4086 => x"51ffa6cc",
          4087 => x"3f84b8e4",
          4088 => x"0856800b",
          4089 => x"84b8e408",
          4090 => x"2580e338",
          4091 => x"84b8e408",
          4092 => x"ff05701b",
          4093 => x"58568077",
          4094 => x"347581ff",
          4095 => x"0683f2d4",
          4096 => x"33701010",
          4097 => x"83f1fc05",
          4098 => x"70085840",
          4099 => x"58597480",
          4100 => x"f2387682",
          4101 => x"2b87fc06",
          4102 => x"83f1fc05",
          4103 => x"811a7053",
          4104 => x"585580da",
          4105 => x"cb3f84b8",
          4106 => x"e408750c",
          4107 => x"83f2d433",
          4108 => x"70101083",
          4109 => x"f1fc0570",
          4110 => x"08574041",
          4111 => x"74a03881",
          4112 => x"1d7081ff",
          4113 => x"065e5793",
          4114 => x"7d278338",
          4115 => x"805d75ff",
          4116 => x"2e098106",
          4117 => x"fedf3877",
          4118 => x"e8ed38f9",
          4119 => x"e6397653",
          4120 => x"79527451",
          4121 => x"ffa6833f",
          4122 => x"83f2d433",
          4123 => x"81057081",
          4124 => x"ff065b57",
          4125 => x"937a2780",
          4126 => x"c838800b",
          4127 => x"83f2d434",
          4128 => x"ffbd3974",
          4129 => x"5180d3f8",
          4130 => x"3f83f2d4",
          4131 => x"3370822b",
          4132 => x"87fc0683",
          4133 => x"f1fc0581",
          4134 => x"1b705452",
          4135 => x"565780d9",
          4136 => x"cf3f84b8",
          4137 => x"e408750c",
          4138 => x"83f2d433",
          4139 => x"70101083",
          4140 => x"f1fc0570",
          4141 => x"08574041",
          4142 => x"74802eff",
          4143 => x"8238ff9e",
          4144 => x"397683f2",
          4145 => x"d434fef7",
          4146 => x"397583f2",
          4147 => x"d434f1c0",
          4148 => x"3983e0cc",
          4149 => x"51ff9f9b",
          4150 => x"3f77e7eb",
          4151 => x"38f8e439",
          4152 => x"f23d0d02",
          4153 => x"80c30533",
          4154 => x"02840580",
          4155 => x"c705335b",
          4156 => x"53728326",
          4157 => x"818d3872",
          4158 => x"812e818b",
          4159 => x"38817325",
          4160 => x"839e3872",
          4161 => x"822e82a8",
          4162 => x"3886a7a0",
          4163 => x"805986a7",
          4164 => x"b080705e",
          4165 => x"5780569f",
          4166 => x"a0587976",
          4167 => x"2e903875",
          4168 => x"83f89434",
          4169 => x"7583f895",
          4170 => x"347583f8",
          4171 => x"922383f8",
          4172 => x"90337098",
          4173 => x"2b71902b",
          4174 => x"0771882b",
          4175 => x"0771077a",
          4176 => x"7f565656",
          4177 => x"5b787727",
          4178 => x"94388074",
          4179 => x"70840556",
          4180 => x"0c747370",
          4181 => x"8405550c",
          4182 => x"767426ee",
          4183 => x"38757827",
          4184 => x"a23883f8",
          4185 => x"90338497",
          4186 => x"b6177978",
          4187 => x"31555555",
          4188 => x"a00be0e0",
          4189 => x"15347474",
          4190 => x"70810556",
          4191 => x"34ff1353",
          4192 => x"72ee3890",
          4193 => x"3d0d0486",
          4194 => x"a7a0800b",
          4195 => x"83f89433",
          4196 => x"70101011",
          4197 => x"83f89533",
          4198 => x"71902911",
          4199 => x"74055b41",
          4200 => x"58405986",
          4201 => x"a7b0800b",
          4202 => x"84b6d833",
          4203 => x"7081ff06",
          4204 => x"84b6d733",
          4205 => x"7081ff06",
          4206 => x"83f89222",
          4207 => x"7083ffff",
          4208 => x"06707529",
          4209 => x"5d595d58",
          4210 => x"5e575b5d",
          4211 => x"73732687",
          4212 => x"38727431",
          4213 => x"75295679",
          4214 => x"81ff067e",
          4215 => x"81ff067c",
          4216 => x"81ff067a",
          4217 => x"83ffff06",
          4218 => x"6281ff06",
          4219 => x"70752914",
          4220 => x"5d425757",
          4221 => x"5b5c7474",
          4222 => x"268f3883",
          4223 => x"f8943374",
          4224 => x"76310570",
          4225 => x"7d291b59",
          4226 => x"5f768306",
          4227 => x"5c7b802e",
          4228 => x"fe9c3878",
          4229 => x"7d555372",
          4230 => x"7726fec1",
          4231 => x"38807370",
          4232 => x"81055534",
          4233 => x"83f89033",
          4234 => x"74708105",
          4235 => x"5634e839",
          4236 => x"86a7a080",
          4237 => x"5986a7b0",
          4238 => x"807084b6",
          4239 => x"d8337081",
          4240 => x"ff0684b6",
          4241 => x"d7337081",
          4242 => x"ff0683f8",
          4243 => x"92227074",
          4244 => x"295d5b5d",
          4245 => x"575e565e",
          4246 => x"57747827",
          4247 => x"81df3873",
          4248 => x"81ff0673",
          4249 => x"81ff0671",
          4250 => x"7129185a",
          4251 => x"54547980",
          4252 => x"2efdbb38",
          4253 => x"800b83f8",
          4254 => x"9434800b",
          4255 => x"83f89534",
          4256 => x"83f89033",
          4257 => x"70982b71",
          4258 => x"902b0771",
          4259 => x"882b0771",
          4260 => x"077a7f56",
          4261 => x"56565b76",
          4262 => x"7926fdae",
          4263 => x"38fdbe39",
          4264 => x"72fce638",
          4265 => x"83f89433",
          4266 => x"7081ff06",
          4267 => x"70101011",
          4268 => x"83f89533",
          4269 => x"71902911",
          4270 => x"86a7a080",
          4271 => x"115e575b",
          4272 => x"56565f86",
          4273 => x"a7b08070",
          4274 => x"1484b6d8",
          4275 => x"337081ff",
          4276 => x"0684b6d7",
          4277 => x"337081ff",
          4278 => x"0683f892",
          4279 => x"227083ff",
          4280 => x"ff067c75",
          4281 => x"2960055e",
          4282 => x"5a415f58",
          4283 => x"5f405e57",
          4284 => x"7973268b",
          4285 => x"38727a31",
          4286 => x"15707d29",
          4287 => x"1957537d",
          4288 => x"81ff0674",
          4289 => x"81ff0671",
          4290 => x"71297d83",
          4291 => x"ffff0662",
          4292 => x"81ff0670",
          4293 => x"7529585f",
          4294 => x"5b5c5d55",
          4295 => x"7b782685",
          4296 => x"38777529",
          4297 => x"53797331",
          4298 => x"16798306",
          4299 => x"5b5879fd",
          4300 => x"e2387683",
          4301 => x"065c7bfd",
          4302 => x"da38fbf2",
          4303 => x"39747831",
          4304 => x"7b2956fe",
          4305 => x"9a39fb3d",
          4306 => x"0d86ee80",
          4307 => x"8c53ff8a",
          4308 => x"73348773",
          4309 => x"34857334",
          4310 => x"81733486",
          4311 => x"ee809c55",
          4312 => x"80f47534",
          4313 => x"ffb07534",
          4314 => x"86ee8098",
          4315 => x"56807634",
          4316 => x"80763486",
          4317 => x"ee809454",
          4318 => x"8a743480",
          4319 => x"7434ff80",
          4320 => x"75348152",
          4321 => x"8351fad8",
          4322 => x"3f86a087",
          4323 => x"e0700854",
          4324 => x"5481f856",
          4325 => x"86a081f8",
          4326 => x"73770684",
          4327 => x"07545572",
          4328 => x"75347308",
          4329 => x"7080ff06",
          4330 => x"80c00751",
          4331 => x"53727534",
          4332 => x"86a087cc",
          4333 => x"08707706",
          4334 => x"81075153",
          4335 => x"7286a081",
          4336 => x"f3347308",
          4337 => x"81f70688",
          4338 => x"07537275",
          4339 => x"3480d00b",
          4340 => x"84b6d834",
          4341 => x"800b84b8",
          4342 => x"e40c873d",
          4343 => x"0d0484b6",
          4344 => x"d83384b8",
          4345 => x"e40c04f7",
          4346 => x"3d0d02af",
          4347 => x"05330284",
          4348 => x"05b30533",
          4349 => x"84b6d733",
          4350 => x"5b595681",
          4351 => x"53757926",
          4352 => x"82da3884",
          4353 => x"b6d83383",
          4354 => x"f8953383",
          4355 => x"f8943372",
          4356 => x"71291286",
          4357 => x"a7a08011",
          4358 => x"83f89222",
          4359 => x"5f515759",
          4360 => x"717c2905",
          4361 => x"7083ffff",
          4362 => x"0683f6ea",
          4363 => x"33535758",
          4364 => x"5372812e",
          4365 => x"83c43883",
          4366 => x"f8922276",
          4367 => x"05557483",
          4368 => x"f8922383",
          4369 => x"f8943376",
          4370 => x"057081ff",
          4371 => x"067a81ff",
          4372 => x"06555b55",
          4373 => x"727a2682",
          4374 => x"8c38ff19",
          4375 => x"537283f8",
          4376 => x"943483f8",
          4377 => x"92227083",
          4378 => x"ffff0684",
          4379 => x"b6d6335c",
          4380 => x"55577974",
          4381 => x"26828938",
          4382 => x"84b6d833",
          4383 => x"76712954",
          4384 => x"58805472",
          4385 => x"9f9f26ac",
          4386 => x"388497b6",
          4387 => x"70145455",
          4388 => x"e0e01333",
          4389 => x"e0e01634",
          4390 => x"72708105",
          4391 => x"54337570",
          4392 => x"81055734",
          4393 => x"81145484",
          4394 => x"b6d57327",
          4395 => x"e338739f",
          4396 => x"9f26a138",
          4397 => x"83f89033",
          4398 => x"8497b615",
          4399 => x"5455a00b",
          4400 => x"e0e01434",
          4401 => x"74737081",
          4402 => x"05553481",
          4403 => x"14549f9f",
          4404 => x"7427eb38",
          4405 => x"84b6d633",
          4406 => x"ff055675",
          4407 => x"83f89223",
          4408 => x"75577881",
          4409 => x"ff067783",
          4410 => x"ffff0654",
          4411 => x"54737326",
          4412 => x"81fd3872",
          4413 => x"74318105",
          4414 => x"84b6d833",
          4415 => x"71712958",
          4416 => x"55577555",
          4417 => x"86a7a080",
          4418 => x"5886a7b0",
          4419 => x"807981ff",
          4420 => x"067581ff",
          4421 => x"06717129",
          4422 => x"195c5c54",
          4423 => x"57757927",
          4424 => x"b9388497",
          4425 => x"b61654e0",
          4426 => x"e0143353",
          4427 => x"84b6e013",
          4428 => x"33787081",
          4429 => x"055a3473",
          4430 => x"70810555",
          4431 => x"33777081",
          4432 => x"05593481",
          4433 => x"1584b6d8",
          4434 => x"3384b6d7",
          4435 => x"33717129",
          4436 => x"19565c5a",
          4437 => x"55727526",
          4438 => x"ce388053",
          4439 => x"7284b8e4",
          4440 => x"0c8b3d0d",
          4441 => x"047483f8",
          4442 => x"943483f8",
          4443 => x"92227083",
          4444 => x"ffff0684",
          4445 => x"b6d6335c",
          4446 => x"5557737a",
          4447 => x"27fdf938",
          4448 => x"77802efe",
          4449 => x"dd387881",
          4450 => x"ff06ff05",
          4451 => x"83f89433",
          4452 => x"56537275",
          4453 => x"2e098106",
          4454 => x"fec83873",
          4455 => x"76318105",
          4456 => x"84b6d833",
          4457 => x"71712978",
          4458 => x"72291156",
          4459 => x"52595473",
          4460 => x"7327feae",
          4461 => x"3883f890",
          4462 => x"338497b6",
          4463 => x"15747631",
          4464 => x"555656a0",
          4465 => x"0be0e016",
          4466 => x"34757570",
          4467 => x"81055734",
          4468 => x"ff135372",
          4469 => x"802efe8a",
          4470 => x"38a00be0",
          4471 => x"e0163475",
          4472 => x"75708105",
          4473 => x"5734ff13",
          4474 => x"5372d838",
          4475 => x"fdf43980",
          4476 => x"0b84b6d8",
          4477 => x"335556fe",
          4478 => x"893983f8",
          4479 => x"96153359",
          4480 => x"84b6e019",
          4481 => x"33743484",
          4482 => x"b6d73359",
          4483 => x"fca939fc",
          4484 => x"3d0d7602",
          4485 => x"84059f05",
          4486 => x"33535170",
          4487 => x"86269b38",
          4488 => x"70101083",
          4489 => x"c3dc0551",
          4490 => x"70080484",
          4491 => x"b6d83351",
          4492 => x"71712786",
          4493 => x"387183f8",
          4494 => x"9534800b",
          4495 => x"84b8e40c",
          4496 => x"863d0d04",
          4497 => x"800b83f8",
          4498 => x"953483f8",
          4499 => x"94337081",
          4500 => x"ff065452",
          4501 => x"72802ee2",
          4502 => x"38ff1251",
          4503 => x"7083f894",
          4504 => x"34800b84",
          4505 => x"b8e40c86",
          4506 => x"3d0d0483",
          4507 => x"f8943370",
          4508 => x"73317009",
          4509 => x"709f2c72",
          4510 => x"06545553",
          4511 => x"547083f8",
          4512 => x"9434de39",
          4513 => x"83f89433",
          4514 => x"720584b6",
          4515 => x"d733ff11",
          4516 => x"55565170",
          4517 => x"75258338",
          4518 => x"70537283",
          4519 => x"f8943480",
          4520 => x"0b84b8e4",
          4521 => x"0c863d0d",
          4522 => x"0483f895",
          4523 => x"33707331",
          4524 => x"7009709f",
          4525 => x"2c720654",
          4526 => x"56535570",
          4527 => x"83f89534",
          4528 => x"800b84b8",
          4529 => x"e40c863d",
          4530 => x"0d0483f8",
          4531 => x"95337205",
          4532 => x"84b6d833",
          4533 => x"ff115555",
          4534 => x"51707425",
          4535 => x"83387053",
          4536 => x"7283f895",
          4537 => x"34800b84",
          4538 => x"b8e40c86",
          4539 => x"3d0d0480",
          4540 => x"0b83f895",
          4541 => x"3483f894",
          4542 => x"3384b6d7",
          4543 => x"33ff0556",
          4544 => x"52717525",
          4545 => x"feb43881",
          4546 => x"12517083",
          4547 => x"f89434fe",
          4548 => x"d039ff3d",
          4549 => x"0d028f05",
          4550 => x"335170b1",
          4551 => x"26b33870",
          4552 => x"101083c3",
          4553 => x"f8055170",
          4554 => x"080483f8",
          4555 => x"90337080",
          4556 => x"f0067184",
          4557 => x"2b80f006",
          4558 => x"7072842a",
          4559 => x"07515253",
          4560 => x"517180f0",
          4561 => x"2e098106",
          4562 => x"9c3880f2",
          4563 => x"0b83f890",
          4564 => x"34800b84",
          4565 => x"b8e40c83",
          4566 => x"3d0d0483",
          4567 => x"f8903381",
          4568 => x"9f069007",
          4569 => x"517083f8",
          4570 => x"9034800b",
          4571 => x"84b8e40c",
          4572 => x"833d0d04",
          4573 => x"83f89033",
          4574 => x"80f00751",
          4575 => x"7083f890",
          4576 => x"34e83983",
          4577 => x"f8903381",
          4578 => x"fe068607",
          4579 => x"517083f8",
          4580 => x"9034d739",
          4581 => x"80f10b83",
          4582 => x"f8903480",
          4583 => x"0b84b8e4",
          4584 => x"0c833d0d",
          4585 => x"0483f890",
          4586 => x"3381fc06",
          4587 => x"84075170",
          4588 => x"83f89034",
          4589 => x"ffb43983",
          4590 => x"f8903387",
          4591 => x"07517083",
          4592 => x"f89034ff",
          4593 => x"a53983f8",
          4594 => x"903381fd",
          4595 => x"06850751",
          4596 => x"7083f890",
          4597 => x"34ff9339",
          4598 => x"83f89033",
          4599 => x"81fb0683",
          4600 => x"07517083",
          4601 => x"f89034ff",
          4602 => x"813983f8",
          4603 => x"903381f9",
          4604 => x"06810751",
          4605 => x"7083f890",
          4606 => x"34feef39",
          4607 => x"83f89033",
          4608 => x"81f80651",
          4609 => x"7083f890",
          4610 => x"34fedf39",
          4611 => x"83f89033",
          4612 => x"81df0680",
          4613 => x"d0075170",
          4614 => x"83f89034",
          4615 => x"fecc3983",
          4616 => x"f8903381",
          4617 => x"bf06b007",
          4618 => x"517083f8",
          4619 => x"9034feba",
          4620 => x"3983f890",
          4621 => x"3381ef06",
          4622 => x"80e00751",
          4623 => x"7083f890",
          4624 => x"34fea739",
          4625 => x"83f89033",
          4626 => x"81cf0680",
          4627 => x"c0075170",
          4628 => x"83f89034",
          4629 => x"fe943983",
          4630 => x"f8903381",
          4631 => x"af06a007",
          4632 => x"517083f8",
          4633 => x"9034fe82",
          4634 => x"3983f890",
          4635 => x"33818f06",
          4636 => x"517083f8",
          4637 => x"9034fdf2",
          4638 => x"3983f890",
          4639 => x"3381fa06",
          4640 => x"82075170",
          4641 => x"83f89034",
          4642 => x"fde039f3",
          4643 => x"3d0d02bf",
          4644 => x"05330284",
          4645 => x"0580c305",
          4646 => x"3383f894",
          4647 => x"3383f893",
          4648 => x"3383f895",
          4649 => x"3384b6da",
          4650 => x"3343415f",
          4651 => x"5d5b5978",
          4652 => x"822e82a1",
          4653 => x"38788224",
          4654 => x"a5387881",
          4655 => x"2e818238",
          4656 => x"7d84b6da",
          4657 => x"34800b84",
          4658 => x"b6dc347a",
          4659 => x"83f89434",
          4660 => x"7b83f892",
          4661 => x"237c83f8",
          4662 => x"95348f3d",
          4663 => x"0d047883",
          4664 => x"2e098106",
          4665 => x"db38800b",
          4666 => x"84b6da34",
          4667 => x"810b84b6",
          4668 => x"dc34820b",
          4669 => x"83f89434",
          4670 => x"a80b83f8",
          4671 => x"9534820b",
          4672 => x"83f89223",
          4673 => x"795884b6",
          4674 => x"d8335784",
          4675 => x"b6d73356",
          4676 => x"84b6d633",
          4677 => x"557b547c",
          4678 => x"537a5283",
          4679 => x"e2d851ff",
          4680 => x"81e63f7d",
          4681 => x"84b6da34",
          4682 => x"800b84b6",
          4683 => x"dc347a83",
          4684 => x"f894347b",
          4685 => x"83f89223",
          4686 => x"7c83f895",
          4687 => x"348f3d0d",
          4688 => x"04800b84",
          4689 => x"b6da3481",
          4690 => x"0b84b6dc",
          4691 => x"34800b83",
          4692 => x"f89434a8",
          4693 => x"0b83f895",
          4694 => x"34800b83",
          4695 => x"f8922384",
          4696 => x"b7e73358",
          4697 => x"84b7e633",
          4698 => x"5784b7e5",
          4699 => x"33567955",
          4700 => x"7b547c53",
          4701 => x"7a5283e2",
          4702 => x"f451ff81",
          4703 => x"8b3f800b",
          4704 => x"84b7e533",
          4705 => x"5a5a7979",
          4706 => x"27a53879",
          4707 => x"1084b8b8",
          4708 => x"05702253",
          4709 => x"5983e38c",
          4710 => x"51ff80ec",
          4711 => x"3f811a70",
          4712 => x"81ff0684",
          4713 => x"b7e53352",
          4714 => x"5b59787a",
          4715 => x"26dd3883",
          4716 => x"d29451ff",
          4717 => x"80d23f7d",
          4718 => x"84b6da34",
          4719 => x"800b84b6",
          4720 => x"dc347a83",
          4721 => x"f894347b",
          4722 => x"83f89223",
          4723 => x"7c83f895",
          4724 => x"348f3d0d",
          4725 => x"04800b84",
          4726 => x"b6da3481",
          4727 => x"0b84b6dc",
          4728 => x"34810b83",
          4729 => x"f89434a8",
          4730 => x"0b83f895",
          4731 => x"34810b83",
          4732 => x"f8922383",
          4733 => x"f6c851ff",
          4734 => x"92ae3f84",
          4735 => x"b8e40852",
          4736 => x"83e39051",
          4737 => x"ff80813f",
          4738 => x"805983f6",
          4739 => x"c851ff92",
          4740 => x"973f7884",
          4741 => x"b8e40827",
          4742 => x"fda63883",
          4743 => x"f6c81933",
          4744 => x"5283e398",
          4745 => x"51feffe0",
          4746 => x"3f811970",
          4747 => x"81ff065a",
          4748 => x"5ad839f9",
          4749 => x"3d0d7a02",
          4750 => x"8405a705",
          4751 => x"3384b6d8",
          4752 => x"3383f895",
          4753 => x"3383f894",
          4754 => x"33727129",
          4755 => x"1286a7a0",
          4756 => x"801183f8",
          4757 => x"92225351",
          4758 => x"595c717c",
          4759 => x"29057083",
          4760 => x"ffff0683",
          4761 => x"f6ea3352",
          4762 => x"59515557",
          4763 => x"5772812e",
          4764 => x"81e93875",
          4765 => x"892e81f9",
          4766 => x"38758924",
          4767 => x"81b93875",
          4768 => x"812e8385",
          4769 => x"3875882e",
          4770 => x"82d53884",
          4771 => x"b6d83383",
          4772 => x"f8943383",
          4773 => x"f8953372",
          4774 => x"72290555",
          4775 => x"565484b6",
          4776 => x"e0163386",
          4777 => x"a7a08014",
          4778 => x"3484b6d8",
          4779 => x"3383f895",
          4780 => x"3383f892",
          4781 => x"22727129",
          4782 => x"125a5a56",
          4783 => x"537583f8",
          4784 => x"96183483",
          4785 => x"f8943373",
          4786 => x"71291658",
          4787 => x"5483f890",
          4788 => x"3386a7b0",
          4789 => x"80183484",
          4790 => x"b6d83370",
          4791 => x"81ff0683",
          4792 => x"f8922283",
          4793 => x"f8953372",
          4794 => x"72291157",
          4795 => x"5b575557",
          4796 => x"83f89033",
          4797 => x"8497b614",
          4798 => x"34811870",
          4799 => x"81ff0659",
          4800 => x"55737826",
          4801 => x"81993884",
          4802 => x"b6d93358",
          4803 => x"7781ea38",
          4804 => x"ff175372",
          4805 => x"83f89534",
          4806 => x"84b6db33",
          4807 => x"5372802e",
          4808 => x"8c3884b6",
          4809 => x"dc335776",
          4810 => x"802e80fb",
          4811 => x"38800b84",
          4812 => x"b8e40c89",
          4813 => x"3d0d0475",
          4814 => x"8d2e9738",
          4815 => x"758d2480",
          4816 => x"f738758a",
          4817 => x"2e098106",
          4818 => x"fec13881",
          4819 => x"528151f1",
          4820 => x"963f800b",
          4821 => x"83f89534",
          4822 => x"ffbe3983",
          4823 => x"f8961533",
          4824 => x"5384b6e0",
          4825 => x"13337434",
          4826 => x"75892e09",
          4827 => x"8106fe89",
          4828 => x"38805376",
          4829 => x"52a051fd",
          4830 => x"ba3f8113",
          4831 => x"7081ff06",
          4832 => x"54547283",
          4833 => x"26ff9138",
          4834 => x"7652a051",
          4835 => x"fda53f81",
          4836 => x"137081ff",
          4837 => x"06545483",
          4838 => x"7327d838",
          4839 => x"fefa3974",
          4840 => x"83f89534",
          4841 => x"fef23975",
          4842 => x"528351f9",
          4843 => x"de3f800b",
          4844 => x"84b8e40c",
          4845 => x"893d0d04",
          4846 => x"7580ff2e",
          4847 => x"098106fd",
          4848 => x"ca3883f8",
          4849 => x"95337081",
          4850 => x"ff0655ff",
          4851 => x"05537383",
          4852 => x"38735372",
          4853 => x"83f89534",
          4854 => x"7652a051",
          4855 => x"fcd53f83",
          4856 => x"f8953370",
          4857 => x"81ff0655",
          4858 => x"ff055373",
          4859 => x"fea53873",
          4860 => x"537283f8",
          4861 => x"9534fea0",
          4862 => x"39800b83",
          4863 => x"f8953481",
          4864 => x"528151ef",
          4865 => x"e23ffe90",
          4866 => x"39805275",
          4867 => x"51efd83f",
          4868 => x"fe8639e6",
          4869 => x"3d0d0280",
          4870 => x"f3053384",
          4871 => x"b7e00857",
          4872 => x"5975812e",
          4873 => x"81b83875",
          4874 => x"822e8382",
          4875 => x"38788a2e",
          4876 => x"84b53878",
          4877 => x"8a2482d1",
          4878 => x"3878882e",
          4879 => x"84b93878",
          4880 => x"892e888f",
          4881 => x"3884b6d8",
          4882 => x"3383f894",
          4883 => x"3383f895",
          4884 => x"33727229",
          4885 => x"05585e5c",
          4886 => x"84b6e019",
          4887 => x"3386a7a0",
          4888 => x"80173484",
          4889 => x"b6d83383",
          4890 => x"f8953383",
          4891 => x"f8922272",
          4892 => x"7129125a",
          4893 => x"5a424078",
          4894 => x"83f89618",
          4895 => x"3483f894",
          4896 => x"33607129",
          4897 => x"6205405a",
          4898 => x"83f89033",
          4899 => x"7f86a7b0",
          4900 => x"80053484",
          4901 => x"b6d83370",
          4902 => x"81ff0683",
          4903 => x"f8922283",
          4904 => x"f8953372",
          4905 => x"72291142",
          4906 => x"405d5859",
          4907 => x"83f89033",
          4908 => x"8497b61f",
          4909 => x"34811d70",
          4910 => x"81ff0642",
          4911 => x"58766126",
          4912 => x"81b83884",
          4913 => x"b6d9335a",
          4914 => x"7986f138",
          4915 => x"ff195675",
          4916 => x"83f89534",
          4917 => x"800b84b8",
          4918 => x"e40c9c3d",
          4919 => x"0d0478b7",
          4920 => x"2e848a38",
          4921 => x"b7792581",
          4922 => x"fd3878b8",
          4923 => x"2e9bb338",
          4924 => x"7880db2e",
          4925 => x"89cc3880",
          4926 => x"0b84b7e0",
          4927 => x"0c84b6d8",
          4928 => x"3383f894",
          4929 => x"3383f895",
          4930 => x"33727229",
          4931 => x"055e4040",
          4932 => x"84b6e019",
          4933 => x"3386a7a0",
          4934 => x"801d3484",
          4935 => x"b6d83383",
          4936 => x"f8953383",
          4937 => x"f8922272",
          4938 => x"71291241",
          4939 => x"5f595678",
          4940 => x"83f8961f",
          4941 => x"3483f894",
          4942 => x"33767129",
          4943 => x"195b5783",
          4944 => x"f8903386",
          4945 => x"a7b0801b",
          4946 => x"3484b6d8",
          4947 => x"337081ff",
          4948 => x"0683f892",
          4949 => x"2283f895",
          4950 => x"33727229",
          4951 => x"11444243",
          4952 => x"585983f8",
          4953 => x"90336084",
          4954 => x"97b60534",
          4955 => x"811f5877",
          4956 => x"81ff0641",
          4957 => x"607727fe",
          4958 => x"ca387783",
          4959 => x"f8953480",
          4960 => x"0b84b8e4",
          4961 => x"0c9c3d0d",
          4962 => x"04789b2e",
          4963 => x"82b73878",
          4964 => x"9b248381",
          4965 => x"38788d2e",
          4966 => x"098106fd",
          4967 => x"a838800b",
          4968 => x"83f89534",
          4969 => x"800b84b8",
          4970 => x"e40c9c3d",
          4971 => x"0d04789b",
          4972 => x"2e82aa38",
          4973 => x"d0195675",
          4974 => x"892684d0",
          4975 => x"3884b7e4",
          4976 => x"33811159",
          4977 => x"577784b7",
          4978 => x"e4347884",
          4979 => x"b7e81834",
          4980 => x"7781ff06",
          4981 => x"59800b84",
          4982 => x"b7e81a34",
          4983 => x"800b84b8",
          4984 => x"e40c9c3d",
          4985 => x"0d04789b",
          4986 => x"2efde938",
          4987 => x"800b84b7",
          4988 => x"e00c84b6",
          4989 => x"d83383f8",
          4990 => x"943383f8",
          4991 => x"95337272",
          4992 => x"29055e40",
          4993 => x"4084b6e0",
          4994 => x"193386a7",
          4995 => x"a0801d34",
          4996 => x"84b6d833",
          4997 => x"83f89533",
          4998 => x"83f89222",
          4999 => x"72712912",
          5000 => x"415f5956",
          5001 => x"7883f896",
          5002 => x"1f3483f8",
          5003 => x"94337671",
          5004 => x"29195b57",
          5005 => x"83f89033",
          5006 => x"86a7b080",
          5007 => x"1b3484b6",
          5008 => x"d8337081",
          5009 => x"ff0683f8",
          5010 => x"922283f8",
          5011 => x"95337272",
          5012 => x"29114442",
          5013 => x"43585983",
          5014 => x"f8903360",
          5015 => x"8497b605",
          5016 => x"34811f58",
          5017 => x"fe893981",
          5018 => x"528151ea",
          5019 => x"fa3f800b",
          5020 => x"83f89534",
          5021 => x"feae3984",
          5022 => x"b6d83383",
          5023 => x"f8953370",
          5024 => x"81ff0683",
          5025 => x"f8943373",
          5026 => x"71291286",
          5027 => x"a7a08005",
          5028 => x"83f89222",
          5029 => x"40515d72",
          5030 => x"7e290570",
          5031 => x"83ffff06",
          5032 => x"83f6ea33",
          5033 => x"5a51595a",
          5034 => x"5c75812e",
          5035 => x"86a43878",
          5036 => x"81ff06ff",
          5037 => x"1a575776",
          5038 => x"fc953876",
          5039 => x"567583f8",
          5040 => x"9534fc90",
          5041 => x"39800b84",
          5042 => x"b7e43480",
          5043 => x"0b84b7e5",
          5044 => x"34800b84",
          5045 => x"b7e63480",
          5046 => x"0b84b7e7",
          5047 => x"34810b84",
          5048 => x"b7e00c80",
          5049 => x"0b84b8e4",
          5050 => x"0c9c3d0d",
          5051 => x"0483f894",
          5052 => x"3384b8cc",
          5053 => x"3483f895",
          5054 => x"3384b8cd",
          5055 => x"3483f893",
          5056 => x"3384b8ce",
          5057 => x"34800b84",
          5058 => x"b7e00c80",
          5059 => x"0b84b8e4",
          5060 => x"0c9c3d0d",
          5061 => x"047880ff",
          5062 => x"2e098106",
          5063 => x"faa73883",
          5064 => x"f8943384",
          5065 => x"b6d83370",
          5066 => x"81ff0683",
          5067 => x"f8953370",
          5068 => x"81ff0672",
          5069 => x"75291186",
          5070 => x"a7a08005",
          5071 => x"83f89222",
          5072 => x"5c40727b",
          5073 => x"29057083",
          5074 => x"ffff0683",
          5075 => x"f6ea3344",
          5076 => x"5c435c42",
          5077 => x"5b5c7d81",
          5078 => x"2e85fe38",
          5079 => x"7881ff06",
          5080 => x"ff1a5856",
          5081 => x"75833875",
          5082 => x"577683f8",
          5083 => x"95347b81",
          5084 => x"ff067a81",
          5085 => x"ff067881",
          5086 => x"ff067272",
          5087 => x"29055f40",
          5088 => x"5b84b780",
          5089 => x"3386a7a0",
          5090 => x"801e3484",
          5091 => x"b6d83383",
          5092 => x"f8953383",
          5093 => x"f8922272",
          5094 => x"7129125a",
          5095 => x"5e4240a0",
          5096 => x"0b83f896",
          5097 => x"183483f8",
          5098 => x"94336071",
          5099 => x"2962055a",
          5100 => x"5683f890",
          5101 => x"3386a7b0",
          5102 => x"801a3484",
          5103 => x"b6d83370",
          5104 => x"81ff0683",
          5105 => x"f8922283",
          5106 => x"f8953372",
          5107 => x"72291143",
          5108 => x"5d5a5e59",
          5109 => x"83f89033",
          5110 => x"7f8497b6",
          5111 => x"0534811a",
          5112 => x"7081ff06",
          5113 => x"5c587c7b",
          5114 => x"2695ea38",
          5115 => x"84b6d933",
          5116 => x"5a7996d0",
          5117 => x"38ff1958",
          5118 => x"7783f895",
          5119 => x"3483f895",
          5120 => x"337081ff",
          5121 => x"0658ff05",
          5122 => x"56fdac39",
          5123 => x"78bb2e95",
          5124 => x"d83878bd",
          5125 => x"2e83d738",
          5126 => x"78bf2e95",
          5127 => x"a83884b7",
          5128 => x"e4335f7e",
          5129 => x"83f938ff",
          5130 => x"bf195675",
          5131 => x"b42684c8",
          5132 => x"38751010",
          5133 => x"83c5c005",
          5134 => x"58770804",
          5135 => x"800b83f8",
          5136 => x"95348052",
          5137 => x"8151e79f",
          5138 => x"3f800b84",
          5139 => x"b8e40c9c",
          5140 => x"3d0d0483",
          5141 => x"f8943384",
          5142 => x"b6d83370",
          5143 => x"81ff0683",
          5144 => x"f8953370",
          5145 => x"81ff0672",
          5146 => x"75291186",
          5147 => x"a7a08005",
          5148 => x"83f89222",
          5149 => x"5c41727b",
          5150 => x"29057083",
          5151 => x"ffff0683",
          5152 => x"f6ea3346",
          5153 => x"53455c59",
          5154 => x"5b5b7f81",
          5155 => x"2e82ef38",
          5156 => x"805c7a81",
          5157 => x"ff067a81",
          5158 => x"ff067a81",
          5159 => x"ff067272",
          5160 => x"29055c58",
          5161 => x"4084b780",
          5162 => x"3386a7a0",
          5163 => x"801b3484",
          5164 => x"b6d83383",
          5165 => x"f8953383",
          5166 => x"f8922272",
          5167 => x"7129125e",
          5168 => x"415e56a0",
          5169 => x"0b83f896",
          5170 => x"1c3483f8",
          5171 => x"94337671",
          5172 => x"291e5a5e",
          5173 => x"83f89033",
          5174 => x"86a7b080",
          5175 => x"1a3484b6",
          5176 => x"d8337081",
          5177 => x"ff0683f8",
          5178 => x"922283f8",
          5179 => x"95337272",
          5180 => x"29115b44",
          5181 => x"5a405983",
          5182 => x"f8903384",
          5183 => x"97b61834",
          5184 => x"60810570",
          5185 => x"81ff065b",
          5186 => x"587e7a26",
          5187 => x"81ac3884",
          5188 => x"b6d93358",
          5189 => x"7792fb38",
          5190 => x"ff195675",
          5191 => x"83f89534",
          5192 => x"811c7081",
          5193 => x"ff065d59",
          5194 => x"7b8326f7",
          5195 => x"a73883f8",
          5196 => x"943384b6",
          5197 => x"d83383f8",
          5198 => x"95337281",
          5199 => x"ff067281",
          5200 => x"ff067281",
          5201 => x"ff067272",
          5202 => x"2905545b",
          5203 => x"435b5b5b",
          5204 => x"84b78033",
          5205 => x"86a7a080",
          5206 => x"1b3484b6",
          5207 => x"d83383f8",
          5208 => x"953383f8",
          5209 => x"92227271",
          5210 => x"29125e41",
          5211 => x"5e56a00b",
          5212 => x"83f8961c",
          5213 => x"3483f894",
          5214 => x"33767129",
          5215 => x"1e5a5e83",
          5216 => x"f8903386",
          5217 => x"a7b0801a",
          5218 => x"3484b6d8",
          5219 => x"337081ff",
          5220 => x"0683f892",
          5221 => x"2283f895",
          5222 => x"33727229",
          5223 => x"115b445a",
          5224 => x"405983f8",
          5225 => x"90338497",
          5226 => x"b6183460",
          5227 => x"81057081",
          5228 => x"ff065b58",
          5229 => x"797f27fe",
          5230 => x"d6387783",
          5231 => x"f89534fe",
          5232 => x"df39820b",
          5233 => x"84b7e00c",
          5234 => x"800b84b8",
          5235 => x"e40c9c3d",
          5236 => x"0d0483f8",
          5237 => x"96173359",
          5238 => x"84b6e019",
          5239 => x"337a3483",
          5240 => x"f8953370",
          5241 => x"81ff0658",
          5242 => x"ff0556f9",
          5243 => x"ca39810b",
          5244 => x"84b7e634",
          5245 => x"800b84b8",
          5246 => x"e40c9c3d",
          5247 => x"0d0483f8",
          5248 => x"9617335b",
          5249 => x"84b6e01b",
          5250 => x"337c3483",
          5251 => x"f8943384",
          5252 => x"b6d83383",
          5253 => x"f895335b",
          5254 => x"5b5b805c",
          5255 => x"fcf43984",
          5256 => x"b7e8429c",
          5257 => x"3ddc1153",
          5258 => x"d80551ff",
          5259 => x"8ad83f84",
          5260 => x"b8e40880",
          5261 => x"2efbf038",
          5262 => x"84b7e533",
          5263 => x"8111575a",
          5264 => x"7584b7e5",
          5265 => x"34791083",
          5266 => x"fe064102",
          5267 => x"80ca0522",
          5268 => x"6184b8b8",
          5269 => x"0523fbcf",
          5270 => x"3983f896",
          5271 => x"17335c84",
          5272 => x"b6e01c33",
          5273 => x"7b3483f8",
          5274 => x"943384b6",
          5275 => x"d83383f8",
          5276 => x"95335b5b",
          5277 => x"5cf9e539",
          5278 => x"84b6d833",
          5279 => x"83f89433",
          5280 => x"83f89533",
          5281 => x"72722905",
          5282 => x"415d5b84",
          5283 => x"b6e01933",
          5284 => x"7f86a7a0",
          5285 => x"80053484",
          5286 => x"b6d83383",
          5287 => x"f8953383",
          5288 => x"f8922272",
          5289 => x"7129125a",
          5290 => x"435b5678",
          5291 => x"83f89618",
          5292 => x"3483f894",
          5293 => x"33767129",
          5294 => x"1b415e83",
          5295 => x"f8903360",
          5296 => x"86a7b080",
          5297 => x"053484b6",
          5298 => x"d8337081",
          5299 => x"ff0683f8",
          5300 => x"922283f8",
          5301 => x"95337272",
          5302 => x"2911415f",
          5303 => x"5a425a83",
          5304 => x"f8903384",
          5305 => x"97b61e34",
          5306 => x"811c7081",
          5307 => x"ff065c58",
          5308 => x"607b2690",
          5309 => x"a23884b6",
          5310 => x"d9335877",
          5311 => x"90e238ff",
          5312 => x"1a567583",
          5313 => x"f8953480",
          5314 => x"0b84b7e0",
          5315 => x"0c84b6db",
          5316 => x"33407f80",
          5317 => x"2ef3bd38",
          5318 => x"84b6dc33",
          5319 => x"5675f3b4",
          5320 => x"38785281",
          5321 => x"51eae43f",
          5322 => x"800b84b8",
          5323 => x"e40c9c3d",
          5324 => x"0d0484b8",
          5325 => x"cc3383f8",
          5326 => x"943484b8",
          5327 => x"cd3383f8",
          5328 => x"953484b8",
          5329 => x"ce335776",
          5330 => x"83f89223",
          5331 => x"ffb93983",
          5332 => x"f8943384",
          5333 => x"b8cc3483",
          5334 => x"f8953384",
          5335 => x"b8cd3483",
          5336 => x"f8933384",
          5337 => x"b8ce34ff",
          5338 => x"9e3984b7",
          5339 => x"e5335b7a",
          5340 => x"802eff93",
          5341 => x"3884b8b8",
          5342 => x"225d7c86",
          5343 => x"2e098106",
          5344 => x"ff853883",
          5345 => x"f8953381",
          5346 => x"055583f8",
          5347 => x"94338105",
          5348 => x"549b5383",
          5349 => x"e3a05294",
          5350 => x"3d705257",
          5351 => x"feee893f",
          5352 => x"7651feff",
          5353 => x"833f84b8",
          5354 => x"e40881ff",
          5355 => x"0683f6e8",
          5356 => x"33577605",
          5357 => x"4160a024",
          5358 => x"fecd3876",
          5359 => x"5283f6c8",
          5360 => x"51fefdce",
          5361 => x"3ffec039",
          5362 => x"800b84b7",
          5363 => x"e5335b58",
          5364 => x"7981ff06",
          5365 => x"5b777b27",
          5366 => x"fead3877",
          5367 => x"1084b8b8",
          5368 => x"05811133",
          5369 => x"574175b1",
          5370 => x"268aa538",
          5371 => x"75101083",
          5372 => x"c794055f",
          5373 => x"7e080484",
          5374 => x"b7e5335e",
          5375 => x"7d802e8f",
          5376 => x"a43883f8",
          5377 => x"943384b8",
          5378 => x"b9337171",
          5379 => x"31700970",
          5380 => x"9f2c7206",
          5381 => x"5a42595e",
          5382 => x"5c7583f8",
          5383 => x"9434fde7",
          5384 => x"3984b7e5",
          5385 => x"33567580",
          5386 => x"2e8ee738",
          5387 => x"84b8b933",
          5388 => x"ff057081",
          5389 => x"ff0684b6",
          5390 => x"d8335d57",
          5391 => x"5f757b27",
          5392 => x"fdc53875",
          5393 => x"83f89534",
          5394 => x"fdbd3980",
          5395 => x"0b83f895",
          5396 => x"3483f894",
          5397 => x"337081ff",
          5398 => x"065d577b",
          5399 => x"802efda7",
          5400 => x"38ff1756",
          5401 => x"7583f894",
          5402 => x"34fd9c39",
          5403 => x"800b83f8",
          5404 => x"953483f8",
          5405 => x"943384b6",
          5406 => x"d733ff05",
          5407 => x"57577676",
          5408 => x"25fd8438",
          5409 => x"81175675",
          5410 => x"83f89434",
          5411 => x"fcf93984",
          5412 => x"b7e53340",
          5413 => x"7f802e8d",
          5414 => x"e03883f8",
          5415 => x"953384b8",
          5416 => x"b9337171",
          5417 => x"31700970",
          5418 => x"9f2c7206",
          5419 => x"5a415942",
          5420 => x"5a7583f8",
          5421 => x"9534fccf",
          5422 => x"3984b7e5",
          5423 => x"335b7a80",
          5424 => x"2efcc438",
          5425 => x"84b8b822",
          5426 => x"4160992e",
          5427 => x"098106fc",
          5428 => x"b63884b6",
          5429 => x"d83383f8",
          5430 => x"953383f8",
          5431 => x"94337271",
          5432 => x"291286a7",
          5433 => x"a0801183",
          5434 => x"f8922243",
          5435 => x"515a5871",
          5436 => x"60290570",
          5437 => x"83ffff06",
          5438 => x"83f6e808",
          5439 => x"87fffe80",
          5440 => x"06425a5d",
          5441 => x"5d7e8482",
          5442 => x"802e92bf",
          5443 => x"38800b83",
          5444 => x"f6e934fb",
          5445 => x"f23984b7",
          5446 => x"e5335a79",
          5447 => x"802efbe7",
          5448 => x"3884b8b8",
          5449 => x"22587799",
          5450 => x"2e098106",
          5451 => x"fbd93881",
          5452 => x"0b83f6e9",
          5453 => x"34fbd039",
          5454 => x"84b7e533",
          5455 => x"5675802e",
          5456 => x"90be3884",
          5457 => x"b8b93383",
          5458 => x"f895335d",
          5459 => x"7c0584b6",
          5460 => x"d833ff11",
          5461 => x"595e5675",
          5462 => x"7d258338",
          5463 => x"75577683",
          5464 => x"f89534fb",
          5465 => x"a23984b7",
          5466 => x"e5335776",
          5467 => x"802e8cc8",
          5468 => x"3884b8b9",
          5469 => x"3383f894",
          5470 => x"33426105",
          5471 => x"84b6d733",
          5472 => x"ff115941",
          5473 => x"56756025",
          5474 => x"83387557",
          5475 => x"7683f894",
          5476 => x"34faf439",
          5477 => x"83e3ac51",
          5478 => x"fee8ed3f",
          5479 => x"800b84b7",
          5480 => x"e5335757",
          5481 => x"7676278b",
          5482 => x"c7387610",
          5483 => x"84b8b805",
          5484 => x"7022535a",
          5485 => x"83e38c51",
          5486 => x"fee8cd3f",
          5487 => x"81177081",
          5488 => x"ff0684b7",
          5489 => x"e5335858",
          5490 => x"58da3982",
          5491 => x"0b84b7e5",
          5492 => x"335f577d",
          5493 => x"802e8d38",
          5494 => x"84b8b822",
          5495 => x"56758326",
          5496 => x"83387557",
          5497 => x"81527681",
          5498 => x"ff0651d5",
          5499 => x"f33ffa97",
          5500 => x"3984b7e5",
          5501 => x"33578177",
          5502 => x"278eb738",
          5503 => x"84b8bb33",
          5504 => x"ff057081",
          5505 => x"ff0684b8",
          5506 => x"b933ff05",
          5507 => x"7081ff06",
          5508 => x"84b6d733",
          5509 => x"7081ff06",
          5510 => x"ff114043",
          5511 => x"525b595c",
          5512 => x"5c777e27",
          5513 => x"8338775a",
          5514 => x"7983f892",
          5515 => x"237681ff",
          5516 => x"06ff1858",
          5517 => x"5f777f27",
          5518 => x"83387757",
          5519 => x"7683f894",
          5520 => x"3484b6d8",
          5521 => x"33ff1157",
          5522 => x"407a6027",
          5523 => x"f9b4387a",
          5524 => x"567583f8",
          5525 => x"9534f9af",
          5526 => x"3984b7e5",
          5527 => x"335f7e80",
          5528 => x"2e8aef38",
          5529 => x"84b8b933",
          5530 => x"84b6d733",
          5531 => x"405b7a7f",
          5532 => x"26f99438",
          5533 => x"83f89433",
          5534 => x"84b6d833",
          5535 => x"7081ff06",
          5536 => x"83f89533",
          5537 => x"71742911",
          5538 => x"86a7a080",
          5539 => x"0583f892",
          5540 => x"225f4071",
          5541 => x"7e290570",
          5542 => x"83ffff06",
          5543 => x"83f6ea33",
          5544 => x"46525959",
          5545 => x"5f5d6081",
          5546 => x"2e84f038",
          5547 => x"7983ffff",
          5548 => x"06707c31",
          5549 => x"5d57807c",
          5550 => x"248efe38",
          5551 => x"84b6d733",
          5552 => x"56767627",
          5553 => x"8ed638ff",
          5554 => x"16567583",
          5555 => x"f892237c",
          5556 => x"81ff0670",
          5557 => x"7c314157",
          5558 => x"8060248e",
          5559 => x"e53884b6",
          5560 => x"d7335676",
          5561 => x"76278dee",
          5562 => x"38ff1656",
          5563 => x"7583f894",
          5564 => x"347e81ff",
          5565 => x"0683f892",
          5566 => x"22575780",
          5567 => x"5a767626",
          5568 => x"90387577",
          5569 => x"3181057e",
          5570 => x"81ff0671",
          5571 => x"71295c5e",
          5572 => x"5b795886",
          5573 => x"a7a0805b",
          5574 => x"86a7b080",
          5575 => x"7f81ff06",
          5576 => x"7f81ff06",
          5577 => x"7171291d",
          5578 => x"4258425c",
          5579 => x"797f27f7",
          5580 => x"d6388497",
          5581 => x"b61a57e0",
          5582 => x"e017335f",
          5583 => x"84b6e01f",
          5584 => x"337b7081",
          5585 => x"055d3476",
          5586 => x"70810558",
          5587 => x"337c7081",
          5588 => x"055e3481",
          5589 => x"1884b6d8",
          5590 => x"3384b6d7",
          5591 => x"33717129",
          5592 => x"1d43405e",
          5593 => x"58776027",
          5594 => x"f79d38e0",
          5595 => x"e017335f",
          5596 => x"84b6e01f",
          5597 => x"337b7081",
          5598 => x"055d3476",
          5599 => x"70810558",
          5600 => x"337c7081",
          5601 => x"055e3481",
          5602 => x"1884b6d8",
          5603 => x"3384b6d7",
          5604 => x"33717129",
          5605 => x"1d43405e",
          5606 => x"587f7826",
          5607 => x"ff9938f6",
          5608 => x"e63984b7",
          5609 => x"e5335675",
          5610 => x"802e87e0",
          5611 => x"38805284",
          5612 => x"b8b93351",
          5613 => x"d8b13ff6",
          5614 => x"ce39800b",
          5615 => x"84b6d833",
          5616 => x"ff1184b7",
          5617 => x"e5335d59",
          5618 => x"40587978",
          5619 => x"2e943884",
          5620 => x"b8b82256",
          5621 => x"75782e09",
          5622 => x"81068bbe",
          5623 => x"3883f895",
          5624 => x"33587681",
          5625 => x"ff0683f8",
          5626 => x"94337943",
          5627 => x"5c5c76ff",
          5628 => x"2e81ed38",
          5629 => x"84b6d733",
          5630 => x"407a6026",
          5631 => x"f689387e",
          5632 => x"81ff0656",
          5633 => x"607626f5",
          5634 => x"fe387b76",
          5635 => x"26617d27",
          5636 => x"075776f5",
          5637 => x"f2387a10",
          5638 => x"101b7090",
          5639 => x"29620586",
          5640 => x"a7a08011",
          5641 => x"701f5d5a",
          5642 => x"86a7b080",
          5643 => x"05798306",
          5644 => x"58515d75",
          5645 => x"8bac3879",
          5646 => x"83065776",
          5647 => x"8ba43883",
          5648 => x"f8903370",
          5649 => x"982b7190",
          5650 => x"2b077188",
          5651 => x"2b077107",
          5652 => x"797f5952",
          5653 => x"5f57777a",
          5654 => x"279e3880",
          5655 => x"77708405",
          5656 => x"590c7d76",
          5657 => x"70840558",
          5658 => x"0c797726",
          5659 => x"ee3884b6",
          5660 => x"d83384b6",
          5661 => x"d733415f",
          5662 => x"7e81ff06",
          5663 => x"6081ff06",
          5664 => x"83f89222",
          5665 => x"7d732964",
          5666 => x"05595959",
          5667 => x"5a777726",
          5668 => x"8c387678",
          5669 => x"311b707b",
          5670 => x"29620557",
          5671 => x"4075761d",
          5672 => x"57577676",
          5673 => x"26f4e038",
          5674 => x"83f89033",
          5675 => x"8497b618",
          5676 => x"595aa00b",
          5677 => x"e0e01934",
          5678 => x"79787081",
          5679 => x"055a3481",
          5680 => x"17577676",
          5681 => x"26f4c038",
          5682 => x"a00be0e0",
          5683 => x"19347978",
          5684 => x"7081055a",
          5685 => x"34811757",
          5686 => x"757727d6",
          5687 => x"38f4a839",
          5688 => x"ff1f7081",
          5689 => x"ff065d58",
          5690 => x"fe8a3983",
          5691 => x"f8903370",
          5692 => x"80f00671",
          5693 => x"842b80f0",
          5694 => x"0671842a",
          5695 => x"07585d57",
          5696 => x"7b80f02e",
          5697 => x"098106be",
          5698 => x"3880f20b",
          5699 => x"83f89034",
          5700 => x"81187081",
          5701 => x"ff065956",
          5702 => x"f5b63983",
          5703 => x"f8961733",
          5704 => x"5e84b6e0",
          5705 => x"1e337c34",
          5706 => x"83f89433",
          5707 => x"84b6d833",
          5708 => x"83f89222",
          5709 => x"84b6d733",
          5710 => x"425c5f5d",
          5711 => x"faee3983",
          5712 => x"f8903387",
          5713 => x"07567583",
          5714 => x"f8903481",
          5715 => x"187081ff",
          5716 => x"065956f4",
          5717 => x"fb3983f8",
          5718 => x"903381fd",
          5719 => x"06850756",
          5720 => x"7583f890",
          5721 => x"34e53983",
          5722 => x"f8903381",
          5723 => x"fb068307",
          5724 => x"567583f8",
          5725 => x"9034d439",
          5726 => x"83f89033",
          5727 => x"81f90681",
          5728 => x"07567583",
          5729 => x"f89034c3",
          5730 => x"3983f890",
          5731 => x"33819f06",
          5732 => x"90075675",
          5733 => x"83f89034",
          5734 => x"ffb13980",
          5735 => x"f10b83f8",
          5736 => x"90348118",
          5737 => x"7081ff06",
          5738 => x"5956f4a4",
          5739 => x"3983f890",
          5740 => x"33818f06",
          5741 => x"567583f8",
          5742 => x"9034ff8f",
          5743 => x"3983f890",
          5744 => x"33819f06",
          5745 => x"90075675",
          5746 => x"83f89034",
          5747 => x"fefd3983",
          5748 => x"f8903381",
          5749 => x"ef0680e0",
          5750 => x"07567583",
          5751 => x"f89034fe",
          5752 => x"ea3983f8",
          5753 => x"903381cf",
          5754 => x"0680c007",
          5755 => x"567583f8",
          5756 => x"9034fed7",
          5757 => x"3983f890",
          5758 => x"3381af06",
          5759 => x"a0075675",
          5760 => x"83f89034",
          5761 => x"fec53983",
          5762 => x"f8903381",
          5763 => x"fe068607",
          5764 => x"567583f8",
          5765 => x"9034feb3",
          5766 => x"3983f890",
          5767 => x"3381fc06",
          5768 => x"84075675",
          5769 => x"83f89034",
          5770 => x"fea13983",
          5771 => x"f8903381",
          5772 => x"fa068207",
          5773 => x"567583f8",
          5774 => x"9034fe8f",
          5775 => x"3983f890",
          5776 => x"3381f806",
          5777 => x"567583f8",
          5778 => x"9034fdff",
          5779 => x"3983f890",
          5780 => x"3380f007",
          5781 => x"567583f8",
          5782 => x"9034fdef",
          5783 => x"3983f890",
          5784 => x"3380f007",
          5785 => x"567583f8",
          5786 => x"9034fddf",
          5787 => x"3983f890",
          5788 => x"3381df06",
          5789 => x"80d00756",
          5790 => x"7583f890",
          5791 => x"34fdcc39",
          5792 => x"83f89033",
          5793 => x"81bf06b0",
          5794 => x"07567583",
          5795 => x"f89034fd",
          5796 => x"ba39800b",
          5797 => x"83f89534",
          5798 => x"80528151",
          5799 => x"d2c93fec",
          5800 => x"ff3984b8",
          5801 => x"cc3383f8",
          5802 => x"943484b8",
          5803 => x"cd3383f8",
          5804 => x"953484b8",
          5805 => x"ce335978",
          5806 => x"83f89223",
          5807 => x"800b84b7",
          5808 => x"e00ce8c7",
          5809 => x"39810b84",
          5810 => x"b7e73480",
          5811 => x"0b84b8e4",
          5812 => x"0c9c3d0d",
          5813 => x"047783f8",
          5814 => x"953483f8",
          5815 => x"95337081",
          5816 => x"ff0658ff",
          5817 => x"0556e7cf",
          5818 => x"3984b7e8",
          5819 => x"429c3ddc",
          5820 => x"1153d805",
          5821 => x"51fef98e",
          5822 => x"3f84b8e4",
          5823 => x"08a13884",
          5824 => x"b8e40884",
          5825 => x"b7e00c80",
          5826 => x"0b84b7e4",
          5827 => x"34800b84",
          5828 => x"b8e40c9c",
          5829 => x"3d0d0477",
          5830 => x"83f89534",
          5831 => x"efe93984",
          5832 => x"b7e53381",
          5833 => x"115c5c7a",
          5834 => x"84b7e534",
          5835 => x"7b1083fe",
          5836 => x"065d0280",
          5837 => x"ca052284",
          5838 => x"b8b81e23",
          5839 => x"800b84b7",
          5840 => x"e434ca39",
          5841 => x"800b83f8",
          5842 => x"95348052",
          5843 => x"8151d197",
          5844 => x"3f83f895",
          5845 => x"337081ff",
          5846 => x"0658ff05",
          5847 => x"56e6d839",
          5848 => x"800b83f8",
          5849 => x"95348052",
          5850 => x"8151d0fb",
          5851 => x"3fef9839",
          5852 => x"8a51feeb",
          5853 => x"e93fef8f",
          5854 => x"3983f895",
          5855 => x"33ff0570",
          5856 => x"09709f2c",
          5857 => x"7206585f",
          5858 => x"57f2a639",
          5859 => x"75528151",
          5860 => x"d93984b6",
          5861 => x"d8334075",
          5862 => x"6027eeeb",
          5863 => x"387583f8",
          5864 => x"9534eee3",
          5865 => x"3983f894",
          5866 => x"33ff0570",
          5867 => x"09709f2c",
          5868 => x"72065840",
          5869 => x"57f0e239",
          5870 => x"83f89433",
          5871 => x"810584b6",
          5872 => x"d733ff11",
          5873 => x"59595675",
          5874 => x"7825f3c0",
          5875 => x"387557f3",
          5876 => x"bb3984b6",
          5877 => x"d7337081",
          5878 => x"ff06585c",
          5879 => x"817726ee",
          5880 => x"a63883f8",
          5881 => x"943384b6",
          5882 => x"d8337081",
          5883 => x"ff0683f8",
          5884 => x"95337174",
          5885 => x"291186a7",
          5886 => x"a0800583",
          5887 => x"f892225f",
          5888 => x"5f717e29",
          5889 => x"057083ff",
          5890 => x"ff0683f6",
          5891 => x"ea335d5b",
          5892 => x"44425f5d",
          5893 => x"77812e81",
          5894 => x"f5387983",
          5895 => x"ffff06ff",
          5896 => x"115c5780",
          5897 => x"7b248489",
          5898 => x"3884b6d7",
          5899 => x"33567676",
          5900 => x"27839838",
          5901 => x"ff165675",
          5902 => x"83f89223",
          5903 => x"7c81ff06",
          5904 => x"ff115757",
          5905 => x"80762483",
          5906 => x"df3884b6",
          5907 => x"d7335676",
          5908 => x"762782ec",
          5909 => x"38ff1656",
          5910 => x"7583f894",
          5911 => x"347b81ff",
          5912 => x"0683f892",
          5913 => x"22575780",
          5914 => x"5a767626",
          5915 => x"90387577",
          5916 => x"3181057e",
          5917 => x"81ff0671",
          5918 => x"71295c5e",
          5919 => x"5f795886",
          5920 => x"a7a0805b",
          5921 => x"86a7b080",
          5922 => x"7c81ff06",
          5923 => x"7f81ff06",
          5924 => x"7171291d",
          5925 => x"4142425d",
          5926 => x"797e27ec",
          5927 => x"ea388497",
          5928 => x"b61a57e0",
          5929 => x"e017335e",
          5930 => x"84b6e01e",
          5931 => x"337b7081",
          5932 => x"055d3476",
          5933 => x"70810558",
          5934 => x"337d7081",
          5935 => x"055f3481",
          5936 => x"1884b6d8",
          5937 => x"3384b6d7",
          5938 => x"33717129",
          5939 => x"1d59415d",
          5940 => x"58777627",
          5941 => x"ecb138e0",
          5942 => x"e017335e",
          5943 => x"84b6e01e",
          5944 => x"337b7081",
          5945 => x"055d3476",
          5946 => x"70810558",
          5947 => x"337d7081",
          5948 => x"055f3481",
          5949 => x"1884b6d8",
          5950 => x"3384b6d7",
          5951 => x"33717129",
          5952 => x"1d59415d",
          5953 => x"58757826",
          5954 => x"ff9938eb",
          5955 => x"fa3983f8",
          5956 => x"9617335c",
          5957 => x"84b6e01c",
          5958 => x"337b3483",
          5959 => x"f8943384",
          5960 => x"b6d83383",
          5961 => x"f8922284",
          5962 => x"b6d7335f",
          5963 => x"5c5f5dfd",
          5964 => x"e93976eb",
          5965 => x"d23884b6",
          5966 => x"d7337081",
          5967 => x"ff06ff11",
          5968 => x"5c425876",
          5969 => x"61278338",
          5970 => x"765a7983",
          5971 => x"f8922377",
          5972 => x"81ff06ff",
          5973 => x"19585a80",
          5974 => x"7a278338",
          5975 => x"80577683",
          5976 => x"f8943484",
          5977 => x"b6d83370",
          5978 => x"81ff06ff",
          5979 => x"12525956",
          5980 => x"807827eb",
          5981 => x"8d388056",
          5982 => x"7583f895",
          5983 => x"34eb8839",
          5984 => x"83f89533",
          5985 => x"810584b6",
          5986 => x"d833ff11",
          5987 => x"59405675",
          5988 => x"7f25efca",
          5989 => x"387557ef",
          5990 => x"c5397581",
          5991 => x"2e098106",
          5992 => x"f4c03883",
          5993 => x"f8953370",
          5994 => x"81ff0683",
          5995 => x"f894337a",
          5996 => x"445d5d57",
          5997 => x"76ff2e09",
          5998 => x"8106f4b8",
          5999 => x"38f6a139",
          6000 => x"ff1d5675",
          6001 => x"83f89434",
          6002 => x"fd9339ff",
          6003 => x"1a567583",
          6004 => x"f89223fc",
          6005 => x"e7397c7b",
          6006 => x"31567583",
          6007 => x"f89434f2",
          6008 => x"9039777d",
          6009 => x"5856777a",
          6010 => x"26f58d38",
          6011 => x"80767081",
          6012 => x"05583483",
          6013 => x"f8903377",
          6014 => x"70810559",
          6015 => x"34757a26",
          6016 => x"f4ec3880",
          6017 => x"76708105",
          6018 => x"583483f8",
          6019 => x"90337770",
          6020 => x"81055934",
          6021 => x"797627d4",
          6022 => x"38f4d339",
          6023 => x"797b3156",
          6024 => x"7583f892",
          6025 => x"23f1a839",
          6026 => x"800b83f8",
          6027 => x"9434fcad",
          6028 => x"397e83f8",
          6029 => x"9223fc84",
          6030 => x"39800b83",
          6031 => x"f89223f1",
          6032 => x"8e39800b",
          6033 => x"83f89434",
          6034 => x"f1a73983",
          6035 => x"f8961833",
          6036 => x"5a84b6e0",
          6037 => x"1a337734",
          6038 => x"800b83f6",
          6039 => x"e934e9a7",
          6040 => x"39fd3d0d",
          6041 => x"02970533",
          6042 => x"84b6da33",
          6043 => x"54547280",
          6044 => x"2e903873",
          6045 => x"51db9c3f",
          6046 => x"800b84b8",
          6047 => x"e40c853d",
          6048 => x"0d047652",
          6049 => x"7351d7ab",
          6050 => x"3f800b84",
          6051 => x"b8e40c85",
          6052 => x"3d0d04f3",
          6053 => x"3d0d02bf",
          6054 => x"05335cff",
          6055 => x"0b83f6e8",
          6056 => x"337081ff",
          6057 => x"0683f6c8",
          6058 => x"11335855",
          6059 => x"55597480",
          6060 => x"2e80d638",
          6061 => x"81145675",
          6062 => x"83f6e834",
          6063 => x"74597884",
          6064 => x"b8e40c8f",
          6065 => x"3d0d0483",
          6066 => x"f6c40854",
          6067 => x"82537380",
          6068 => x"2e913873",
          6069 => x"73327030",
          6070 => x"71077009",
          6071 => x"709f2a56",
          6072 => x"5d5e5872",
          6073 => x"83f6c40c",
          6074 => x"ff598054",
          6075 => x"7b812e09",
          6076 => x"81068338",
          6077 => x"7b547b83",
          6078 => x"32703070",
          6079 => x"80257607",
          6080 => x"5c5c5d79",
          6081 => x"802e85c4",
          6082 => x"3884b6d8",
          6083 => x"3383f895",
          6084 => x"3383f894",
          6085 => x"33727129",
          6086 => x"1286a7a0",
          6087 => x"800583f8",
          6088 => x"92225b59",
          6089 => x"5d717929",
          6090 => x"057083ff",
          6091 => x"ff0683f6",
          6092 => x"e9335859",
          6093 => x"55587481",
          6094 => x"2e838c38",
          6095 => x"81f05473",
          6096 => x"86ee8080",
          6097 => x"34800b87",
          6098 => x"c098880c",
          6099 => x"87c09888",
          6100 => x"08567580",
          6101 => x"2ef63886",
          6102 => x"ee808408",
          6103 => x"577683f4",
          6104 => x"94153481",
          6105 => x"147081ff",
          6106 => x"06555581",
          6107 => x"f97427cf",
          6108 => x"38805483",
          6109 => x"f6841433",
          6110 => x"7081ff06",
          6111 => x"83f68e16",
          6112 => x"33585455",
          6113 => x"72762e85",
          6114 => x"c1387281",
          6115 => x"ff2e86b4",
          6116 => x"387483f6",
          6117 => x"98153475",
          6118 => x"81ff065a",
          6119 => x"7981ff2e",
          6120 => x"85cd3875",
          6121 => x"83f6a215",
          6122 => x"3483f684",
          6123 => x"143383f6",
          6124 => x"8e153481",
          6125 => x"147081ff",
          6126 => x"06555e89",
          6127 => x"7427ffb3",
          6128 => x"3883f68c",
          6129 => x"3370982b",
          6130 => x"70802558",
          6131 => x"56547583",
          6132 => x"f6bc3473",
          6133 => x"81ff0670",
          6134 => x"862a8132",
          6135 => x"70810651",
          6136 => x"54587280",
          6137 => x"2e85e738",
          6138 => x"810b83f6",
          6139 => x"bd347309",
          6140 => x"81065372",
          6141 => x"802e85e4",
          6142 => x"38810b83",
          6143 => x"f6be3480",
          6144 => x"0b83f6bd",
          6145 => x"3383f6c4",
          6146 => x"0883f6be",
          6147 => x"337083f6",
          6148 => x"c03383f6",
          6149 => x"bf335d5d",
          6150 => x"425e5c5e",
          6151 => x"5683f698",
          6152 => x"16335574",
          6153 => x"81ff2e8d",
          6154 => x"3883f6ac",
          6155 => x"16335473",
          6156 => x"802e8282",
          6157 => x"3883f6a2",
          6158 => x"16335372",
          6159 => x"81ff2e8b",
          6160 => x"3883f6ac",
          6161 => x"16335473",
          6162 => x"81ec3874",
          6163 => x"81ff0654",
          6164 => x"7381ff2e",
          6165 => x"8d3883f6",
          6166 => x"ac163353",
          6167 => x"72812e81",
          6168 => x"da387481",
          6169 => x"ff065372",
          6170 => x"81ff2e84",
          6171 => x"8c3883f6",
          6172 => x"ac163354",
          6173 => x"81742784",
          6174 => x"803883f6",
          6175 => x"b80887e8",
          6176 => x"0587c098",
          6177 => x"9c085454",
          6178 => x"73732783",
          6179 => x"ec38810b",
          6180 => x"87c0989c",
          6181 => x"0883f6b8",
          6182 => x"0c588116",
          6183 => x"7081ff06",
          6184 => x"57548976",
          6185 => x"27fef638",
          6186 => x"7683f6bf",
          6187 => x"347783f6",
          6188 => x"c034fe9e",
          6189 => x"1953729c",
          6190 => x"26828b38",
          6191 => x"72101083",
          6192 => x"c8dc055a",
          6193 => x"79080483",
          6194 => x"f6ec0854",
          6195 => x"73802e91",
          6196 => x"3883f414",
          6197 => x"87c0989c",
          6198 => x"085e5e7d",
          6199 => x"7d27fcdc",
          6200 => x"38800b83",
          6201 => x"f6ea3354",
          6202 => x"5472812e",
          6203 => x"83387454",
          6204 => x"7383f6ea",
          6205 => x"3487c098",
          6206 => x"9c0883f6",
          6207 => x"ec0c7381",
          6208 => x"ff065877",
          6209 => x"812e9438",
          6210 => x"83f89617",
          6211 => x"335484b6",
          6212 => x"e0143376",
          6213 => x"3481f054",
          6214 => x"fca53983",
          6215 => x"f6c40853",
          6216 => x"72802e82",
          6217 => x"9c387281",
          6218 => x"2e83f438",
          6219 => x"80c37634",
          6220 => x"81f054fc",
          6221 => x"8a398058",
          6222 => x"fee03980",
          6223 => x"74565783",
          6224 => x"597c812e",
          6225 => x"9b387977",
          6226 => x"2e098106",
          6227 => x"83b4387d",
          6228 => x"812e80ed",
          6229 => x"3879812e",
          6230 => x"80d73879",
          6231 => x"81ff0659",
          6232 => x"87772775",
          6233 => x"982b5454",
          6234 => x"728025a1",
          6235 => x"3873802e",
          6236 => x"9c388117",
          6237 => x"7081ff06",
          6238 => x"761081fe",
          6239 => x"06877227",
          6240 => x"71982b57",
          6241 => x"53575854",
          6242 => x"807324e1",
          6243 => x"38781010",
          6244 => x"10791005",
          6245 => x"7611832b",
          6246 => x"780583f2",
          6247 => x"f4057033",
          6248 => x"5b565478",
          6249 => x"87c0989c",
          6250 => x"0883f6b8",
          6251 => x"0c57fdea",
          6252 => x"3980597d",
          6253 => x"812effa8",
          6254 => x"387981ff",
          6255 => x"0659ffa0",
          6256 => x"398259ff",
          6257 => x"9b3978ff",
          6258 => x"2efa9f38",
          6259 => x"800b84b6",
          6260 => x"da335454",
          6261 => x"72812e83",
          6262 => x"e8387b82",
          6263 => x"32703070",
          6264 => x"80257607",
          6265 => x"4059567d",
          6266 => x"8a387b83",
          6267 => x"2e098106",
          6268 => x"f9cc3878",
          6269 => x"ff2ef9c6",
          6270 => x"38805372",
          6271 => x"10101083",
          6272 => x"f6f00570",
          6273 => x"335d5478",
          6274 => x"7c2e83ba",
          6275 => x"38811370",
          6276 => x"81ff0654",
          6277 => x"57937327",
          6278 => x"e23884b6",
          6279 => x"db335372",
          6280 => x"802ef99a",
          6281 => x"3884b6dc",
          6282 => x"335574f9",
          6283 => x"91387881",
          6284 => x"ff065282",
          6285 => x"51ccd43f",
          6286 => x"7884b8e4",
          6287 => x"0c8f3d0d",
          6288 => x"04be7634",
          6289 => x"81f054f9",
          6290 => x"f6397281",
          6291 => x"ff2e9238",
          6292 => x"83f6ac14",
          6293 => x"3381055b",
          6294 => x"7a83f6ac",
          6295 => x"1534fac9",
          6296 => x"39800b83",
          6297 => x"f6ac1534",
          6298 => x"ff0b83f6",
          6299 => x"981534ff",
          6300 => x"0b83f6a2",
          6301 => x"1534fab1",
          6302 => x"397481ff",
          6303 => x"06537281",
          6304 => x"ff2efc96",
          6305 => x"3883f6ac",
          6306 => x"16335581",
          6307 => x"7527fc8a",
          6308 => x"387781ff",
          6309 => x"06547381",
          6310 => x"2e098106",
          6311 => x"fbfc3883",
          6312 => x"f6b80881",
          6313 => x"fa0587c0",
          6314 => x"989c0854",
          6315 => x"55747327",
          6316 => x"fbe83887",
          6317 => x"c0989c08",
          6318 => x"83f6b80c",
          6319 => x"7681ff06",
          6320 => x"59fbd739",
          6321 => x"ff0b83f6",
          6322 => x"981534f9",
          6323 => x"ca397283",
          6324 => x"f6bd3473",
          6325 => x"09810653",
          6326 => x"72fa9e38",
          6327 => x"7283f6be",
          6328 => x"34800b83",
          6329 => x"f6bd3383",
          6330 => x"f6c40883",
          6331 => x"f6be3370",
          6332 => x"83f6c033",
          6333 => x"83f6bf33",
          6334 => x"5d5d425e",
          6335 => x"5c5e56fa",
          6336 => x"9c397982",
          6337 => x"2e098106",
          6338 => x"fccb387a",
          6339 => x"597a812e",
          6340 => x"fcce3879",
          6341 => x"812e0981",
          6342 => x"06fcc038",
          6343 => x"fd9339ef",
          6344 => x"763481f0",
          6345 => x"54f89839",
          6346 => x"800b84b6",
          6347 => x"db335754",
          6348 => x"75833881",
          6349 => x"547384b6",
          6350 => x"db34ff59",
          6351 => x"f7ac3980",
          6352 => x"0b84b6da",
          6353 => x"33585476",
          6354 => x"83388154",
          6355 => x"7384b6da",
          6356 => x"34ff59f7",
          6357 => x"95398153",
          6358 => x"83f6c408",
          6359 => x"842ef783",
          6360 => x"38840b83",
          6361 => x"f6c40cf6",
          6362 => x"ff3984b6",
          6363 => x"d7337081",
          6364 => x"ff06ff11",
          6365 => x"575a5480",
          6366 => x"79278338",
          6367 => x"80557483",
          6368 => x"f8922373",
          6369 => x"81ff06ff",
          6370 => x"15555380",
          6371 => x"73278338",
          6372 => x"80547383",
          6373 => x"f8943484",
          6374 => x"b6d83370",
          6375 => x"81ff0656",
          6376 => x"ff055380",
          6377 => x"75278338",
          6378 => x"80537283",
          6379 => x"f89534ff",
          6380 => x"59f6b739",
          6381 => x"81528351",
          6382 => x"ffbaa53f",
          6383 => x"ff59f6aa",
          6384 => x"397254fc",
          6385 => x"95398414",
          6386 => x"085283f6",
          6387 => x"c851fede",
          6388 => x"f63f810b",
          6389 => x"83f6e834",
          6390 => x"83f6c833",
          6391 => x"59fcbb39",
          6392 => x"803d0d81",
          6393 => x"51f5ac3f",
          6394 => x"823d0d04",
          6395 => x"fa3d0d80",
          6396 => x"0b83f2f0",
          6397 => x"08535702",
          6398 => x"a3053382",
          6399 => x"133483f2",
          6400 => x"f0085180",
          6401 => x"e0713485",
          6402 => x"0b83f2f0",
          6403 => x"085556fe",
          6404 => x"0b811534",
          6405 => x"800b86f0",
          6406 => x"80e83487",
          6407 => x"c0989c08",
          6408 => x"83f2f008",
          6409 => x"5580ce90",
          6410 => x"055387c0",
          6411 => x"989c0852",
          6412 => x"87c0989c",
          6413 => x"08517072",
          6414 => x"2ef63881",
          6415 => x"143387c0",
          6416 => x"989c0856",
          6417 => x"52747327",
          6418 => x"87387181",
          6419 => x"fe2edb38",
          6420 => x"87c098a4",
          6421 => x"0851ff55",
          6422 => x"70732780",
          6423 => x"c8387155",
          6424 => x"71ff2e80",
          6425 => x"c03887c0",
          6426 => x"989c0880",
          6427 => x"ce900553",
          6428 => x"87c0989c",
          6429 => x"085287c0",
          6430 => x"989c0855",
          6431 => x"74722ef6",
          6432 => x"38811433",
          6433 => x"87c0989c",
          6434 => x"08525270",
          6435 => x"73278738",
          6436 => x"7181ff2e",
          6437 => x"db3887c0",
          6438 => x"98a40855",
          6439 => x"72752683",
          6440 => x"38ff5271",
          6441 => x"55ff1670",
          6442 => x"81ff0657",
          6443 => x"5375802e",
          6444 => x"98387481",
          6445 => x"ff065271",
          6446 => x"fed53874",
          6447 => x"ff2e8a38",
          6448 => x"7684b8e4",
          6449 => x"0c883d0d",
          6450 => x"04810b84",
          6451 => x"b8e40c88",
          6452 => x"3d0d04fa",
          6453 => x"3d0d7902",
          6454 => x"8405a305",
          6455 => x"33565280",
          6456 => x"0b83f2f0",
          6457 => x"0873882b",
          6458 => x"87fc8080",
          6459 => x"06707598",
          6460 => x"2a075155",
          6461 => x"55577183",
          6462 => x"15347290",
          6463 => x"2a517084",
          6464 => x"15347190",
          6465 => x"2a567585",
          6466 => x"15347286",
          6467 => x"153483f2",
          6468 => x"f0085274",
          6469 => x"82133483",
          6470 => x"f2f00851",
          6471 => x"80e17134",
          6472 => x"850b83f2",
          6473 => x"f0085556",
          6474 => x"fe0b8115",
          6475 => x"34800b86",
          6476 => x"f080e834",
          6477 => x"87c0989c",
          6478 => x"0883f2f0",
          6479 => x"085580ce",
          6480 => x"90055387",
          6481 => x"c0989c08",
          6482 => x"5287c098",
          6483 => x"9c085170",
          6484 => x"722ef638",
          6485 => x"81143387",
          6486 => x"c0989c08",
          6487 => x"56527473",
          6488 => x"27873871",
          6489 => x"81fe2edb",
          6490 => x"3887c098",
          6491 => x"a40851ff",
          6492 => x"55707327",
          6493 => x"80c83871",
          6494 => x"5571ff2e",
          6495 => x"80c03887",
          6496 => x"c0989c08",
          6497 => x"80ce9005",
          6498 => x"5387c098",
          6499 => x"9c085287",
          6500 => x"c0989c08",
          6501 => x"5574722e",
          6502 => x"f6388114",
          6503 => x"3387c098",
          6504 => x"9c085252",
          6505 => x"70732787",
          6506 => x"387181ff",
          6507 => x"2edb3887",
          6508 => x"c098a408",
          6509 => x"55727526",
          6510 => x"8338ff52",
          6511 => x"7155ff16",
          6512 => x"7081ff06",
          6513 => x"57537580",
          6514 => x"2e80c738",
          6515 => x"7481ff06",
          6516 => x"5271fed4",
          6517 => x"38745170",
          6518 => x"81ff0656",
          6519 => x"75aa3880",
          6520 => x"c6147b84",
          6521 => x"80115552",
          6522 => x"52707327",
          6523 => x"92387170",
          6524 => x"81055333",
          6525 => x"71708105",
          6526 => x"53347271",
          6527 => x"26f03876",
          6528 => x"84b8e40c",
          6529 => x"883d0d04",
          6530 => x"810b84b8",
          6531 => x"e40c883d",
          6532 => x"0d04ff51",
          6533 => x"c239fa3d",
          6534 => x"0d790284",
          6535 => x"05a30533",
          6536 => x"5656800b",
          6537 => x"83f2f008",
          6538 => x"77882b87",
          6539 => x"fc808006",
          6540 => x"7079982a",
          6541 => x"07515555",
          6542 => x"57758315",
          6543 => x"3472902a",
          6544 => x"51708415",
          6545 => x"3475902a",
          6546 => x"52718515",
          6547 => x"34728615",
          6548 => x"347a83f2",
          6549 => x"f00880c6",
          6550 => x"11848013",
          6551 => x"56545551",
          6552 => x"70732797",
          6553 => x"38707081",
          6554 => x"05523372",
          6555 => x"70810554",
          6556 => x"34727126",
          6557 => x"f03883f2",
          6558 => x"f0085474",
          6559 => x"82153483",
          6560 => x"f2f00855",
          6561 => x"80e27534",
          6562 => x"850b83f2",
          6563 => x"f0085556",
          6564 => x"fe0b8115",
          6565 => x"34800b86",
          6566 => x"f080e834",
          6567 => x"87c0989c",
          6568 => x"0883f2f0",
          6569 => x"085580ce",
          6570 => x"90055387",
          6571 => x"c0989c08",
          6572 => x"5287c098",
          6573 => x"9c085170",
          6574 => x"722ef638",
          6575 => x"81143387",
          6576 => x"c0989c08",
          6577 => x"56527473",
          6578 => x"27873871",
          6579 => x"81fe2edb",
          6580 => x"3887c098",
          6581 => x"a40851ff",
          6582 => x"55707327",
          6583 => x"80c83871",
          6584 => x"5571ff2e",
          6585 => x"80c03887",
          6586 => x"c0989c08",
          6587 => x"80ce9005",
          6588 => x"5387c098",
          6589 => x"9c085287",
          6590 => x"c0989c08",
          6591 => x"5574722e",
          6592 => x"f6388114",
          6593 => x"3387c098",
          6594 => x"9c085252",
          6595 => x"70732787",
          6596 => x"387181ff",
          6597 => x"2edb3887",
          6598 => x"c098a408",
          6599 => x"55727526",
          6600 => x"8338ff52",
          6601 => x"7155ff16",
          6602 => x"7081ff06",
          6603 => x"57537580",
          6604 => x"2ea13874",
          6605 => x"81ff0652",
          6606 => x"71fed538",
          6607 => x"74517081",
          6608 => x"ff065473",
          6609 => x"802e8338",
          6610 => x"81577684",
          6611 => x"b8e40c88",
          6612 => x"3d0d04ff",
          6613 => x"51e839fb",
          6614 => x"3d0d83f2",
          6615 => x"f0085180",
          6616 => x"d0713485",
          6617 => x"0b83f2f0",
          6618 => x"085656fe",
          6619 => x"0b811634",
          6620 => x"800b86f0",
          6621 => x"80e83487",
          6622 => x"c0989c08",
          6623 => x"83f2f008",
          6624 => x"5680ce90",
          6625 => x"055487c0",
          6626 => x"989c0852",
          6627 => x"87c0989c",
          6628 => x"08537272",
          6629 => x"2ef63881",
          6630 => x"153387c0",
          6631 => x"989c0852",
          6632 => x"52707427",
          6633 => x"87387181",
          6634 => x"fe2edb38",
          6635 => x"87c098a4",
          6636 => x"0851ff53",
          6637 => x"70742780",
          6638 => x"c8387153",
          6639 => x"71ff2e80",
          6640 => x"c03887c0",
          6641 => x"989c0880",
          6642 => x"ce900553",
          6643 => x"87c0989c",
          6644 => x"085287c0",
          6645 => x"989c0851",
          6646 => x"70722ef6",
          6647 => x"38811533",
          6648 => x"87c0989c",
          6649 => x"08555273",
          6650 => x"73278738",
          6651 => x"7181ff2e",
          6652 => x"db3887c0",
          6653 => x"98a40851",
          6654 => x"72712683",
          6655 => x"38ff5271",
          6656 => x"53ff1670",
          6657 => x"81ff0657",
          6658 => x"5275802e",
          6659 => x"8a387281",
          6660 => x"ff065473",
          6661 => x"fed538ff",
          6662 => x"39803d0d",
          6663 => x"83e3e851",
          6664 => x"fed0d03f",
          6665 => x"823d0d04",
          6666 => x"f93d0d84",
          6667 => x"b8d4087a",
          6668 => x"7131832a",
          6669 => x"7083ffff",
          6670 => x"0670832b",
          6671 => x"73117033",
          6672 => x"81123371",
          6673 => x"8b2b7183",
          6674 => x"2b077711",
          6675 => x"70338112",
          6676 => x"3371982b",
          6677 => x"71902b07",
          6678 => x"5c544153",
          6679 => x"535d5759",
          6680 => x"52565753",
          6681 => x"80712481",
          6682 => x"af387216",
          6683 => x"82113383",
          6684 => x"1233718b",
          6685 => x"2b71832b",
          6686 => x"07760570",
          6687 => x"33811233",
          6688 => x"71982b71",
          6689 => x"902b0757",
          6690 => x"535c5259",
          6691 => x"56528071",
          6692 => x"24839e38",
          6693 => x"84133385",
          6694 => x"1433718b",
          6695 => x"2b71832b",
          6696 => x"07750576",
          6697 => x"882a5254",
          6698 => x"56577486",
          6699 => x"13347381",
          6700 => x"ff065473",
          6701 => x"87133484",
          6702 => x"b8d40870",
          6703 => x"17841233",
          6704 => x"85133371",
          6705 => x"882b0770",
          6706 => x"882a5c55",
          6707 => x"59545177",
          6708 => x"84143471",
          6709 => x"85143484",
          6710 => x"b8d40816",
          6711 => x"52800b86",
          6712 => x"1334800b",
          6713 => x"87133484",
          6714 => x"b8d40853",
          6715 => x"74841434",
          6716 => x"73851434",
          6717 => x"84b8d408",
          6718 => x"16703381",
          6719 => x"12337188",
          6720 => x"2b078280",
          6721 => x"80077088",
          6722 => x"2a585852",
          6723 => x"52747234",
          6724 => x"75811334",
          6725 => x"893d0d04",
          6726 => x"86123387",
          6727 => x"1333718b",
          6728 => x"2b71832b",
          6729 => x"07751184",
          6730 => x"16338517",
          6731 => x"3371882b",
          6732 => x"0770882a",
          6733 => x"58585451",
          6734 => x"53585871",
          6735 => x"84123472",
          6736 => x"85123484",
          6737 => x"b8d40870",
          6738 => x"16841133",
          6739 => x"85123371",
          6740 => x"8b2b7183",
          6741 => x"2b07565a",
          6742 => x"5a527205",
          6743 => x"86123387",
          6744 => x"13337188",
          6745 => x"2b077088",
          6746 => x"2a525559",
          6747 => x"52778613",
          6748 => x"34728713",
          6749 => x"3484b8d4",
          6750 => x"08157033",
          6751 => x"81123371",
          6752 => x"882b0781",
          6753 => x"ffff0670",
          6754 => x"882a5a5a",
          6755 => x"54527672",
          6756 => x"34778113",
          6757 => x"3484b8d4",
          6758 => x"08701770",
          6759 => x"33811233",
          6760 => x"718b2b71",
          6761 => x"832b0774",
          6762 => x"05703381",
          6763 => x"12337188",
          6764 => x"2b077083",
          6765 => x"2b8ffff8",
          6766 => x"0677057b",
          6767 => x"882a5452",
          6768 => x"53545c5a",
          6769 => x"57545277",
          6770 => x"82143473",
          6771 => x"83143484",
          6772 => x"b8d40870",
          6773 => x"17703381",
          6774 => x"1233718b",
          6775 => x"2b71832b",
          6776 => x"07740570",
          6777 => x"33811233",
          6778 => x"71882b07",
          6779 => x"81ffff06",
          6780 => x"70882a5f",
          6781 => x"5253555a",
          6782 => x"57545277",
          6783 => x"73347081",
          6784 => x"143484b8",
          6785 => x"d4087017",
          6786 => x"82113383",
          6787 => x"1233718b",
          6788 => x"2b71832b",
          6789 => x"07740570",
          6790 => x"33811233",
          6791 => x"71982b71",
          6792 => x"902b0758",
          6793 => x"535d525a",
          6794 => x"57535370",
          6795 => x"8025fce4",
          6796 => x"38713381",
          6797 => x"13337188",
          6798 => x"2b078280",
          6799 => x"80077088",
          6800 => x"2a595954",
          6801 => x"76753477",
          6802 => x"81163484",
          6803 => x"b8d40870",
          6804 => x"17703381",
          6805 => x"1233718b",
          6806 => x"2b71832b",
          6807 => x"07740582",
          6808 => x"14338315",
          6809 => x"3371882b",
          6810 => x"0770882a",
          6811 => x"575c5c52",
          6812 => x"58565253",
          6813 => x"72821534",
          6814 => x"75831534",
          6815 => x"893d0d04",
          6816 => x"f93d0d79",
          6817 => x"84b8d408",
          6818 => x"58587680",
          6819 => x"2e8f3877",
          6820 => x"802e8638",
          6821 => x"7751fb90",
          6822 => x"3f893d0d",
          6823 => x"0484fff4",
          6824 => x"0b84b8d4",
          6825 => x"0ca0800b",
          6826 => x"84b8d023",
          6827 => x"82808053",
          6828 => x"765284ff",
          6829 => x"f451fed3",
          6830 => x"c63f84b8",
          6831 => x"d4085576",
          6832 => x"7534810b",
          6833 => x"81163484",
          6834 => x"b8d40854",
          6835 => x"76841534",
          6836 => x"810b8515",
          6837 => x"3484b8d4",
          6838 => x"08567686",
          6839 => x"1734810b",
          6840 => x"87173484",
          6841 => x"b8d40884",
          6842 => x"b8d022ff",
          6843 => x"05fe8080",
          6844 => x"077083ff",
          6845 => x"ff067088",
          6846 => x"2a585155",
          6847 => x"56748817",
          6848 => x"34738917",
          6849 => x"3484b8d0",
          6850 => x"22701010",
          6851 => x"1084b8d4",
          6852 => x"0805f805",
          6853 => x"55557682",
          6854 => x"1534810b",
          6855 => x"831534fe",
          6856 => x"ee39f73d",
          6857 => x"0d7b5280",
          6858 => x"53815184",
          6859 => x"72278e38",
          6860 => x"fb12832a",
          6861 => x"82057083",
          6862 => x"ffff0651",
          6863 => x"517083ff",
          6864 => x"ff0684b8",
          6865 => x"d4088411",
          6866 => x"33851233",
          6867 => x"71882b07",
          6868 => x"7052595a",
          6869 => x"585581ff",
          6870 => x"ff547580",
          6871 => x"2e80cc38",
          6872 => x"75101010",
          6873 => x"17703381",
          6874 => x"12337188",
          6875 => x"2b077081",
          6876 => x"ffff0679",
          6877 => x"317083ff",
          6878 => x"ff06707a",
          6879 => x"2756535c",
          6880 => x"5c545272",
          6881 => x"74278a38",
          6882 => x"70802e85",
          6883 => x"38757355",
          6884 => x"58841233",
          6885 => x"85133371",
          6886 => x"882b0757",
          6887 => x"5a75c138",
          6888 => x"7381ffff",
          6889 => x"2e853877",
          6890 => x"74545680",
          6891 => x"76832b78",
          6892 => x"11703381",
          6893 => x"12337188",
          6894 => x"2b077081",
          6895 => x"ffff0656",
          6896 => x"565d5659",
          6897 => x"5970792e",
          6898 => x"83388159",
          6899 => x"80517473",
          6900 => x"26828d38",
          6901 => x"78517880",
          6902 => x"2e828538",
          6903 => x"72752e82",
          6904 => x"88387416",
          6905 => x"70832b78",
          6906 => x"11748280",
          6907 => x"80077088",
          6908 => x"2a5b5c56",
          6909 => x"565a7674",
          6910 => x"34788115",
          6911 => x"3484b8d4",
          6912 => x"08157688",
          6913 => x"2a535371",
          6914 => x"82143475",
          6915 => x"83143484",
          6916 => x"b8d40870",
          6917 => x"19703381",
          6918 => x"12337188",
          6919 => x"2b077083",
          6920 => x"2b8ffff8",
          6921 => x"0674057e",
          6922 => x"83ffff06",
          6923 => x"70882a5c",
          6924 => x"58535759",
          6925 => x"52527582",
          6926 => x"12347281",
          6927 => x"ff065372",
          6928 => x"83123484",
          6929 => x"b8d40818",
          6930 => x"54757434",
          6931 => x"72811534",
          6932 => x"84b8d408",
          6933 => x"70198611",
          6934 => x"33871233",
          6935 => x"718b2b71",
          6936 => x"832b0774",
          6937 => x"05585c5c",
          6938 => x"53577584",
          6939 => x"15347285",
          6940 => x"153484b8",
          6941 => x"d4087016",
          6942 => x"55780586",
          6943 => x"11338712",
          6944 => x"3371882b",
          6945 => x"0770882a",
          6946 => x"54545859",
          6947 => x"70861534",
          6948 => x"71871534",
          6949 => x"84b8d408",
          6950 => x"70198411",
          6951 => x"33851233",
          6952 => x"718b2b71",
          6953 => x"832b0774",
          6954 => x"05585a5c",
          6955 => x"5a527586",
          6956 => x"15347287",
          6957 => x"153484b8",
          6958 => x"d4087016",
          6959 => x"55780584",
          6960 => x"11338512",
          6961 => x"3371882b",
          6962 => x"0770882a",
          6963 => x"545c5759",
          6964 => x"70841534",
          6965 => x"79851534",
          6966 => x"84b8d408",
          6967 => x"18840551",
          6968 => x"7084b8e4",
          6969 => x"0c8b3d0d",
          6970 => x"04861433",
          6971 => x"87153371",
          6972 => x"8b2b7183",
          6973 => x"2b077905",
          6974 => x"84173385",
          6975 => x"18337188",
          6976 => x"2b077088",
          6977 => x"2a5a5b59",
          6978 => x"53545274",
          6979 => x"84123476",
          6980 => x"85123484",
          6981 => x"b8d40870",
          6982 => x"19841133",
          6983 => x"85123371",
          6984 => x"8b2b7183",
          6985 => x"2b077405",
          6986 => x"86143387",
          6987 => x"15337188",
          6988 => x"2b077088",
          6989 => x"2a585d5f",
          6990 => x"52565b57",
          6991 => x"5270861a",
          6992 => x"3476871a",
          6993 => x"3484b8d4",
          6994 => x"08187033",
          6995 => x"81123371",
          6996 => x"882b0781",
          6997 => x"ffff0670",
          6998 => x"882a5957",
          6999 => x"54577577",
          7000 => x"34748118",
          7001 => x"3484b8d4",
          7002 => x"08188405",
          7003 => x"51fef139",
          7004 => x"f93d0d79",
          7005 => x"84b8d408",
          7006 => x"58587680",
          7007 => x"2ea03877",
          7008 => x"54778a38",
          7009 => x"7384b8e4",
          7010 => x"0c893d0d",
          7011 => x"047751fb",
          7012 => x"913f84b8",
          7013 => x"e40884b8",
          7014 => x"e40c893d",
          7015 => x"0d0484ff",
          7016 => x"f40b84b8",
          7017 => x"d40ca080",
          7018 => x"0b84b8d0",
          7019 => x"23828080",
          7020 => x"53765284",
          7021 => x"fff451fe",
          7022 => x"cdc53f84",
          7023 => x"b8d40855",
          7024 => x"76753481",
          7025 => x"0b811634",
          7026 => x"84b8d408",
          7027 => x"54768415",
          7028 => x"34810b85",
          7029 => x"153484b8",
          7030 => x"d4085676",
          7031 => x"86173481",
          7032 => x"0b871734",
          7033 => x"84b8d408",
          7034 => x"84b8d022",
          7035 => x"ff05fe80",
          7036 => x"80077083",
          7037 => x"ffff0670",
          7038 => x"882a5851",
          7039 => x"55567488",
          7040 => x"17347389",
          7041 => x"173484b8",
          7042 => x"d0227010",
          7043 => x"101084b8",
          7044 => x"d40805f8",
          7045 => x"05555576",
          7046 => x"82153481",
          7047 => x"0b831534",
          7048 => x"77547780",
          7049 => x"2efedd38",
          7050 => x"fee339ed",
          7051 => x"3d0d6567",
          7052 => x"415f8070",
          7053 => x"84b8d408",
          7054 => x"59454176",
          7055 => x"612e84aa",
          7056 => x"387e802e",
          7057 => x"85af387f",
          7058 => x"802e88d7",
          7059 => x"38815484",
          7060 => x"60278f38",
          7061 => x"7ffb0583",
          7062 => x"2a820570",
          7063 => x"83ffff06",
          7064 => x"55587383",
          7065 => x"ffff067f",
          7066 => x"7831832a",
          7067 => x"7083ffff",
          7068 => x"0670832b",
          7069 => x"7a117033",
          7070 => x"81123371",
          7071 => x"882b0770",
          7072 => x"75317083",
          7073 => x"ffff0670",
          7074 => x"101010fc",
          7075 => x"0573832b",
          7076 => x"61117033",
          7077 => x"81123371",
          7078 => x"882b0770",
          7079 => x"902b7090",
          7080 => x"2c534245",
          7081 => x"46445354",
          7082 => x"43445c48",
          7083 => x"59525e5f",
          7084 => x"42807a24",
          7085 => x"85fd3882",
          7086 => x"15338316",
          7087 => x"3371882b",
          7088 => x"07701010",
          7089 => x"10197033",
          7090 => x"81123371",
          7091 => x"982b7190",
          7092 => x"2b07535c",
          7093 => x"53565656",
          7094 => x"80742485",
          7095 => x"c9387a62",
          7096 => x"2782f638",
          7097 => x"631b5877",
          7098 => x"622e87a2",
          7099 => x"3860802e",
          7100 => x"85f93860",
          7101 => x"1b587762",
          7102 => x"2587be38",
          7103 => x"63185961",
          7104 => x"792492f7",
          7105 => x"38761e70",
          7106 => x"33811233",
          7107 => x"718b2b71",
          7108 => x"832b077a",
          7109 => x"11703381",
          7110 => x"12337198",
          7111 => x"2b71902b",
          7112 => x"07474359",
          7113 => x"5253575b",
          7114 => x"58806024",
          7115 => x"8cba3876",
          7116 => x"1e821133",
          7117 => x"83123371",
          7118 => x"8b2b7183",
          7119 => x"2b077a11",
          7120 => x"86113387",
          7121 => x"1233718b",
          7122 => x"2b71832b",
          7123 => x"077e0584",
          7124 => x"14338515",
          7125 => x"3371882b",
          7126 => x"0770882a",
          7127 => x"59574852",
          7128 => x"5b415853",
          7129 => x"5c595677",
          7130 => x"841d3479",
          7131 => x"851d3484",
          7132 => x"b8d40870",
          7133 => x"17841133",
          7134 => x"85123371",
          7135 => x"8b2b7183",
          7136 => x"2b077405",
          7137 => x"86143387",
          7138 => x"15337188",
          7139 => x"2b077088",
          7140 => x"2a5f425e",
          7141 => x"52405741",
          7142 => x"57778616",
          7143 => x"347b8716",
          7144 => x"3484b8d4",
          7145 => x"08167033",
          7146 => x"81123371",
          7147 => x"882b0781",
          7148 => x"ffff0670",
          7149 => x"882a5a5c",
          7150 => x"5e597679",
          7151 => x"3479811a",
          7152 => x"3484b8d4",
          7153 => x"08701f82",
          7154 => x"11338312",
          7155 => x"33718b2b",
          7156 => x"71832b07",
          7157 => x"74057333",
          7158 => x"81153371",
          7159 => x"882b0770",
          7160 => x"882a415c",
          7161 => x"455d5f5a",
          7162 => x"55557979",
          7163 => x"3475811a",
          7164 => x"3484b8d4",
          7165 => x"08701f70",
          7166 => x"33811233",
          7167 => x"718b2b71",
          7168 => x"832b0774",
          7169 => x"05821433",
          7170 => x"83153371",
          7171 => x"882b0770",
          7172 => x"882a415c",
          7173 => x"455d5f5a",
          7174 => x"55557982",
          7175 => x"1a347583",
          7176 => x"1a3484b8",
          7177 => x"d408701f",
          7178 => x"82113383",
          7179 => x"12337188",
          7180 => x"2b076657",
          7181 => x"62567083",
          7182 => x"2b42525a",
          7183 => x"5d7e0584",
          7184 => x"0551fec4",
          7185 => x"fd3f84b8",
          7186 => x"d4081e84",
          7187 => x"05616505",
          7188 => x"1c7083ff",
          7189 => x"ff065d44",
          7190 => x"5f7a6226",
          7191 => x"81b6387e",
          7192 => x"547384b8",
          7193 => x"e40c953d",
          7194 => x"0d0484ff",
          7195 => x"f40b84b8",
          7196 => x"d40ca080",
          7197 => x"0b84b8d0",
          7198 => x"23828080",
          7199 => x"53605284",
          7200 => x"fff451fe",
          7201 => x"c7f93f84",
          7202 => x"b8d4085e",
          7203 => x"607e3481",
          7204 => x"0b811f34",
          7205 => x"84b8d408",
          7206 => x"5d60841e",
          7207 => x"34810b85",
          7208 => x"1e3484b8",
          7209 => x"d4085c60",
          7210 => x"861d3481",
          7211 => x"0b871d34",
          7212 => x"84b8d408",
          7213 => x"84b8d022",
          7214 => x"ff05fe80",
          7215 => x"80077083",
          7216 => x"ffff0670",
          7217 => x"882a5c5a",
          7218 => x"5b577888",
          7219 => x"18347789",
          7220 => x"183484b8",
          7221 => x"d0227010",
          7222 => x"101084b8",
          7223 => x"d40805f8",
          7224 => x"05555660",
          7225 => x"82153481",
          7226 => x"0b831534",
          7227 => x"84b8d408",
          7228 => x"577efad3",
          7229 => x"3876802e",
          7230 => x"828c387e",
          7231 => x"547f802e",
          7232 => x"fedf387f",
          7233 => x"51f49b3f",
          7234 => x"84b8e408",
          7235 => x"84b8e40c",
          7236 => x"953d0d04",
          7237 => x"611c84b8",
          7238 => x"d4087183",
          7239 => x"2b71115e",
          7240 => x"447f0570",
          7241 => x"33811233",
          7242 => x"71882b07",
          7243 => x"81ffff06",
          7244 => x"70882a48",
          7245 => x"445b5e40",
          7246 => x"637b3460",
          7247 => x"811c3461",
          7248 => x"84b8d408",
          7249 => x"057c882a",
          7250 => x"57587582",
          7251 => x"19347b83",
          7252 => x"193484b8",
          7253 => x"d408701f",
          7254 => x"70338112",
          7255 => x"3371882b",
          7256 => x"0770832b",
          7257 => x"8ffff806",
          7258 => x"74056483",
          7259 => x"ffff0670",
          7260 => x"882a4a5c",
          7261 => x"47575e5b",
          7262 => x"5d636382",
          7263 => x"05347681",
          7264 => x"ff064160",
          7265 => x"63830534",
          7266 => x"84b8d408",
          7267 => x"1e5b637b",
          7268 => x"3460811c",
          7269 => x"346184b8",
          7270 => x"d4080584",
          7271 => x"0551ed88",
          7272 => x"3f7e54fd",
          7273 => x"bc397b75",
          7274 => x"317083ff",
          7275 => x"ff064254",
          7276 => x"faac3977",
          7277 => x"81ffff06",
          7278 => x"76317083",
          7279 => x"ffff0682",
          7280 => x"17338318",
          7281 => x"3371882b",
          7282 => x"07701010",
          7283 => x"101b7033",
          7284 => x"81123371",
          7285 => x"982b7190",
          7286 => x"2b07535e",
          7287 => x"53545858",
          7288 => x"45547380",
          7289 => x"25f9f738",
          7290 => x"ffbc3961",
          7291 => x"7824fa83",
          7292 => x"38807a24",
          7293 => x"8b8f3877",
          7294 => x"83ffff06",
          7295 => x"5b617b27",
          7296 => x"fcdd38fe",
          7297 => x"8f3984ff",
          7298 => x"f40b84b8",
          7299 => x"d40ca080",
          7300 => x"0b84b8d0",
          7301 => x"23828080",
          7302 => x"537e5284",
          7303 => x"fff451fe",
          7304 => x"c4dd3f84",
          7305 => x"b8d4085a",
          7306 => x"7e7a3481",
          7307 => x"0b811b34",
          7308 => x"84b8d408",
          7309 => x"597e841a",
          7310 => x"34810b85",
          7311 => x"1a3484b8",
          7312 => x"d408587e",
          7313 => x"86193481",
          7314 => x"0b871934",
          7315 => x"84b8d408",
          7316 => x"84b8d022",
          7317 => x"ff05fe80",
          7318 => x"80077083",
          7319 => x"ffff0670",
          7320 => x"882a5856",
          7321 => x"57447464",
          7322 => x"88053473",
          7323 => x"64890534",
          7324 => x"84b8d022",
          7325 => x"70101010",
          7326 => x"84b8d408",
          7327 => x"05f80542",
          7328 => x"437e6182",
          7329 => x"05348161",
          7330 => x"830534fc",
          7331 => x"ee39807a",
          7332 => x"2483de38",
          7333 => x"6183ffff",
          7334 => x"065b617b",
          7335 => x"27fbc038",
          7336 => x"fcf23976",
          7337 => x"802e82bd",
          7338 => x"387e51ea",
          7339 => x"fb3f7f54",
          7340 => x"7384b8e4",
          7341 => x"0c953d0d",
          7342 => x"04761e82",
          7343 => x"11338312",
          7344 => x"33718b2b",
          7345 => x"71832b07",
          7346 => x"7a118611",
          7347 => x"33871233",
          7348 => x"718b2b71",
          7349 => x"832b077e",
          7350 => x"05841433",
          7351 => x"85153371",
          7352 => x"882b0770",
          7353 => x"882a4344",
          7354 => x"45565b46",
          7355 => x"58535c45",
          7356 => x"56786484",
          7357 => x"05347a64",
          7358 => x"85053484",
          7359 => x"b8d40870",
          7360 => x"17841133",
          7361 => x"85123371",
          7362 => x"8b2b7183",
          7363 => x"2b077405",
          7364 => x"86143387",
          7365 => x"15337188",
          7366 => x"2b077088",
          7367 => x"2a5b4142",
          7368 => x"485d595d",
          7369 => x"41736486",
          7370 => x"05347a64",
          7371 => x"87053484",
          7372 => x"b8d40816",
          7373 => x"70338112",
          7374 => x"3371882b",
          7375 => x"0781ffff",
          7376 => x"0670882a",
          7377 => x"5f5c5a5d",
          7378 => x"7b7d3479",
          7379 => x"811e3484",
          7380 => x"b8d40870",
          7381 => x"1f821133",
          7382 => x"83123371",
          7383 => x"8b2b7183",
          7384 => x"2b077405",
          7385 => x"73338115",
          7386 => x"3371882b",
          7387 => x"0770882a",
          7388 => x"5e5c5e40",
          7389 => x"43574554",
          7390 => x"767c3475",
          7391 => x"811d3484",
          7392 => x"b8d40870",
          7393 => x"1f703381",
          7394 => x"1233718b",
          7395 => x"2b71832b",
          7396 => x"07740582",
          7397 => x"14338315",
          7398 => x"3371882b",
          7399 => x"0770882a",
          7400 => x"4047405b",
          7401 => x"405c5555",
          7402 => x"78821834",
          7403 => x"60831834",
          7404 => x"84b8d408",
          7405 => x"701f8211",
          7406 => x"33831233",
          7407 => x"71882b07",
          7408 => x"66576256",
          7409 => x"70832b42",
          7410 => x"52585d7e",
          7411 => x"05840551",
          7412 => x"febdef3f",
          7413 => x"84b8d408",
          7414 => x"1e840578",
          7415 => x"83ffff06",
          7416 => x"5c5ffc99",
          7417 => x"3984fff4",
          7418 => x"0b84b8d4",
          7419 => x"0ca0800b",
          7420 => x"84b8d023",
          7421 => x"82808053",
          7422 => x"7f5284ff",
          7423 => x"f451fec0",
          7424 => x"fe3f84b8",
          7425 => x"d408567f",
          7426 => x"7634810b",
          7427 => x"81173484",
          7428 => x"b8d40855",
          7429 => x"7f841634",
          7430 => x"810b8516",
          7431 => x"3484b8d4",
          7432 => x"08547f86",
          7433 => x"1534810b",
          7434 => x"87153484",
          7435 => x"b8d40884",
          7436 => x"b8d022ff",
          7437 => x"05fe8080",
          7438 => x"077083ff",
          7439 => x"ff067088",
          7440 => x"2a454344",
          7441 => x"5e61881f",
          7442 => x"3460891f",
          7443 => x"3484b8d0",
          7444 => x"22701010",
          7445 => x"1084b8d4",
          7446 => x"0805f805",
          7447 => x"5c5d7f82",
          7448 => x"1c34810b",
          7449 => x"831c347e",
          7450 => x"51e7bd3f",
          7451 => x"7f54fcc0",
          7452 => x"39861933",
          7453 => x"871a3371",
          7454 => x"8b2b7183",
          7455 => x"2b077905",
          7456 => x"841c3385",
          7457 => x"1d337188",
          7458 => x"2b077088",
          7459 => x"2a5c485e",
          7460 => x"43595576",
          7461 => x"61840534",
          7462 => x"63618505",
          7463 => x"3484b8d4",
          7464 => x"08701e84",
          7465 => x"11338512",
          7466 => x"33718b2b",
          7467 => x"71832b07",
          7468 => x"74058614",
          7469 => x"33871533",
          7470 => x"71882b07",
          7471 => x"70882a41",
          7472 => x"5f484859",
          7473 => x"56594079",
          7474 => x"64860534",
          7475 => x"78648705",
          7476 => x"3484b8d4",
          7477 => x"081d7033",
          7478 => x"81123371",
          7479 => x"882b0781",
          7480 => x"ffff0670",
          7481 => x"882a5942",
          7482 => x"58587578",
          7483 => x"347f8119",
          7484 => x"3484b8d4",
          7485 => x"08701f70",
          7486 => x"33811233",
          7487 => x"718b2b71",
          7488 => x"832b0774",
          7489 => x"05703381",
          7490 => x"12337188",
          7491 => x"2b077083",
          7492 => x"2b8ffff8",
          7493 => x"06770563",
          7494 => x"882a485d",
          7495 => x"5d5a5d40",
          7496 => x"5d44417f",
          7497 => x"8217347b",
          7498 => x"83173484",
          7499 => x"b8d40870",
          7500 => x"1f703381",
          7501 => x"1233718b",
          7502 => x"2b71832b",
          7503 => x"07740570",
          7504 => x"33811233",
          7505 => x"71882b07",
          7506 => x"81ffff06",
          7507 => x"70882a48",
          7508 => x"5d5e5e46",
          7509 => x"5a415b60",
          7510 => x"60347660",
          7511 => x"81053461",
          7512 => x"83ffff06",
          7513 => x"5bfab339",
          7514 => x"86153387",
          7515 => x"1633718b",
          7516 => x"2b71832b",
          7517 => x"07790584",
          7518 => x"18338519",
          7519 => x"3371882b",
          7520 => x"0770882a",
          7521 => x"5e5e5a52",
          7522 => x"415d7884",
          7523 => x"1e347985",
          7524 => x"1e3484b8",
          7525 => x"d4087019",
          7526 => x"84113385",
          7527 => x"1233718b",
          7528 => x"2b71832b",
          7529 => x"07740586",
          7530 => x"14338715",
          7531 => x"3371882b",
          7532 => x"0770882a",
          7533 => x"44565e52",
          7534 => x"5a425556",
          7535 => x"7c608605",
          7536 => x"34756087",
          7537 => x"053484b8",
          7538 => x"d4081870",
          7539 => x"33811233",
          7540 => x"71882b07",
          7541 => x"81ffff06",
          7542 => x"70882a5b",
          7543 => x"5b585577",
          7544 => x"75347881",
          7545 => x"163484b8",
          7546 => x"d408701f",
          7547 => x"70338112",
          7548 => x"33718b2b",
          7549 => x"71832b07",
          7550 => x"74057033",
          7551 => x"81123371",
          7552 => x"882b0770",
          7553 => x"832b8fff",
          7554 => x"f8067705",
          7555 => x"63882a56",
          7556 => x"545f5f58",
          7557 => x"59425e55",
          7558 => x"7f821734",
          7559 => x"7b831734",
          7560 => x"84b8d408",
          7561 => x"701f7033",
          7562 => x"81123371",
          7563 => x"8b2b7183",
          7564 => x"2b077405",
          7565 => x"70338112",
          7566 => x"3371882b",
          7567 => x"0781ffff",
          7568 => x"0670882a",
          7569 => x"5d545e58",
          7570 => x"5b595d55",
          7571 => x"757c3476",
          7572 => x"811d3484",
          7573 => x"b8d40870",
          7574 => x"1f821133",
          7575 => x"83123371",
          7576 => x"8b2b7183",
          7577 => x"2b077411",
          7578 => x"86113387",
          7579 => x"1233718b",
          7580 => x"2b71832b",
          7581 => x"07780584",
          7582 => x"14338515",
          7583 => x"3371882b",
          7584 => x"0770882a",
          7585 => x"59574952",
          7586 => x"5c425953",
          7587 => x"5d5a5757",
          7588 => x"77841d34",
          7589 => x"79851d34",
          7590 => x"84b8d408",
          7591 => x"70178411",
          7592 => x"33851233",
          7593 => x"718b2b71",
          7594 => x"832b0774",
          7595 => x"05861433",
          7596 => x"87153371",
          7597 => x"882b0770",
          7598 => x"882a5f42",
          7599 => x"5e524057",
          7600 => x"41577786",
          7601 => x"16347b87",
          7602 => x"163484b8",
          7603 => x"d4081670",
          7604 => x"33811233",
          7605 => x"71882b07",
          7606 => x"81ffff06",
          7607 => x"70882a5a",
          7608 => x"5c5e5976",
          7609 => x"79347981",
          7610 => x"1a3484b8",
          7611 => x"d408701f",
          7612 => x"82113383",
          7613 => x"1233718b",
          7614 => x"2b71832b",
          7615 => x"07740573",
          7616 => x"33811533",
          7617 => x"71882b07",
          7618 => x"70882a41",
          7619 => x"5c455d5f",
          7620 => x"5a555579",
          7621 => x"79347581",
          7622 => x"1a3484b8",
          7623 => x"d408701f",
          7624 => x"70338112",
          7625 => x"33718b2b",
          7626 => x"71832b07",
          7627 => x"74058214",
          7628 => x"33831533",
          7629 => x"71882b07",
          7630 => x"70882a41",
          7631 => x"5c455d5f",
          7632 => x"5a555579",
          7633 => x"821a3475",
          7634 => x"831a3484",
          7635 => x"b8d40870",
          7636 => x"1f821133",
          7637 => x"83123371",
          7638 => x"882b0766",
          7639 => x"57625670",
          7640 => x"832b4252",
          7641 => x"5a5d7e05",
          7642 => x"840551fe",
          7643 => x"b6d43f84",
          7644 => x"b8d4081e",
          7645 => x"84056165",
          7646 => x"051c7083",
          7647 => x"ffff065d",
          7648 => x"445ff1d5",
          7649 => x"39861933",
          7650 => x"871a3371",
          7651 => x"8b2b7183",
          7652 => x"2b077905",
          7653 => x"841c3385",
          7654 => x"1d337188",
          7655 => x"2b077088",
          7656 => x"2a40485d",
          7657 => x"4341557a",
          7658 => x"61840534",
          7659 => x"63618505",
          7660 => x"3484b8d4",
          7661 => x"08701e84",
          7662 => x"11338512",
          7663 => x"33718b2b",
          7664 => x"71832b07",
          7665 => x"74058614",
          7666 => x"33871533",
          7667 => x"71882b07",
          7668 => x"70882a5b",
          7669 => x"415f485c",
          7670 => x"59415673",
          7671 => x"64860534",
          7672 => x"7a648705",
          7673 => x"3484b8d4",
          7674 => x"081d7033",
          7675 => x"81123371",
          7676 => x"882b0781",
          7677 => x"ffff0670",
          7678 => x"882a5c5f",
          7679 => x"42557875",
          7680 => x"347c8116",
          7681 => x"3484b8d4",
          7682 => x"08701f70",
          7683 => x"33811233",
          7684 => x"718b2b71",
          7685 => x"832b0774",
          7686 => x"05703381",
          7687 => x"12337188",
          7688 => x"2b077083",
          7689 => x"2b8ffff8",
          7690 => x"06770563",
          7691 => x"882a5d44",
          7692 => x"5c49585e",
          7693 => x"45584074",
          7694 => x"821e347b",
          7695 => x"831e3484",
          7696 => x"b8d40870",
          7697 => x"1f703381",
          7698 => x"1233718b",
          7699 => x"2b71832b",
          7700 => x"07740570",
          7701 => x"33811233",
          7702 => x"71882b07",
          7703 => x"81ffff06",
          7704 => x"70882a47",
          7705 => x"5f495846",
          7706 => x"595e5b7f",
          7707 => x"7d347881",
          7708 => x"1e347783",
          7709 => x"ffff065b",
          7710 => x"f383397e",
          7711 => x"605254e5",
          7712 => x"a13f84b8",
          7713 => x"e4085f84",
          7714 => x"b8e40880",
          7715 => x"2e933862",
          7716 => x"53735284",
          7717 => x"b8e40851",
          7718 => x"feb5cf3f",
          7719 => x"7351df88",
          7720 => x"3f615b61",
          7721 => x"7b27efb7",
          7722 => x"38f0e939",
          7723 => x"f93d0d7a",
          7724 => x"7a2984b8",
          7725 => x"d4085858",
          7726 => x"76802eb7",
          7727 => x"38775477",
          7728 => x"8a387384",
          7729 => x"b8e40c89",
          7730 => x"3d0d0477",
          7731 => x"51e4d33f",
          7732 => x"84b8e408",
          7733 => x"5484b8e4",
          7734 => x"08802ee6",
          7735 => x"38775380",
          7736 => x"5284b8e4",
          7737 => x"0851feb7",
          7738 => x"963f7384",
          7739 => x"b8e40c89",
          7740 => x"3d0d0484",
          7741 => x"fff40b84",
          7742 => x"b8d40ca0",
          7743 => x"800b84b8",
          7744 => x"d0238280",
          7745 => x"80537652",
          7746 => x"84fff451",
          7747 => x"feb6f03f",
          7748 => x"84b8d408",
          7749 => x"55767534",
          7750 => x"810b8116",
          7751 => x"3484b8d4",
          7752 => x"08547684",
          7753 => x"1534810b",
          7754 => x"85153484",
          7755 => x"b8d40856",
          7756 => x"76861734",
          7757 => x"810b8717",
          7758 => x"3484b8d4",
          7759 => x"0884b8d0",
          7760 => x"22ff05fe",
          7761 => x"80800770",
          7762 => x"83ffff06",
          7763 => x"70882a58",
          7764 => x"51555674",
          7765 => x"88173473",
          7766 => x"89173484",
          7767 => x"b8d02270",
          7768 => x"10101084",
          7769 => x"b8d40805",
          7770 => x"f8055555",
          7771 => x"76821534",
          7772 => x"810b8315",
          7773 => x"34775477",
          7774 => x"802efec6",
          7775 => x"38fecc39",
          7776 => x"ff3d0d02",
          7777 => x"8f053351",
          7778 => x"81527072",
          7779 => x"26873884",
          7780 => x"b8e01133",
          7781 => x"527184b8",
          7782 => x"e40c833d",
          7783 => x"0d04fe3d",
          7784 => x"0d029305",
          7785 => x"33528353",
          7786 => x"7181269d",
          7787 => x"387151d4",
          7788 => x"bb3f84b8",
          7789 => x"e40881ff",
          7790 => x"06537287",
          7791 => x"387284b8",
          7792 => x"e0133484",
          7793 => x"b8e01233",
          7794 => x"537284b8",
          7795 => x"e40c843d",
          7796 => x"0d04f73d",
          7797 => x"0d7c7e60",
          7798 => x"028c05af",
          7799 => x"05335a5c",
          7800 => x"57598154",
          7801 => x"76742687",
          7802 => x"3884b8e0",
          7803 => x"17335473",
          7804 => x"81065483",
          7805 => x"5573bd38",
          7806 => x"7358850b",
          7807 => x"87c0988c",
          7808 => x"0c785375",
          7809 => x"527651d5",
          7810 => x"ca3f84b8",
          7811 => x"e40881ff",
          7812 => x"06557480",
          7813 => x"2ea73887",
          7814 => x"c0988c08",
          7815 => x"5473e238",
          7816 => x"797826d6",
          7817 => x"3874fc80",
          7818 => x"80065473",
          7819 => x"802e8338",
          7820 => x"81547355",
          7821 => x"7484b8e4",
          7822 => x"0c8b3d0d",
          7823 => x"04848016",
          7824 => x"81197081",
          7825 => x"ff065a55",
          7826 => x"56797826",
          7827 => x"ffac38d5",
          7828 => x"39f73d0d",
          7829 => x"7c7e6002",
          7830 => x"8c05af05",
          7831 => x"335a5c57",
          7832 => x"59815476",
          7833 => x"74268738",
          7834 => x"84b8e017",
          7835 => x"33547381",
          7836 => x"06548355",
          7837 => x"73bd3873",
          7838 => x"58850b87",
          7839 => x"c0988c0c",
          7840 => x"78537552",
          7841 => x"7651d78e",
          7842 => x"3f84b8e4",
          7843 => x"0881ff06",
          7844 => x"5574802e",
          7845 => x"a73887c0",
          7846 => x"988c0854",
          7847 => x"73e23879",
          7848 => x"7826d638",
          7849 => x"74fc8080",
          7850 => x"06547380",
          7851 => x"2e833881",
          7852 => x"54735574",
          7853 => x"84b8e40c",
          7854 => x"8b3d0d04",
          7855 => x"84801681",
          7856 => x"197081ff",
          7857 => x"065a5556",
          7858 => x"797826ff",
          7859 => x"ac38d539",
          7860 => x"fc3d0d78",
          7861 => x"0284059b",
          7862 => x"05330288",
          7863 => x"059f0533",
          7864 => x"53535581",
          7865 => x"53717326",
          7866 => x"873884b8",
          7867 => x"e0123353",
          7868 => x"72810654",
          7869 => x"8353739b",
          7870 => x"38850b87",
          7871 => x"c0988c0c",
          7872 => x"81537073",
          7873 => x"2e963872",
          7874 => x"7125ad38",
          7875 => x"70832e9a",
          7876 => x"38845372",
          7877 => x"84b8e40c",
          7878 => x"863d0d04",
          7879 => x"88800a75",
          7880 => x"0c7384b8",
          7881 => x"e40c863d",
          7882 => x"0d048180",
          7883 => x"750c800b",
          7884 => x"84b8e40c",
          7885 => x"863d0d04",
          7886 => x"71842b87",
          7887 => x"c0928c11",
          7888 => x"535470cd",
          7889 => x"38710870",
          7890 => x"812a8106",
          7891 => x"51517080",
          7892 => x"2e8a3887",
          7893 => x"c0988c08",
          7894 => x"5574ea38",
          7895 => x"87c0988c",
          7896 => x"085170ca",
          7897 => x"3881720c",
          7898 => x"87c0928c",
          7899 => x"14527108",
          7900 => x"82065473",
          7901 => x"802eff9b",
          7902 => x"38710882",
          7903 => x"065473ee",
          7904 => x"38ff9039",
          7905 => x"f63d0d7c",
          7906 => x"58800b83",
          7907 => x"1933715b",
          7908 => x"56577477",
          7909 => x"2e098106",
          7910 => x"a8387733",
          7911 => x"5675832e",
          7912 => x"81873880",
          7913 => x"53805281",
          7914 => x"183351fe",
          7915 => x"a33f84b8",
          7916 => x"e408802e",
          7917 => x"83388159",
          7918 => x"7884b8e4",
          7919 => x"0c8c3d0d",
          7920 => x"048154b4",
          7921 => x"180853b8",
          7922 => x"18705381",
          7923 => x"1933525a",
          7924 => x"fcff3f81",
          7925 => x"5984b8e4",
          7926 => x"08772e09",
          7927 => x"8106d938",
          7928 => x"84b8e408",
          7929 => x"831934b4",
          7930 => x"180870a8",
          7931 => x"1a0831a0",
          7932 => x"1a0884b8",
          7933 => x"e4085c58",
          7934 => x"565b7476",
          7935 => x"27ff9b38",
          7936 => x"82183355",
          7937 => x"74822e09",
          7938 => x"8106ff8e",
          7939 => x"38815475",
          7940 => x"1b537952",
          7941 => x"81183351",
          7942 => x"fcb73f76",
          7943 => x"78335759",
          7944 => x"75832e09",
          7945 => x"8106fefb",
          7946 => x"38841833",
          7947 => x"5776812e",
          7948 => x"098106fe",
          7949 => x"ee38b818",
          7950 => x"5a84807a",
          7951 => x"56578075",
          7952 => x"70810557",
          7953 => x"34ff1757",
          7954 => x"76f43880",
          7955 => x"d50b84b6",
          7956 => x"1934ffaa",
          7957 => x"0b84b719",
          7958 => x"3480d27a",
          7959 => x"3480d20b",
          7960 => x"b9193480",
          7961 => x"e10bba19",
          7962 => x"3480c10b",
          7963 => x"bb193480",
          7964 => x"f20b849c",
          7965 => x"193480f2",
          7966 => x"0b849d19",
          7967 => x"3480c10b",
          7968 => x"849e1934",
          7969 => x"80e10b84",
          7970 => x"9f193494",
          7971 => x"18085574",
          7972 => x"84a01934",
          7973 => x"74882a5b",
          7974 => x"7a84a119",
          7975 => x"3474902a",
          7976 => x"567584a2",
          7977 => x"19347498",
          7978 => x"2a5b7a84",
          7979 => x"a3193490",
          7980 => x"18085b7a",
          7981 => x"84a41934",
          7982 => x"7a882a55",
          7983 => x"7484a519",
          7984 => x"347a902a",
          7985 => x"567584a6",
          7986 => x"19347a98",
          7987 => x"2a557484",
          7988 => x"a71934a4",
          7989 => x"18088105",
          7990 => x"70b41a0c",
          7991 => x"5b81547a",
          7992 => x"53795281",
          7993 => x"183351fa",
          7994 => x"e83f7684",
          7995 => x"19348053",
          7996 => x"80528118",
          7997 => x"3351fbd8",
          7998 => x"3f84b8e4",
          7999 => x"08802efd",
          8000 => x"b738fdb2",
          8001 => x"39f33d0d",
          8002 => x"60607008",
          8003 => x"59565681",
          8004 => x"76278838",
          8005 => x"9c170876",
          8006 => x"268c3881",
          8007 => x"587784b8",
          8008 => x"e40c8f3d",
          8009 => x"0d04ff77",
          8010 => x"33565874",
          8011 => x"822e81cc",
          8012 => x"38748224",
          8013 => x"82a53874",
          8014 => x"812e0981",
          8015 => x"06dd3875",
          8016 => x"812a1670",
          8017 => x"892aa819",
          8018 => x"08055a5a",
          8019 => x"805bb417",
          8020 => x"08792eb0",
          8021 => x"38831733",
          8022 => x"5c7b7b2e",
          8023 => x"09810683",
          8024 => x"de388154",
          8025 => x"7853b817",
          8026 => x"52811733",
          8027 => x"51f8e33f",
          8028 => x"84b8e408",
          8029 => x"802e8538",
          8030 => x"ff59815b",
          8031 => x"78b4180c",
          8032 => x"7aff9a38",
          8033 => x"7983ff06",
          8034 => x"17b81133",
          8035 => x"811c7089",
          8036 => x"2aa81b08",
          8037 => x"05535d5d",
          8038 => x"59b41708",
          8039 => x"792eb538",
          8040 => x"800b8318",
          8041 => x"33715c56",
          8042 => x"5d747d2e",
          8043 => x"09810684",
          8044 => x"b5388154",
          8045 => x"7853b817",
          8046 => x"52811733",
          8047 => x"51f8933f",
          8048 => x"84b8e408",
          8049 => x"802e8538",
          8050 => x"ff59815a",
          8051 => x"78b4180c",
          8052 => x"79feca38",
          8053 => x"7a83ff06",
          8054 => x"17b81133",
          8055 => x"70882b7e",
          8056 => x"07788106",
          8057 => x"71842a53",
          8058 => x"5d59595d",
          8059 => x"79feae38",
          8060 => x"769fff06",
          8061 => x"84b8e40c",
          8062 => x"8f3d0d04",
          8063 => x"75882aa8",
          8064 => x"18080559",
          8065 => x"b4170879",
          8066 => x"2eb53880",
          8067 => x"0b831833",
          8068 => x"715c5d5b",
          8069 => x"7b7b2e09",
          8070 => x"810681c2",
          8071 => x"38815478",
          8072 => x"53b81752",
          8073 => x"81173351",
          8074 => x"f7a83f84",
          8075 => x"b8e40880",
          8076 => x"2e8538ff",
          8077 => x"59815a78",
          8078 => x"b4180c79",
          8079 => x"fddf3875",
          8080 => x"1083fe06",
          8081 => x"7705b805",
          8082 => x"81113371",
          8083 => x"3371882b",
          8084 => x"0784b8e4",
          8085 => x"0c575b8f",
          8086 => x"3d0d0474",
          8087 => x"832e0981",
          8088 => x"06fdb838",
          8089 => x"75872aa8",
          8090 => x"18080559",
          8091 => x"b4170879",
          8092 => x"2eb53880",
          8093 => x"0b831833",
          8094 => x"715c5e5b",
          8095 => x"7c7b2e09",
          8096 => x"81068281",
          8097 => x"38815478",
          8098 => x"53b81752",
          8099 => x"81173351",
          8100 => x"f6c03f84",
          8101 => x"b8e40880",
          8102 => x"2e8538ff",
          8103 => x"59815a78",
          8104 => x"b4180c79",
          8105 => x"fcf73875",
          8106 => x"822b83fc",
          8107 => x"067705b8",
          8108 => x"05831133",
          8109 => x"82123371",
          8110 => x"902b7188",
          8111 => x"2b078114",
          8112 => x"33707207",
          8113 => x"882b7533",
          8114 => x"7180ffff",
          8115 => x"fe800607",
          8116 => x"84b8e40c",
          8117 => x"415c5e59",
          8118 => x"5a568f3d",
          8119 => x"0d048154",
          8120 => x"b4170853",
          8121 => x"b8177053",
          8122 => x"81183352",
          8123 => x"5cf6e23f",
          8124 => x"815a84b8",
          8125 => x"e4087b2e",
          8126 => x"098106fe",
          8127 => x"be3884b8",
          8128 => x"e4088318",
          8129 => x"34b41708",
          8130 => x"a8180831",
          8131 => x"84b8e408",
          8132 => x"5b5e7da0",
          8133 => x"180827fe",
          8134 => x"84388217",
          8135 => x"33557482",
          8136 => x"2e098106",
          8137 => x"fdf73881",
          8138 => x"54b41708",
          8139 => x"a0180805",
          8140 => x"537b5281",
          8141 => x"173351f6",
          8142 => x"983f7a5a",
          8143 => x"fddf3981",
          8144 => x"54b41708",
          8145 => x"53b81770",
          8146 => x"53811833",
          8147 => x"525cf681",
          8148 => x"3f84b8e4",
          8149 => x"087b2e09",
          8150 => x"81068281",
          8151 => x"3884b8e4",
          8152 => x"08831834",
          8153 => x"b41708a8",
          8154 => x"1808315d",
          8155 => x"7ca01808",
          8156 => x"278b3882",
          8157 => x"17335e7d",
          8158 => x"822e81cb",
          8159 => x"3884b8e4",
          8160 => x"085bfbde",
          8161 => x"398154b4",
          8162 => x"170853b8",
          8163 => x"17705381",
          8164 => x"1833525c",
          8165 => x"f5bb3f81",
          8166 => x"5a84b8e4",
          8167 => x"087b2e09",
          8168 => x"8106fdff",
          8169 => x"3884b8e4",
          8170 => x"08831834",
          8171 => x"b41708a8",
          8172 => x"18083184",
          8173 => x"b8e4085b",
          8174 => x"5e7da018",
          8175 => x"0827fdc5",
          8176 => x"38821733",
          8177 => x"5574822e",
          8178 => x"098106fd",
          8179 => x"b8388154",
          8180 => x"b41708a0",
          8181 => x"18080553",
          8182 => x"7b528117",
          8183 => x"3351f4f1",
          8184 => x"3f7a5afd",
          8185 => x"a0398154",
          8186 => x"b4170853",
          8187 => x"b8177053",
          8188 => x"81183352",
          8189 => x"5ef4da3f",
          8190 => x"815a84b8",
          8191 => x"e4087d2e",
          8192 => x"098106fb",
          8193 => x"cb3884b8",
          8194 => x"e4088318",
          8195 => x"34b41708",
          8196 => x"a8180831",
          8197 => x"84b8e408",
          8198 => x"5b5574a0",
          8199 => x"180827fb",
          8200 => x"91388217",
          8201 => x"33557482",
          8202 => x"2e098106",
          8203 => x"fb843881",
          8204 => x"54b41708",
          8205 => x"a0180805",
          8206 => x"537d5281",
          8207 => x"173351f4",
          8208 => x"903f7c5a",
          8209 => x"faec3981",
          8210 => x"54b41708",
          8211 => x"a0180805",
          8212 => x"537b5281",
          8213 => x"173351f3",
          8214 => x"f83ffa86",
          8215 => x"39815b7a",
          8216 => x"f9bb38fa",
          8217 => x"9f39f23d",
          8218 => x"0d606264",
          8219 => x"5d575982",
          8220 => x"58817627",
          8221 => x"9c38759c",
          8222 => x"1a082795",
          8223 => x"38783355",
          8224 => x"74782e96",
          8225 => x"38747824",
          8226 => x"81803874",
          8227 => x"812e828a",
          8228 => x"387784b8",
          8229 => x"e40c903d",
          8230 => x"0d047588",
          8231 => x"2aa81a08",
          8232 => x"0558800b",
          8233 => x"b41a0858",
          8234 => x"5c76782e",
          8235 => x"86b63883",
          8236 => x"19337c5b",
          8237 => x"5d7c7c2e",
          8238 => x"09810683",
          8239 => x"fa388154",
          8240 => x"7753b819",
          8241 => x"52811933",
          8242 => x"51f2873f",
          8243 => x"84b8e408",
          8244 => x"802e8538",
          8245 => x"ff58815a",
          8246 => x"77b41a0c",
          8247 => x"795879ff",
          8248 => x"b0387510",
          8249 => x"83fe0679",
          8250 => x"057b83ff",
          8251 => x"ff06585e",
          8252 => x"76b81f34",
          8253 => x"76882a5a",
          8254 => x"79b91f34",
          8255 => x"810b831a",
          8256 => x"347784b8",
          8257 => x"e40c903d",
          8258 => x"0d047483",
          8259 => x"2e098106",
          8260 => x"feff3875",
          8261 => x"872aa81a",
          8262 => x"08055880",
          8263 => x"0bb41a08",
          8264 => x"585c7678",
          8265 => x"2e85e138",
          8266 => x"8319337c",
          8267 => x"5b5d7c7c",
          8268 => x"2e098106",
          8269 => x"84bd3881",
          8270 => x"547753b8",
          8271 => x"19528119",
          8272 => x"3351f18e",
          8273 => x"3f84b8e4",
          8274 => x"08802e85",
          8275 => x"38ff5881",
          8276 => x"5a77b41a",
          8277 => x"0c795879",
          8278 => x"feb73875",
          8279 => x"822b83fc",
          8280 => x"067905b8",
          8281 => x"11831133",
          8282 => x"70982b8f",
          8283 => x"0a067ef0",
          8284 => x"0a060741",
          8285 => x"575e5c7d",
          8286 => x"7d347d88",
          8287 => x"2a5675b9",
          8288 => x"1d347d90",
          8289 => x"2a5a79ba",
          8290 => x"1d347d98",
          8291 => x"2a5b7abb",
          8292 => x"1d34810b",
          8293 => x"831a34fe",
          8294 => x"e8397581",
          8295 => x"2a167089",
          8296 => x"2aa81b08",
          8297 => x"05b41b08",
          8298 => x"59595a76",
          8299 => x"782eb738",
          8300 => x"800b831a",
          8301 => x"33715e56",
          8302 => x"5d747d2e",
          8303 => x"09810682",
          8304 => x"d4388154",
          8305 => x"7753b819",
          8306 => x"52811933",
          8307 => x"51f0833f",
          8308 => x"84b8e408",
          8309 => x"802e8538",
          8310 => x"ff58815c",
          8311 => x"77b41a0c",
          8312 => x"7b587bfd",
          8313 => x"ac387983",
          8314 => x"ff0619b8",
          8315 => x"05811b77",
          8316 => x"81065f5f",
          8317 => x"577a557c",
          8318 => x"802e8f38",
          8319 => x"7a842b9f",
          8320 => x"f0067733",
          8321 => x"8f067107",
          8322 => x"565a7477",
          8323 => x"34810b83",
          8324 => x"1a347d89",
          8325 => x"2aa81a08",
          8326 => x"0556800b",
          8327 => x"b41a0856",
          8328 => x"5f74762e",
          8329 => x"83dd3881",
          8330 => x"547453b8",
          8331 => x"19705381",
          8332 => x"1a335257",
          8333 => x"f09b3f81",
          8334 => x"5884b8e4",
          8335 => x"087f2e09",
          8336 => x"810680c7",
          8337 => x"3884b8e4",
          8338 => x"08831a34",
          8339 => x"b4190870",
          8340 => x"a81b0831",
          8341 => x"a01b0884",
          8342 => x"b8e4085b",
          8343 => x"5c565c74",
          8344 => x"7a278b38",
          8345 => x"82193355",
          8346 => x"74822e82",
          8347 => x"e4388154",
          8348 => x"75537652",
          8349 => x"81193351",
          8350 => x"eed83f84",
          8351 => x"b8e40880",
          8352 => x"2e8538ff",
          8353 => x"56815875",
          8354 => x"b41a0c77",
          8355 => x"fc83387d",
          8356 => x"83ff0619",
          8357 => x"b8057b84",
          8358 => x"2a56567c",
          8359 => x"8f387a88",
          8360 => x"2a763381",
          8361 => x"f006718f",
          8362 => x"0607565c",
          8363 => x"74763481",
          8364 => x"0b831a34",
          8365 => x"fccb3981",
          8366 => x"547653b8",
          8367 => x"19705381",
          8368 => x"1a33525d",
          8369 => x"ef8b3f81",
          8370 => x"5a84b8e4",
          8371 => x"087c2e09",
          8372 => x"8106fc88",
          8373 => x"3884b8e4",
          8374 => x"08831a34",
          8375 => x"b4190870",
          8376 => x"a81b0831",
          8377 => x"a01b0884",
          8378 => x"b8e4085d",
          8379 => x"59405e7e",
          8380 => x"7727fbca",
          8381 => x"38821933",
          8382 => x"5574822e",
          8383 => x"098106fb",
          8384 => x"bd388154",
          8385 => x"761e537c",
          8386 => x"52811933",
          8387 => x"51eec23f",
          8388 => x"7b5afbaa",
          8389 => x"39815476",
          8390 => x"53b81970",
          8391 => x"53811a33",
          8392 => x"5257eead",
          8393 => x"3f815c84",
          8394 => x"b8e4087d",
          8395 => x"2e098106",
          8396 => x"fdae3884",
          8397 => x"b8e40883",
          8398 => x"1a34b419",
          8399 => x"0870a81b",
          8400 => x"0831a01b",
          8401 => x"0884b8e4",
          8402 => x"085f4056",
          8403 => x"5f747e27",
          8404 => x"fcf03882",
          8405 => x"19335574",
          8406 => x"822e0981",
          8407 => x"06fce338",
          8408 => x"81547d1f",
          8409 => x"53765281",
          8410 => x"193351ed",
          8411 => x"e43f7c5c",
          8412 => x"fcd03981",
          8413 => x"547653b8",
          8414 => x"19705381",
          8415 => x"1a335257",
          8416 => x"edcf3f81",
          8417 => x"5a84b8e4",
          8418 => x"087c2e09",
          8419 => x"8106fbc5",
          8420 => x"3884b8e4",
          8421 => x"08831a34",
          8422 => x"b4190870",
          8423 => x"a81b0831",
          8424 => x"a01b0884",
          8425 => x"b8e4085d",
          8426 => x"5f405e7e",
          8427 => x"7d27fb87",
          8428 => x"38821933",
          8429 => x"5574822e",
          8430 => x"098106fa",
          8431 => x"fa388154",
          8432 => x"7c1e5376",
          8433 => x"52811933",
          8434 => x"51ed863f",
          8435 => x"7b5afae7",
          8436 => x"39815479",
          8437 => x"1c537652",
          8438 => x"81193351",
          8439 => x"ecf33f7e",
          8440 => x"58fd8b39",
          8441 => x"7b761083",
          8442 => x"fe067a05",
          8443 => x"7c83ffff",
          8444 => x"06595f58",
          8445 => x"76b81f34",
          8446 => x"76882a5a",
          8447 => x"79b91f34",
          8448 => x"f9fa397e",
          8449 => x"58fd8839",
          8450 => x"7b76822b",
          8451 => x"83fc067a",
          8452 => x"05b81183",
          8453 => x"11337098",
          8454 => x"2b8f0a06",
          8455 => x"7ff00a06",
          8456 => x"0742585f",
          8457 => x"5d587d7d",
          8458 => x"347d882a",
          8459 => x"5675b91d",
          8460 => x"347d902a",
          8461 => x"5a79ba1d",
          8462 => x"347d982a",
          8463 => x"5b7abb1d",
          8464 => x"34facf39",
          8465 => x"f63d0d7c",
          8466 => x"7e71085b",
          8467 => x"5c5a7a81",
          8468 => x"8a389019",
          8469 => x"08577680",
          8470 => x"2e80f438",
          8471 => x"769c1a08",
          8472 => x"2780ec38",
          8473 => x"94190870",
          8474 => x"56547380",
          8475 => x"2e80d738",
          8476 => x"767b2e81",
          8477 => x"93387656",
          8478 => x"8116569c",
          8479 => x"19087626",
          8480 => x"89388256",
          8481 => x"75772682",
          8482 => x"b2387552",
          8483 => x"7951f0f5",
          8484 => x"3f84b8e4",
          8485 => x"08802e81",
          8486 => x"d0388058",
          8487 => x"84b8e408",
          8488 => x"812eb138",
          8489 => x"84b8e408",
          8490 => x"09703070",
          8491 => x"72078025",
          8492 => x"707b0751",
          8493 => x"51555573",
          8494 => x"82aa3875",
          8495 => x"772e0981",
          8496 => x"06ffb538",
          8497 => x"73557484",
          8498 => x"b8e40c8c",
          8499 => x"3d0d0481",
          8500 => x"57ff9139",
          8501 => x"84b8e408",
          8502 => x"58ca397a",
          8503 => x"527951f0",
          8504 => x"a43f8155",
          8505 => x"7484b8e4",
          8506 => x"0827db38",
          8507 => x"84b8e408",
          8508 => x"5584b8e4",
          8509 => x"08ff2ece",
          8510 => x"389c1908",
          8511 => x"84b8e408",
          8512 => x"26c4387a",
          8513 => x"57fedd39",
          8514 => x"811b569c",
          8515 => x"19087626",
          8516 => x"83388256",
          8517 => x"75527951",
          8518 => x"efeb3f80",
          8519 => x"5884b8e4",
          8520 => x"08812e81",
          8521 => x"a03884b8",
          8522 => x"e4080970",
          8523 => x"30707207",
          8524 => x"8025707b",
          8525 => x"0784b8e4",
          8526 => x"08545151",
          8527 => x"555573ff",
          8528 => x"853884b8",
          8529 => x"e408802e",
          8530 => x"9a389019",
          8531 => x"08548174",
          8532 => x"27fea338",
          8533 => x"739c1a08",
          8534 => x"27fe9b38",
          8535 => x"73705757",
          8536 => x"fe963975",
          8537 => x"802efe8e",
          8538 => x"38ff5375",
          8539 => x"527851f5",
          8540 => x"f53f84b8",
          8541 => x"e40884b8",
          8542 => x"e4083070",
          8543 => x"84b8e408",
          8544 => x"07802556",
          8545 => x"58557a80",
          8546 => x"c4387480",
          8547 => x"e3387590",
          8548 => x"1a0c9c19",
          8549 => x"08fe0594",
          8550 => x"1a085658",
          8551 => x"74782686",
          8552 => x"38ff1594",
          8553 => x"1a0c8419",
          8554 => x"3381075a",
          8555 => x"79841a34",
          8556 => x"75557484",
          8557 => x"b8e40c8c",
          8558 => x"3d0d0480",
          8559 => x"0b84b8e4",
          8560 => x"0c8c3d0d",
          8561 => x"0484b8e4",
          8562 => x"0858feda",
          8563 => x"3973802e",
          8564 => x"ffb83875",
          8565 => x"537a5278",
          8566 => x"51f58b3f",
          8567 => x"84b8e408",
          8568 => x"55ffa739",
          8569 => x"84b8e408",
          8570 => x"84b8e40c",
          8571 => x"8c3d0d04",
          8572 => x"ff567481",
          8573 => x"2effb938",
          8574 => x"8155ffb6",
          8575 => x"39f83d0d",
          8576 => x"7a7c7108",
          8577 => x"59555873",
          8578 => x"f0800a26",
          8579 => x"80df3873",
          8580 => x"9f065372",
          8581 => x"80d73873",
          8582 => x"90190c88",
          8583 => x"18085574",
          8584 => x"80df3876",
          8585 => x"33567582",
          8586 => x"2680cc38",
          8587 => x"73852a53",
          8588 => x"820b8818",
          8589 => x"225a5672",
          8590 => x"7927a938",
          8591 => x"ac170898",
          8592 => x"190c7494",
          8593 => x"190c9818",
          8594 => x"08538256",
          8595 => x"72802e94",
          8596 => x"3873892a",
          8597 => x"1398190c",
          8598 => x"7383ff06",
          8599 => x"17b8059c",
          8600 => x"190c8056",
          8601 => x"7584b8e4",
          8602 => x"0c8a3d0d",
          8603 => x"04820b84",
          8604 => x"b8e40c8a",
          8605 => x"3d0d04ac",
          8606 => x"17085574",
          8607 => x"802effac",
          8608 => x"388a1722",
          8609 => x"70892b57",
          8610 => x"59737627",
          8611 => x"a5389c17",
          8612 => x"0853fe15",
          8613 => x"fe145456",
          8614 => x"80597573",
          8615 => x"278d388a",
          8616 => x"17227671",
          8617 => x"29b01908",
          8618 => x"055a5378",
          8619 => x"98190cff",
          8620 => x"91397452",
          8621 => x"7751eccd",
          8622 => x"3f84b8e4",
          8623 => x"085584b8",
          8624 => x"e408ff2e",
          8625 => x"a438810b",
          8626 => x"84b8e408",
          8627 => x"27ff9e38",
          8628 => x"9c170853",
          8629 => x"84b8e408",
          8630 => x"7327ff91",
          8631 => x"38737631",
          8632 => x"54737627",
          8633 => x"cd38ffaa",
          8634 => x"39810b84",
          8635 => x"b8e40c8a",
          8636 => x"3d0d04f3",
          8637 => x"3d0d7f70",
          8638 => x"08901208",
          8639 => x"a0055c5a",
          8640 => x"57f0800a",
          8641 => x"7a278638",
          8642 => x"800b9818",
          8643 => x"0c981708",
          8644 => x"55845674",
          8645 => x"802eb238",
          8646 => x"7983ff06",
          8647 => x"5b7a9d38",
          8648 => x"81159418",
          8649 => x"08575875",
          8650 => x"a9387985",
          8651 => x"2a881a22",
          8652 => x"57557476",
          8653 => x"2781f538",
          8654 => x"7798180c",
          8655 => x"7990180c",
          8656 => x"781bb805",
          8657 => x"9c180c80",
          8658 => x"567584b8",
          8659 => x"e40c8f3d",
          8660 => x"0d047798",
          8661 => x"180c8a19",
          8662 => x"22ff057a",
          8663 => x"892a065c",
          8664 => x"7bda3875",
          8665 => x"527651eb",
          8666 => x"9c3f84b8",
          8667 => x"e4085d82",
          8668 => x"56810b84",
          8669 => x"b8e40827",
          8670 => x"d0388156",
          8671 => x"84b8e408",
          8672 => x"ff2ec638",
          8673 => x"9c190884",
          8674 => x"b8e40826",
          8675 => x"82913860",
          8676 => x"802e8198",
          8677 => x"38941708",
          8678 => x"527651f9",
          8679 => x"a73f84b8",
          8680 => x"e4085d87",
          8681 => x"5684b8e4",
          8682 => x"08802eff",
          8683 => x"9c388256",
          8684 => x"84b8e408",
          8685 => x"812eff91",
          8686 => x"38815684",
          8687 => x"b8e408ff",
          8688 => x"2eff8638",
          8689 => x"84b8e408",
          8690 => x"831a335f",
          8691 => x"587d80ea",
          8692 => x"38fe189c",
          8693 => x"1a08fe05",
          8694 => x"5956805c",
          8695 => x"7578278d",
          8696 => x"388a1922",
          8697 => x"767129b0",
          8698 => x"1b08055d",
          8699 => x"5e7bb41a",
          8700 => x"0cb81958",
          8701 => x"84807857",
          8702 => x"55807670",
          8703 => x"81055834",
          8704 => x"ff155574",
          8705 => x"f4387456",
          8706 => x"8a192255",
          8707 => x"75752781",
          8708 => x"80388154",
          8709 => x"751c5377",
          8710 => x"52811933",
          8711 => x"51e4b23f",
          8712 => x"84b8e408",
          8713 => x"80e73881",
          8714 => x"1656dd39",
          8715 => x"7a98180c",
          8716 => x"840b84b8",
          8717 => x"e40c8f3d",
          8718 => x"0d047554",
          8719 => x"b4190853",
          8720 => x"b8197053",
          8721 => x"811a3352",
          8722 => x"56e4863f",
          8723 => x"84b8e408",
          8724 => x"80f33884",
          8725 => x"b8e40883",
          8726 => x"1a34b419",
          8727 => x"08a81a08",
          8728 => x"315574a0",
          8729 => x"1a0827fe",
          8730 => x"e8388219",
          8731 => x"335c7b82",
          8732 => x"2e098106",
          8733 => x"fedb3881",
          8734 => x"54b41908",
          8735 => x"a01a0805",
          8736 => x"53755281",
          8737 => x"193351e3",
          8738 => x"c83ffec5",
          8739 => x"398a1922",
          8740 => x"557483ff",
          8741 => x"ff065574",
          8742 => x"762e0981",
          8743 => x"06a7387c",
          8744 => x"94180cfe",
          8745 => x"1d9c1a08",
          8746 => x"fe055e56",
          8747 => x"8058757d",
          8748 => x"27fd8538",
          8749 => x"8a192276",
          8750 => x"7129b01b",
          8751 => x"08059819",
          8752 => x"0c5cfcf8",
          8753 => x"39810b84",
          8754 => x"b8e40c8f",
          8755 => x"3d0d04ee",
          8756 => x"3d0d6466",
          8757 => x"415c847c",
          8758 => x"085a5b81",
          8759 => x"ff70981e",
          8760 => x"08585e5e",
          8761 => x"75802e82",
          8762 => x"d238b819",
          8763 => x"5f755a80",
          8764 => x"58b41908",
          8765 => x"762e82d1",
          8766 => x"38831933",
          8767 => x"78585574",
          8768 => x"782e0981",
          8769 => x"06819438",
          8770 => x"81547553",
          8771 => x"b8195281",
          8772 => x"193351e1",
          8773 => x"bd3f84b8",
          8774 => x"e408802e",
          8775 => x"8538ff5a",
          8776 => x"815779b4",
          8777 => x"1a0c765b",
          8778 => x"76829038",
          8779 => x"9c1c0870",
          8780 => x"33585876",
          8781 => x"802e8281",
          8782 => x"388b1833",
          8783 => x"bf067081",
          8784 => x"ff065b41",
          8785 => x"60861d34",
          8786 => x"7681e532",
          8787 => x"703078ae",
          8788 => x"32703072",
          8789 => x"80257180",
          8790 => x"25075445",
          8791 => x"45575574",
          8792 => x"9338747a",
          8793 => x"df064356",
          8794 => x"61882e81",
          8795 => x"bf387560",
          8796 => x"2e818638",
          8797 => x"81ff5d80",
          8798 => x"527b51fa",
          8799 => x"f63f84b8",
          8800 => x"e4085b84",
          8801 => x"b8e40881",
          8802 => x"b238981c",
          8803 => x"085675fe",
          8804 => x"dc387a84",
          8805 => x"b8e40c94",
          8806 => x"3d0d0481",
          8807 => x"54b41908",
          8808 => x"537e5281",
          8809 => x"193351e1",
          8810 => x"a83f8157",
          8811 => x"84b8e408",
          8812 => x"782e0981",
          8813 => x"06feef38",
          8814 => x"84b8e408",
          8815 => x"831a34b4",
          8816 => x"1908a81a",
          8817 => x"083184b8",
          8818 => x"e408585b",
          8819 => x"7aa01a08",
          8820 => x"27feb538",
          8821 => x"82193341",
          8822 => x"60822e09",
          8823 => x"8106fea8",
          8824 => x"388154b4",
          8825 => x"1908a01a",
          8826 => x"0805537e",
          8827 => x"52811933",
          8828 => x"51e0de3f",
          8829 => x"7757fe90",
          8830 => x"39798f2e",
          8831 => x"09810681",
          8832 => x"e7387686",
          8833 => x"2a81065b",
          8834 => x"7a802e93",
          8835 => x"388d1833",
          8836 => x"7781bf06",
          8837 => x"70901f08",
          8838 => x"7fac050c",
          8839 => x"595e5e76",
          8840 => x"7d2eab38",
          8841 => x"81ff5574",
          8842 => x"5dfecc39",
          8843 => x"81567560",
          8844 => x"2e098106",
          8845 => x"febe38c1",
          8846 => x"39845b80",
          8847 => x"0b981d0c",
          8848 => x"7a84b8e4",
          8849 => x"0c943d0d",
          8850 => x"04775bfd",
          8851 => x"df398d18",
          8852 => x"33577d77",
          8853 => x"2e098106",
          8854 => x"cb388c19",
          8855 => x"089b1933",
          8856 => x"9a1a3371",
          8857 => x"882b0758",
          8858 => x"564175ff",
          8859 => x"b7387733",
          8860 => x"7081bf06",
          8861 => x"8d29f305",
          8862 => x"515a8176",
          8863 => x"585b83e4",
          8864 => x"e4173378",
          8865 => x"05811133",
          8866 => x"71337188",
          8867 => x"2b075244",
          8868 => x"567a802e",
          8869 => x"80c53879",
          8870 => x"81fe26ff",
          8871 => x"87387910",
          8872 => x"6105765c",
          8873 => x"42756223",
          8874 => x"811a5a81",
          8875 => x"17578c77",
          8876 => x"27cc3877",
          8877 => x"3370862a",
          8878 => x"81065957",
          8879 => x"77802e90",
          8880 => x"387981fe",
          8881 => x"26fedd38",
          8882 => x"79106105",
          8883 => x"43806323",
          8884 => x"ff1d7081",
          8885 => x"ff065e41",
          8886 => x"fd9d3975",
          8887 => x"83ffff2e",
          8888 => x"ca3881ff",
          8889 => x"55fec039",
          8890 => x"7ca8387c",
          8891 => x"558b5774",
          8892 => x"812a7581",
          8893 => x"80290578",
          8894 => x"7081055a",
          8895 => x"33407f05",
          8896 => x"7081ff06",
          8897 => x"ff195956",
          8898 => x"5976e438",
          8899 => x"747e2efd",
          8900 => x"8138ff0b",
          8901 => x"ac1d0c7a",
          8902 => x"84b8e40c",
          8903 => x"943d0d04",
          8904 => x"ef3d0d63",
          8905 => x"70085c5c",
          8906 => x"80527b51",
          8907 => x"f5cf3f84",
          8908 => x"b8e4085a",
          8909 => x"84b8e408",
          8910 => x"82803881",
          8911 => x"ff70405d",
          8912 => x"ff0bac1d",
          8913 => x"0cb81b5e",
          8914 => x"981c0856",
          8915 => x"8058b41b",
          8916 => x"08762e82",
          8917 => x"cc38831b",
          8918 => x"33785855",
          8919 => x"74782e09",
          8920 => x"810681df",
          8921 => x"38815475",
          8922 => x"53b81b52",
          8923 => x"811b3351",
          8924 => x"dce03f84",
          8925 => x"b8e40880",
          8926 => x"2e8538ff",
          8927 => x"56815775",
          8928 => x"b41c0c76",
          8929 => x"5a7681b2",
          8930 => x"389c1c08",
          8931 => x"70335859",
          8932 => x"76802e84",
          8933 => x"99388b19",
          8934 => x"33bf0670",
          8935 => x"81ff0657",
          8936 => x"5877861d",
          8937 => x"347681e5",
          8938 => x"2e80f238",
          8939 => x"75832a81",
          8940 => x"0655758f",
          8941 => x"2e81ef38",
          8942 => x"7480e238",
          8943 => x"758f2e81",
          8944 => x"e5387caa",
          8945 => x"38787d56",
          8946 => x"588b5774",
          8947 => x"812a7581",
          8948 => x"80290578",
          8949 => x"7081055a",
          8950 => x"33577605",
          8951 => x"7081ff06",
          8952 => x"ff195956",
          8953 => x"5d76e438",
          8954 => x"747f2e80",
          8955 => x"cd38ab1c",
          8956 => x"33810657",
          8957 => x"76a7388b",
          8958 => x"0ba01d59",
          8959 => x"57787081",
          8960 => x"055a3378",
          8961 => x"7081055a",
          8962 => x"33717131",
          8963 => x"ff1a5a58",
          8964 => x"42407680",
          8965 => x"2e81dc38",
          8966 => x"75802ee1",
          8967 => x"3881ff5d",
          8968 => x"ff0bac1d",
          8969 => x"0c80527b",
          8970 => x"51f5c83f",
          8971 => x"84b8e408",
          8972 => x"5a84b8e4",
          8973 => x"08802efe",
          8974 => x"8f387984",
          8975 => x"b8e40c93",
          8976 => x"3d0d0481",
          8977 => x"54b41b08",
          8978 => x"537d5281",
          8979 => x"1b3351dc",
          8980 => x"803f8157",
          8981 => x"84b8e408",
          8982 => x"782e0981",
          8983 => x"06fea438",
          8984 => x"84b8e408",
          8985 => x"831c34b4",
          8986 => x"1b08a81c",
          8987 => x"083184b8",
          8988 => x"e4085859",
          8989 => x"78a01c08",
          8990 => x"27fdea38",
          8991 => x"821b335a",
          8992 => x"79822e09",
          8993 => x"8106fddd",
          8994 => x"388154b4",
          8995 => x"1b08a01c",
          8996 => x"0805537d",
          8997 => x"52811b33",
          8998 => x"51dbb63f",
          8999 => x"7757fdc5",
          9000 => x"39775afd",
          9001 => x"e439ab1c",
          9002 => x"3370862a",
          9003 => x"81064255",
          9004 => x"60fef238",
          9005 => x"76862a81",
          9006 => x"065a7980",
          9007 => x"2e93388d",
          9008 => x"19337781",
          9009 => x"bf067090",
          9010 => x"1f087fac",
          9011 => x"050c595e",
          9012 => x"5f767d2e",
          9013 => x"af3881ff",
          9014 => x"55745d80",
          9015 => x"527b51f4",
          9016 => x"923f84b8",
          9017 => x"e4085a84",
          9018 => x"b8e40880",
          9019 => x"2efcd938",
          9020 => x"fec83975",
          9021 => x"802efec2",
          9022 => x"3881ff5d",
          9023 => x"ff0bac1d",
          9024 => x"0cfea239",
          9025 => x"8d193357",
          9026 => x"7e772e09",
          9027 => x"8106c738",
          9028 => x"8c1b089b",
          9029 => x"1a339a1b",
          9030 => x"3371882b",
          9031 => x"07594240",
          9032 => x"76ffb338",
          9033 => x"783370bf",
          9034 => x"068d29f3",
          9035 => x"055b5581",
          9036 => x"77595683",
          9037 => x"e4e41833",
          9038 => x"79058111",
          9039 => x"33713371",
          9040 => x"882b0752",
          9041 => x"42577580",
          9042 => x"2e80ed38",
          9043 => x"7981fe26",
          9044 => x"ff843876",
          9045 => x"5181a18a",
          9046 => x"3f84b8e4",
          9047 => x"087a1061",
          9048 => x"05702253",
          9049 => x"43811b5b",
          9050 => x"5681a0f6",
          9051 => x"3f7584b8",
          9052 => x"e4082e09",
          9053 => x"8106fede",
          9054 => x"38765681",
          9055 => x"18588c78",
          9056 => x"27ffb038",
          9057 => x"78337086",
          9058 => x"2a810656",
          9059 => x"5975802e",
          9060 => x"92387480",
          9061 => x"2e8d3879",
          9062 => x"10600570",
          9063 => x"2241417f",
          9064 => x"feb438ff",
          9065 => x"1d7081ff",
          9066 => x"065e5afe",
          9067 => x"ae39840b",
          9068 => x"84b8e40c",
          9069 => x"933d0d04",
          9070 => x"7683ffff",
          9071 => x"2effbc38",
          9072 => x"81ff55fe",
          9073 => x"9439ea3d",
          9074 => x"0d687008",
          9075 => x"70ab1333",
          9076 => x"81a00658",
          9077 => x"5a5d5e86",
          9078 => x"567485b5",
          9079 => x"38748c1d",
          9080 => x"08702257",
          9081 => x"575d7480",
          9082 => x"2e8e3881",
          9083 => x"1d701017",
          9084 => x"70225156",
          9085 => x"5d74f438",
          9086 => x"953da01f",
          9087 => x"5b408c60",
          9088 => x"7b585855",
          9089 => x"75708105",
          9090 => x"57337770",
          9091 => x"81055934",
          9092 => x"ff155574",
          9093 => x"ef380280",
          9094 => x"db053370",
          9095 => x"81065856",
          9096 => x"76802e82",
          9097 => x"aa3880c0",
          9098 => x"0bab1f34",
          9099 => x"810b943d",
          9100 => x"405b8c1c",
          9101 => x"087b5859",
          9102 => x"8b7a615a",
          9103 => x"57557770",
          9104 => x"81055933",
          9105 => x"76708105",
          9106 => x"5834ff15",
          9107 => x"5574ef38",
          9108 => x"857b2780",
          9109 => x"c2387a79",
          9110 => x"22565774",
          9111 => x"802eb838",
          9112 => x"74821a5a",
          9113 => x"568f5875",
          9114 => x"81067710",
          9115 => x"0776812a",
          9116 => x"7083ffff",
          9117 => x"0672902a",
          9118 => x"81064458",
          9119 => x"56576080",
          9120 => x"2e873876",
          9121 => x"84a0a132",
          9122 => x"57ff1858",
          9123 => x"778025d7",
          9124 => x"38782255",
          9125 => x"74ca3887",
          9126 => x"02840580",
          9127 => x"cf055758",
          9128 => x"76b007bf",
          9129 => x"0655b975",
          9130 => x"27843887",
          9131 => x"15557476",
          9132 => x"34ff16ff",
          9133 => x"1978842a",
          9134 => x"59595676",
          9135 => x"e338771f",
          9136 => x"5980fe79",
          9137 => x"34767a58",
          9138 => x"56807827",
          9139 => x"a0387933",
          9140 => x"5574a02e",
          9141 => x"98388116",
          9142 => x"56757827",
          9143 => x"88a23875",
          9144 => x"1a703356",
          9145 => x"5774a02e",
          9146 => x"098106ea",
          9147 => x"38811656",
          9148 => x"a0557787",
          9149 => x"268e3898",
          9150 => x"3d7805ec",
          9151 => x"05811971",
          9152 => x"33575941",
          9153 => x"74773487",
          9154 => x"762787f4",
          9155 => x"387d51f8",
          9156 => x"8f3f84b8",
          9157 => x"e4088b38",
          9158 => x"811b5b80",
          9159 => x"e37b27fe",
          9160 => x"91388756",
          9161 => x"7a80e42e",
          9162 => x"82e73884",
          9163 => x"b8e40856",
          9164 => x"84b8e408",
          9165 => x"842e0981",
          9166 => x"0682d638",
          9167 => x"0280db05",
          9168 => x"33ab1f34",
          9169 => x"7d080284",
          9170 => x"0580db05",
          9171 => x"33575875",
          9172 => x"812a8106",
          9173 => x"5f815b7e",
          9174 => x"802e9038",
          9175 => x"8d528c1d",
          9176 => x"51fe8ac1",
          9177 => x"3f84b8e4",
          9178 => x"081b5b80",
          9179 => x"527d51ed",
          9180 => x"8c3f84b8",
          9181 => x"e4085684",
          9182 => x"b8e40881",
          9183 => x"823884b8",
          9184 => x"e408b819",
          9185 => x"5e59981e",
          9186 => x"08568057",
          9187 => x"b4180876",
          9188 => x"2e85f338",
          9189 => x"83183340",
          9190 => x"7f772e09",
          9191 => x"810682a3",
          9192 => x"38815475",
          9193 => x"53b81852",
          9194 => x"81183351",
          9195 => x"d4a43f84",
          9196 => x"b8e40880",
          9197 => x"2e8538ff",
          9198 => x"56815775",
          9199 => x"b4190c76",
          9200 => x"5676bc38",
          9201 => x"9c1e0870",
          9202 => x"33564274",
          9203 => x"81e52e81",
          9204 => x"c9387430",
          9205 => x"70802578",
          9206 => x"07565f74",
          9207 => x"802e81c9",
          9208 => x"38811959",
          9209 => x"787b2e86",
          9210 => x"89388152",
          9211 => x"7d51ee83",
          9212 => x"3f84b8e4",
          9213 => x"085684b8",
          9214 => x"e408802e",
          9215 => x"ff883887",
          9216 => x"5875842e",
          9217 => x"81893875",
          9218 => x"58758183",
          9219 => x"38ff1b40",
          9220 => x"7f81f338",
          9221 => x"981e0857",
          9222 => x"b41c0877",
          9223 => x"2eaf3883",
          9224 => x"1c337857",
          9225 => x"407f8482",
          9226 => x"38815476",
          9227 => x"53b81c52",
          9228 => x"811c3351",
          9229 => x"d39c3f84",
          9230 => x"b8e40880",
          9231 => x"2e8538ff",
          9232 => x"57815676",
          9233 => x"b41d0c75",
          9234 => x"587580c3",
          9235 => x"38a00b9c",
          9236 => x"1f085755",
          9237 => x"80767081",
          9238 => x"055834ff",
          9239 => x"155574f4",
          9240 => x"388b0b9c",
          9241 => x"1f087b58",
          9242 => x"58557570",
          9243 => x"81055733",
          9244 => x"77708105",
          9245 => x"5934ff15",
          9246 => x"5574ef38",
          9247 => x"9c1e08ab",
          9248 => x"1f339806",
          9249 => x"5e5a7c8c",
          9250 => x"1b34810b",
          9251 => x"831d3477",
          9252 => x"567584b8",
          9253 => x"e40c983d",
          9254 => x"0d048175",
          9255 => x"30708025",
          9256 => x"72075740",
          9257 => x"5774feb9",
          9258 => x"38745981",
          9259 => x"527d51ec",
          9260 => x"c23f84b8",
          9261 => x"e4085684",
          9262 => x"b8e40880",
          9263 => x"2efdc738",
          9264 => x"febd3981",
          9265 => x"54b41808",
          9266 => x"537c5281",
          9267 => x"183351d3",
          9268 => x"803f84b8",
          9269 => x"e408772e",
          9270 => x"09810683",
          9271 => x"bf3884b8",
          9272 => x"e4088319",
          9273 => x"34b41808",
          9274 => x"a8190831",
          9275 => x"5574a019",
          9276 => x"08278b38",
          9277 => x"82183341",
          9278 => x"60822e84",
          9279 => x"ac3884b8",
          9280 => x"e40857fd",
          9281 => x"9c397f85",
          9282 => x"2b901f08",
          9283 => x"71315358",
          9284 => x"7d51e9e9",
          9285 => x"3f84b8e4",
          9286 => x"085884b8",
          9287 => x"e408feef",
          9288 => x"387984b8",
          9289 => x"e4085658",
          9290 => x"8b577481",
          9291 => x"2a758180",
          9292 => x"29057870",
          9293 => x"81055a33",
          9294 => x"57760570",
          9295 => x"81ff06ff",
          9296 => x"1959565d",
          9297 => x"76e43874",
          9298 => x"81ff06b8",
          9299 => x"1d434198",
          9300 => x"1e085780",
          9301 => x"56b41c08",
          9302 => x"772eb238",
          9303 => x"831c335b",
          9304 => x"7a762e09",
          9305 => x"810682c9",
          9306 => x"38815476",
          9307 => x"53b81c52",
          9308 => x"811c3351",
          9309 => x"d0dc3f84",
          9310 => x"b8e40880",
          9311 => x"2e8538ff",
          9312 => x"57815676",
          9313 => x"b41d0c75",
          9314 => x"5875fe83",
          9315 => x"388c1c08",
          9316 => x"9c1f0861",
          9317 => x"81ff065f",
          9318 => x"5c5f608d",
          9319 => x"1c348f0b",
          9320 => x"8b1c3475",
          9321 => x"8c1c3475",
          9322 => x"9a1c3475",
          9323 => x"9b1c347c",
          9324 => x"8d29f305",
          9325 => x"76775a58",
          9326 => x"597683ff",
          9327 => x"ff2e8b38",
          9328 => x"78101f70",
          9329 => x"22811b5b",
          9330 => x"585683e4",
          9331 => x"e418337b",
          9332 => x"05557675",
          9333 => x"70810557",
          9334 => x"3476882a",
          9335 => x"56757534",
          9336 => x"76853883",
          9337 => x"ffff5781",
          9338 => x"18588c78",
          9339 => x"27cb3876",
          9340 => x"83ffff2e",
          9341 => x"81b33878",
          9342 => x"101f7022",
          9343 => x"58587680",
          9344 => x"2e81a638",
          9345 => x"7c7b3481",
          9346 => x"0b831d34",
          9347 => x"80527d51",
          9348 => x"e9e13f84",
          9349 => x"b8e40858",
          9350 => x"84b8e408",
          9351 => x"fcf1387f",
          9352 => x"ff05407f",
          9353 => x"fea938fb",
          9354 => x"eb398154",
          9355 => x"b41c0853",
          9356 => x"b81c7053",
          9357 => x"811d3352",
          9358 => x"59d0963f",
          9359 => x"815684b8",
          9360 => x"e408fc83",
          9361 => x"3884b8e4",
          9362 => x"08831d34",
          9363 => x"b41c08a8",
          9364 => x"1d083184",
          9365 => x"b8e40857",
          9366 => x"4160a01d",
          9367 => x"0827fbc9",
          9368 => x"38821c33",
          9369 => x"4261822e",
          9370 => x"098106fb",
          9371 => x"bc388154",
          9372 => x"b41c08a0",
          9373 => x"1d080553",
          9374 => x"7852811c",
          9375 => x"3351cfd1",
          9376 => x"3f7756fb",
          9377 => x"a439769c",
          9378 => x"1f087033",
          9379 => x"57435674",
          9380 => x"81e52e09",
          9381 => x"8106faba",
          9382 => x"38fbff39",
          9383 => x"81705757",
          9384 => x"76802efa",
          9385 => x"9f38fad7",
          9386 => x"397c80c0",
          9387 => x"075dfed4",
          9388 => x"398154b4",
          9389 => x"1c085361",
          9390 => x"52811c33",
          9391 => x"51cf923f",
          9392 => x"84b8e408",
          9393 => x"762e0981",
          9394 => x"06bc3884",
          9395 => x"b8e40883",
          9396 => x"1d34b41c",
          9397 => x"08a81d08",
          9398 => x"315574a0",
          9399 => x"1d08278a",
          9400 => x"38821c33",
          9401 => x"5f7e822e",
          9402 => x"aa3884b8",
          9403 => x"e40856fc",
          9404 => x"f83975ff",
          9405 => x"1c41587f",
          9406 => x"802efa98",
          9407 => x"38fc8739",
          9408 => x"751a57f7",
          9409 => x"e8398170",
          9410 => x"59567580",
          9411 => x"2efcfe38",
          9412 => x"fafd3981",
          9413 => x"54b41c08",
          9414 => x"a01d0805",
          9415 => x"53615281",
          9416 => x"1c3351ce",
          9417 => x"ac3ffcc1",
          9418 => x"398154b4",
          9419 => x"1808a019",
          9420 => x"0805537c",
          9421 => x"52811833",
          9422 => x"51ce963f",
          9423 => x"f8e339f3",
          9424 => x"3d0d7f61",
          9425 => x"7108405e",
          9426 => x"5c800b96",
          9427 => x"1e34981c",
          9428 => x"08802e82",
          9429 => x"b538ac1c",
          9430 => x"08ff2e80",
          9431 => x"d9388070",
          9432 => x"71608c05",
          9433 => x"08702257",
          9434 => x"585b5c58",
          9435 => x"72782ebc",
          9436 => x"38775474",
          9437 => x"14702281",
          9438 => x"1b5b5556",
          9439 => x"7a829538",
          9440 => x"80d08014",
          9441 => x"7083ffff",
          9442 => x"06585a76",
          9443 => x"8fff2682",
          9444 => x"83387379",
          9445 => x"1a761170",
          9446 => x"225d5855",
          9447 => x"5b79d438",
          9448 => x"7a307080",
          9449 => x"2570307a",
          9450 => x"065a5c5e",
          9451 => x"7c189405",
          9452 => x"57800b82",
          9453 => x"18348070",
          9454 => x"891f5957",
          9455 => x"589c1c08",
          9456 => x"16703381",
          9457 => x"18585653",
          9458 => x"74a02eb2",
          9459 => x"3874852e",
          9460 => x"81bc3875",
          9461 => x"89327030",
          9462 => x"70720780",
          9463 => x"25555b54",
          9464 => x"778b2690",
          9465 => x"3872802e",
          9466 => x"8b38ae77",
          9467 => x"70810559",
          9468 => x"34811858",
          9469 => x"74777081",
          9470 => x"05593481",
          9471 => x"18588a76",
          9472 => x"27ffba38",
          9473 => x"7c188805",
          9474 => x"55800b81",
          9475 => x"1634961d",
          9476 => x"335372a5",
          9477 => x"387781f3",
          9478 => x"38bf0b96",
          9479 => x"1e348157",
          9480 => x"7c179405",
          9481 => x"56800b82",
          9482 => x"17349c1c",
          9483 => x"088c1133",
          9484 => x"55537389",
          9485 => x"3873891e",
          9486 => x"349c1c08",
          9487 => x"538b1333",
          9488 => x"881e349c",
          9489 => x"1c089c11",
          9490 => x"83113382",
          9491 => x"12337190",
          9492 => x"2b71882b",
          9493 => x"07811433",
          9494 => x"70720788",
          9495 => x"2b753371",
          9496 => x"07640c59",
          9497 => x"97163396",
          9498 => x"17337188",
          9499 => x"2b075f41",
          9500 => x"5b405a56",
          9501 => x"5b557786",
          9502 => x"1e239915",
          9503 => x"33981633",
          9504 => x"71882b07",
          9505 => x"5d547b84",
          9506 => x"1e238f3d",
          9507 => x"0d0481e5",
          9508 => x"55fec039",
          9509 => x"771d9611",
          9510 => x"81ff7a31",
          9511 => x"585b5783",
          9512 => x"b5527a90",
          9513 => x"2b740751",
          9514 => x"8191893f",
          9515 => x"84b8e408",
          9516 => x"83ffff06",
          9517 => x"5581ff75",
          9518 => x"27ad3881",
          9519 => x"762781b3",
          9520 => x"3874882a",
          9521 => x"54737a34",
          9522 => x"74971834",
          9523 => x"82780558",
          9524 => x"800b8c1f",
          9525 => x"08565b78",
          9526 => x"19751170",
          9527 => x"225c5754",
          9528 => x"79fd9038",
          9529 => x"fdba3974",
          9530 => x"30763070",
          9531 => x"78078025",
          9532 => x"72802507",
          9533 => x"58555775",
          9534 => x"80f93874",
          9535 => x"7a348178",
          9536 => x"0558800b",
          9537 => x"8c1f0856",
          9538 => x"5bcd3972",
          9539 => x"73891f33",
          9540 => x"5a575777",
          9541 => x"802efe88",
          9542 => x"387c961e",
          9543 => x"7e575954",
          9544 => x"891433ff",
          9545 => x"bf115a54",
          9546 => x"789926a4",
          9547 => x"389c1c08",
          9548 => x"8c113354",
          9549 => x"5b887627",
          9550 => x"b4387284",
          9551 => x"2a537281",
          9552 => x"065e7d80",
          9553 => x"2e8a38a0",
          9554 => x"147083ff",
          9555 => x"ff065553",
          9556 => x"73787081",
          9557 => x"055a3481",
          9558 => x"16811681",
          9559 => x"19718913",
          9560 => x"335e5759",
          9561 => x"565679ff",
          9562 => x"b738fdb4",
          9563 => x"3972832a",
          9564 => x"53cc3980",
          9565 => x"7b307080",
          9566 => x"25703073",
          9567 => x"06535d5f",
          9568 => x"58fca939",
          9569 => x"ef3d0d63",
          9570 => x"70087042",
          9571 => x"575c8065",
          9572 => x"70335755",
          9573 => x"5374af2e",
          9574 => x"83388153",
          9575 => x"7480dc2e",
          9576 => x"81df3872",
          9577 => x"802e81d9",
          9578 => x"38981608",
          9579 => x"881d0c73",
          9580 => x"33963d94",
          9581 => x"3d414255",
          9582 => x"9f752782",
          9583 => x"a7387342",
          9584 => x"8c160858",
          9585 => x"80576170",
          9586 => x"70810552",
          9587 => x"33555373",
          9588 => x"81df3872",
          9589 => x"7f0c73ff",
          9590 => x"2e81ec38",
          9591 => x"83ffff74",
          9592 => x"278b3876",
          9593 => x"10185680",
          9594 => x"76238117",
          9595 => x"577383ff",
          9596 => x"ff0670af",
          9597 => x"3270309f",
          9598 => x"73277180",
          9599 => x"2507575b",
          9600 => x"5b557382",
          9601 => x"90387480",
          9602 => x"dc2e8289",
          9603 => x"387480ff",
          9604 => x"26b23883",
          9605 => x"e4800b83",
          9606 => x"e4803370",
          9607 => x"81ff0656",
          9608 => x"54567380",
          9609 => x"2e81ab38",
          9610 => x"73752e8f",
          9611 => x"38811670",
          9612 => x"337081ff",
          9613 => x"06565456",
          9614 => x"73ee3872",
          9615 => x"81ff065b",
          9616 => x"7a818438",
          9617 => x"7681fe26",
          9618 => x"80fd3876",
          9619 => x"10185d74",
          9620 => x"7d238117",
          9621 => x"62707081",
          9622 => x"05523356",
          9623 => x"54577380",
          9624 => x"2efef038",
          9625 => x"80cb3981",
          9626 => x"7380dc32",
          9627 => x"70307080",
          9628 => x"25730751",
          9629 => x"55585572",
          9630 => x"802ea138",
          9631 => x"81147046",
          9632 => x"54807433",
          9633 => x"545572af",
          9634 => x"2edd3872",
          9635 => x"80dc3270",
          9636 => x"30708025",
          9637 => x"77075154",
          9638 => x"5772e138",
          9639 => x"72881d0c",
          9640 => x"7333963d",
          9641 => x"943d4142",
          9642 => x"55749f26",
          9643 => x"fe9038b4",
          9644 => x"3983b552",
          9645 => x"7351818d",
          9646 => x"e73f84b8",
          9647 => x"e40883ff",
          9648 => x"ff065473",
          9649 => x"fe8d3886",
          9650 => x"547384b8",
          9651 => x"e40c933d",
          9652 => x"0d0483e4",
          9653 => x"80337081",
          9654 => x"ff065c53",
          9655 => x"7a802efe",
          9656 => x"e338e439",
          9657 => x"ff800bab",
          9658 => x"1d348052",
          9659 => x"7b51de8d",
          9660 => x"3f84b8e4",
          9661 => x"0884b8e4",
          9662 => x"0c933d0d",
          9663 => x"04817380",
          9664 => x"dc327030",
          9665 => x"70802573",
          9666 => x"0741555a",
          9667 => x"567d802e",
          9668 => x"a1388114",
          9669 => x"42806270",
          9670 => x"33555556",
          9671 => x"72af2edd",
          9672 => x"387280dc",
          9673 => x"32703070",
          9674 => x"80257807",
          9675 => x"4054597d",
          9676 => x"e1387361",
          9677 => x"0c9f7527",
          9678 => x"822b5a76",
          9679 => x"812e84f8",
          9680 => x"3876822e",
          9681 => x"83d13876",
          9682 => x"17597680",
          9683 => x"2ea73876",
          9684 => x"177811fe",
          9685 => x"05702270",
          9686 => x"a0327030",
          9687 => x"709f2a52",
          9688 => x"42565f56",
          9689 => x"597cae2e",
          9690 => x"84387289",
          9691 => x"38ff1757",
          9692 => x"76dd3876",
          9693 => x"59771956",
          9694 => x"80762376",
          9695 => x"802efec7",
          9696 => x"38807822",
          9697 => x"7083ffff",
          9698 => x"0672585d",
          9699 => x"55567aa0",
          9700 => x"2e82e638",
          9701 => x"7383ffff",
          9702 => x"065372ae",
          9703 => x"2e82f138",
          9704 => x"76802eaa",
          9705 => x"387719fe",
          9706 => x"0570225a",
          9707 => x"5478ae2e",
          9708 => x"9d387610",
          9709 => x"18fe0554",
          9710 => x"ff175776",
          9711 => x"802e8f38",
          9712 => x"fe147022",
          9713 => x"5e547cae",
          9714 => x"2e098106",
          9715 => x"eb388b0b",
          9716 => x"a01d5553",
          9717 => x"a0747081",
          9718 => x"055634ff",
          9719 => x"135372f4",
          9720 => x"3872735c",
          9721 => x"5e887816",
          9722 => x"70228119",
          9723 => x"5957545d",
          9724 => x"74802e80",
          9725 => x"ed3874a0",
          9726 => x"2e83d038",
          9727 => x"74ae3270",
          9728 => x"30708025",
          9729 => x"555a5475",
          9730 => x"772e85ce",
          9731 => x"387283bb",
          9732 => x"3872597c",
          9733 => x"7b268338",
          9734 => x"81597577",
          9735 => x"32703070",
          9736 => x"72078025",
          9737 => x"707c0751",
          9738 => x"51545472",
          9739 => x"802e83e0",
          9740 => x"387c8b2e",
          9741 => x"86833875",
          9742 => x"772e8a38",
          9743 => x"7983075a",
          9744 => x"7577269e",
          9745 => x"38765688",
          9746 => x"5b8b7e82",
          9747 => x"2b81fc06",
          9748 => x"7718575f",
          9749 => x"5d771570",
          9750 => x"22811858",
          9751 => x"565374ff",
          9752 => x"9538a01c",
          9753 => x"33577681",
          9754 => x"e52e8384",
          9755 => x"387c882e",
          9756 => x"82e3387d",
          9757 => x"8c065877",
          9758 => x"8c2e82ed",
          9759 => x"387d8306",
          9760 => x"5574832e",
          9761 => x"82e33879",
          9762 => x"812a8106",
          9763 => x"56759d38",
          9764 => x"7d81065d",
          9765 => x"7c802e85",
          9766 => x"38799007",
          9767 => x"5a7d822a",
          9768 => x"81065e7d",
          9769 => x"802e8538",
          9770 => x"7988075a",
          9771 => x"79ab1d34",
          9772 => x"7b51e4ec",
          9773 => x"3f84b8e4",
          9774 => x"08ab1d33",
          9775 => x"565484b8",
          9776 => x"e408802e",
          9777 => x"81ac3884",
          9778 => x"b8e40884",
          9779 => x"2e098106",
          9780 => x"fbf73874",
          9781 => x"852a8106",
          9782 => x"5a79802e",
          9783 => x"84f03874",
          9784 => x"822a8106",
          9785 => x"59788298",
          9786 => x"387b0865",
          9787 => x"55567342",
          9788 => x"8c160858",
          9789 => x"8057f9ce",
          9790 => x"39811670",
          9791 => x"11791170",
          9792 => x"22404056",
          9793 => x"567ca02e",
          9794 => x"f0387580",
          9795 => x"2efd8538",
          9796 => x"7983075a",
          9797 => x"fd8a3982",
          9798 => x"18225675",
          9799 => x"ae2e0981",
          9800 => x"06fcac38",
          9801 => x"77225473",
          9802 => x"ae2e0981",
          9803 => x"06fca038",
          9804 => x"7610185b",
          9805 => x"807b2380",
          9806 => x"0ba01d56",
          9807 => x"53ae5476",
          9808 => x"73268338",
          9809 => x"a0547375",
          9810 => x"70810557",
          9811 => x"34811353",
          9812 => x"8a7327e9",
          9813 => x"3879a007",
          9814 => x"5877ab1d",
          9815 => x"347b51e3",
          9816 => x"bf3f84b8",
          9817 => x"e408ab1d",
          9818 => x"33565484",
          9819 => x"b8e408fe",
          9820 => x"d6387482",
          9821 => x"2a810658",
          9822 => x"77face38",
          9823 => x"861c3370",
          9824 => x"842a8106",
          9825 => x"565d7480",
          9826 => x"2e83cd38",
          9827 => x"901c0883",
          9828 => x"ff066005",
          9829 => x"80d31133",
          9830 => x"80d21233",
          9831 => x"71882b07",
          9832 => x"62334157",
          9833 => x"54547d83",
          9834 => x"2e82d838",
          9835 => x"74881d0c",
          9836 => x"7b086555",
          9837 => x"56feb739",
          9838 => x"77225574",
          9839 => x"ae2efef0",
          9840 => x"38761759",
          9841 => x"76fb8838",
          9842 => x"fbab3979",
          9843 => x"83077617",
          9844 => x"565afd81",
          9845 => x"397d822b",
          9846 => x"81fc0670",
          9847 => x"8c06595e",
          9848 => x"778c2e09",
          9849 => x"8106fd95",
          9850 => x"38798207",
          9851 => x"5afd9839",
          9852 => x"850ba01d",
          9853 => x"347c882e",
          9854 => x"098106fc",
          9855 => x"f638d639",
          9856 => x"ff800bab",
          9857 => x"1d34800b",
          9858 => x"84b8e40c",
          9859 => x"933d0d04",
          9860 => x"7480ff26",
          9861 => x"9d3881ff",
          9862 => x"752780c9",
          9863 => x"38ff1d59",
          9864 => x"787b2681",
          9865 => x"f7387983",
          9866 => x"077d7718",
          9867 => x"575c5afc",
          9868 => x"a4397982",
          9869 => x"075a83b5",
          9870 => x"52745181",
          9871 => x"85f63f84",
          9872 => x"b8e40883",
          9873 => x"ffff0670",
          9874 => x"872a8106",
          9875 => x"5a557880",
          9876 => x"2ec43874",
          9877 => x"80ff0683",
          9878 => x"e4f41133",
          9879 => x"56547481",
          9880 => x"ff26ffb9",
          9881 => x"3874802e",
          9882 => x"81853883",
          9883 => x"e48c0b83",
          9884 => x"e48c3370",
          9885 => x"81ff0656",
          9886 => x"54597380",
          9887 => x"2e80e038",
          9888 => x"73752e8f",
          9889 => x"38811970",
          9890 => x"337081ff",
          9891 => x"06565459",
          9892 => x"73ee3872",
          9893 => x"81ff0659",
          9894 => x"7880d438",
          9895 => x"ffbf1554",
          9896 => x"7399268a",
          9897 => x"387d8207",
          9898 => x"7081ff06",
          9899 => x"5f53ff9f",
          9900 => x"15597899",
          9901 => x"2693387d",
          9902 => x"81077081",
          9903 => x"ff06e017",
          9904 => x"7083ffff",
          9905 => x"0658565f",
          9906 => x"537b1ba0",
          9907 => x"05597479",
          9908 => x"34811b5b",
          9909 => x"751655fa",
          9910 => x"fc398053",
          9911 => x"fab33983",
          9912 => x"e48c3370",
          9913 => x"81ff065a",
          9914 => x"5378802e",
          9915 => x"ffae3880",
          9916 => x"df7a8307",
          9917 => x"7d1da005",
          9918 => x"5b5b5574",
          9919 => x"7934811b",
          9920 => x"5bd23980",
          9921 => x"cd143380",
          9922 => x"cc153371",
          9923 => x"982b7190",
          9924 => x"2b077707",
          9925 => x"881f0c5a",
          9926 => x"57fd9539",
          9927 => x"7b1ba005",
          9928 => x"75882a54",
          9929 => x"54727434",
          9930 => x"811b7c11",
          9931 => x"a0055a5b",
          9932 => x"74793481",
          9933 => x"1b5bff9c",
          9934 => x"39798307",
          9935 => x"a01d3358",
          9936 => x"5a7681e5",
          9937 => x"2e098106",
          9938 => x"faa338fd",
          9939 => x"a3397482",
          9940 => x"2a81065c",
          9941 => x"7bf6f238",
          9942 => x"850b84b8",
          9943 => x"e40c933d",
          9944 => x"0d04eb3d",
          9945 => x"0d676902",
          9946 => x"880580e7",
          9947 => x"05334242",
          9948 => x"5e80610c",
          9949 => x"ff7e0870",
          9950 => x"595b4279",
          9951 => x"802e85d7",
          9952 => x"38797081",
          9953 => x"055b3370",
          9954 => x"9f265656",
          9955 => x"75ba2e85",
          9956 => x"d03874ed",
          9957 => x"3875ba2e",
          9958 => x"85c73884",
          9959 => x"d0c03356",
          9960 => x"80762485",
          9961 => x"b2387510",
          9962 => x"1084d0ac",
          9963 => x"05700858",
          9964 => x"5a8c5876",
          9965 => x"802e8596",
          9966 => x"3876610c",
          9967 => x"7f81fe06",
          9968 => x"77335d59",
          9969 => x"7b802e9b",
          9970 => x"38811733",
          9971 => x"51ffbbb0",
          9972 => x"3f84b8e4",
          9973 => x"0881ff06",
          9974 => x"7081065e",
          9975 => x"587c802e",
          9976 => x"86963880",
          9977 => x"77347516",
          9978 => x"5d84b8d8",
          9979 => x"1d338118",
          9980 => x"34815281",
          9981 => x"173351ff",
          9982 => x"bba43f84",
          9983 => x"b8e40881",
          9984 => x"ff067081",
          9985 => x"06415683",
          9986 => x"587f84c2",
          9987 => x"3878802e",
          9988 => x"8d387582",
          9989 => x"2a810641",
          9990 => x"8a586084",
          9991 => x"b138805b",
          9992 => x"7a831834",
          9993 => x"ff0bb418",
          9994 => x"0c7a7b5a",
          9995 => x"5581547a",
          9996 => x"53b81770",
          9997 => x"53811833",
          9998 => x"5258ffbb",
          9999 => x"953f84b8",
         10000 => x"e4087b2e",
         10001 => x"8538ff55",
         10002 => x"815974b4",
         10003 => x"180c8456",
         10004 => x"78993884",
         10005 => x"b7173384",
         10006 => x"b6183371",
         10007 => x"882b0756",
         10008 => x"56835674",
         10009 => x"82d4d52e",
         10010 => x"85a53875",
         10011 => x"81268b38",
         10012 => x"84b8d91d",
         10013 => x"33426185",
         10014 => x"bf388158",
         10015 => x"75842e83",
         10016 => x"cd388d58",
         10017 => x"75812683",
         10018 => x"c53880c4",
         10019 => x"173380c3",
         10020 => x"18337188",
         10021 => x"2b075e59",
         10022 => x"7c84802e",
         10023 => x"09810683",
         10024 => x"ad3880cf",
         10025 => x"173380ce",
         10026 => x"18337188",
         10027 => x"2b07575a",
         10028 => x"75a43880",
         10029 => x"dc178311",
         10030 => x"33821233",
         10031 => x"71902b71",
         10032 => x"882b0781",
         10033 => x"14337072",
         10034 => x"07882b75",
         10035 => x"33710756",
         10036 => x"5a45435e",
         10037 => x"5f5675a0",
         10038 => x"180c80c8",
         10039 => x"17338218",
         10040 => x"3480c817",
         10041 => x"33ff1170",
         10042 => x"81ff065f",
         10043 => x"40598d58",
         10044 => x"7c812682",
         10045 => x"d9387881",
         10046 => x"ff067671",
         10047 => x"2980c519",
         10048 => x"335a5f5a",
         10049 => x"778a1823",
         10050 => x"77597780",
         10051 => x"2e87c438",
         10052 => x"ff187806",
         10053 => x"426187bb",
         10054 => x"3880ca17",
         10055 => x"3380c918",
         10056 => x"3371882b",
         10057 => x"07564074",
         10058 => x"88182374",
         10059 => x"758f065e",
         10060 => x"5a8d587c",
         10061 => x"82983880",
         10062 => x"cc173380",
         10063 => x"cb183371",
         10064 => x"882b0756",
         10065 => x"5c74a438",
         10066 => x"80d81783",
         10067 => x"11338212",
         10068 => x"3371902b",
         10069 => x"71882b07",
         10070 => x"81143370",
         10071 => x"7207882b",
         10072 => x"75337107",
         10073 => x"53445a58",
         10074 => x"42424280",
         10075 => x"c7173380",
         10076 => x"c6183371",
         10077 => x"882b075d",
         10078 => x"588d587b",
         10079 => x"802e81ce",
         10080 => x"387d1c7a",
         10081 => x"842a055a",
         10082 => x"79752681",
         10083 => x"c1387852",
         10084 => x"747a3151",
         10085 => x"fdee8e3f",
         10086 => x"84b8e408",
         10087 => x"5684b8e4",
         10088 => x"08802e81",
         10089 => x"a93884b8",
         10090 => x"e40880ff",
         10091 => x"fffff526",
         10092 => x"8338835d",
         10093 => x"7583fff5",
         10094 => x"26833882",
         10095 => x"5d759ff5",
         10096 => x"2685eb38",
         10097 => x"815d8216",
         10098 => x"709c190c",
         10099 => x"7ba4190c",
         10100 => x"7b1d70a8",
         10101 => x"1a0c7b1d",
         10102 => x"b01a0c57",
         10103 => x"597c832e",
         10104 => x"8a873888",
         10105 => x"17225c8d",
         10106 => x"587b802e",
         10107 => x"80e0387d",
         10108 => x"16ac180c",
         10109 => x"7819557c",
         10110 => x"822e8d38",
         10111 => x"78101970",
         10112 => x"812a7a81",
         10113 => x"0605565a",
         10114 => x"83ff1589",
         10115 => x"2a598d58",
         10116 => x"78a01808",
         10117 => x"26b838ff",
         10118 => x"0b94180c",
         10119 => x"ff0b9018",
         10120 => x"0cff800b",
         10121 => x"8418347c",
         10122 => x"832e8696",
         10123 => x"387c7734",
         10124 => x"84d0bc22",
         10125 => x"81055d7c",
         10126 => x"84d0bc23",
         10127 => x"7c861823",
         10128 => x"84d0c40b",
         10129 => x"8c180c80",
         10130 => x"0b98180c",
         10131 => x"80587784",
         10132 => x"b8e40c97",
         10133 => x"3d0d048b",
         10134 => x"0b84b8e4",
         10135 => x"0c973d0d",
         10136 => x"047633d0",
         10137 => x"117081ff",
         10138 => x"06575758",
         10139 => x"74892691",
         10140 => x"38821778",
         10141 => x"81ff06d0",
         10142 => x"055d5978",
         10143 => x"7a2e87fe",
         10144 => x"38807e08",
         10145 => x"83e4d45f",
         10146 => x"405c7c08",
         10147 => x"7f5a5b7a",
         10148 => x"7081055c",
         10149 => x"33797081",
         10150 => x"055b33ff",
         10151 => x"9f125a58",
         10152 => x"56779926",
         10153 => x"8938e016",
         10154 => x"7081ff06",
         10155 => x"5755ff9f",
         10156 => x"17587799",
         10157 => x"268938e0",
         10158 => x"177081ff",
         10159 => x"06585575",
         10160 => x"30709f2a",
         10161 => x"59557577",
         10162 => x"2e098106",
         10163 => x"853877ff",
         10164 => x"be38787a",
         10165 => x"32703070",
         10166 => x"72079f2a",
         10167 => x"7a075d58",
         10168 => x"557a802e",
         10169 => x"87983881",
         10170 => x"1c841e5e",
         10171 => x"5c837c25",
         10172 => x"ff983861",
         10173 => x"56f9a939",
         10174 => x"78802efe",
         10175 => x"cf387782",
         10176 => x"2a81065e",
         10177 => x"8a587dfe",
         10178 => x"c5388058",
         10179 => x"fec0397a",
         10180 => x"78335759",
         10181 => x"7581e92e",
         10182 => x"09810683",
         10183 => x"38815975",
         10184 => x"81eb3270",
         10185 => x"30708025",
         10186 => x"7b075a5b",
         10187 => x"5c7783ad",
         10188 => x"387581e8",
         10189 => x"2e83a638",
         10190 => x"933d7757",
         10191 => x"5a835983",
         10192 => x"fa163370",
         10193 => x"595b7a80",
         10194 => x"2ea53884",
         10195 => x"81163384",
         10196 => x"80173371",
         10197 => x"902b7188",
         10198 => x"2b0783ff",
         10199 => x"19337072",
         10200 => x"07882b83",
         10201 => x"fe1b3371",
         10202 => x"0752595b",
         10203 => x"40404077",
         10204 => x"7a708405",
         10205 => x"5c0cff19",
         10206 => x"90175759",
         10207 => x"788025ff",
         10208 => x"be3884b8",
         10209 => x"d91d3370",
         10210 => x"30709f2a",
         10211 => x"7271319b",
         10212 => x"3d711010",
         10213 => x"05f00584",
         10214 => x"b61c445d",
         10215 => x"52435b42",
         10216 => x"78085b83",
         10217 => x"567a802e",
         10218 => x"80fb3880",
         10219 => x"0b831834",
         10220 => x"ff0bb418",
         10221 => x"0c7a5580",
         10222 => x"567aff2e",
         10223 => x"a5388154",
         10224 => x"7a53b817",
         10225 => x"52811733",
         10226 => x"51ffb486",
         10227 => x"3f84b8e4",
         10228 => x"08762e85",
         10229 => x"38ff5581",
         10230 => x"5674b418",
         10231 => x"0c845875",
         10232 => x"bf38811f",
         10233 => x"337f3371",
         10234 => x"882b075d",
         10235 => x"5e83587b",
         10236 => x"82d4d52e",
         10237 => x"098106a8",
         10238 => x"38800bb8",
         10239 => x"18335758",
         10240 => x"7581e92e",
         10241 => x"82b73875",
         10242 => x"81eb3270",
         10243 => x"30708025",
         10244 => x"7a074242",
         10245 => x"427fbc38",
         10246 => x"7581e82e",
         10247 => x"b6388258",
         10248 => x"7781ff06",
         10249 => x"56800b84",
         10250 => x"b8d91e33",
         10251 => x"5d587b78",
         10252 => x"2e098106",
         10253 => x"83388158",
         10254 => x"817627f8",
         10255 => x"bd387780",
         10256 => x"2ef8b738",
         10257 => x"811a841a",
         10258 => x"5a5a837a",
         10259 => x"27fed138",
         10260 => x"f8a83983",
         10261 => x"0b80ee18",
         10262 => x"83e49440",
         10263 => x"5d587b70",
         10264 => x"81055d33",
         10265 => x"7e708105",
         10266 => x"40337171",
         10267 => x"31ff1b5b",
         10268 => x"52565677",
         10269 => x"802e80c5",
         10270 => x"3875802e",
         10271 => x"e138850b",
         10272 => x"818a1883",
         10273 => x"e498405d",
         10274 => x"587b7081",
         10275 => x"055d337e",
         10276 => x"70810540",
         10277 => x"33717131",
         10278 => x"ff1b5b58",
         10279 => x"42407780",
         10280 => x"2e858e38",
         10281 => x"75802ee1",
         10282 => x"388258fe",
         10283 => x"f3398d58",
         10284 => x"7cfa9338",
         10285 => x"7784b8e4",
         10286 => x"0c973d0d",
         10287 => x"04755875",
         10288 => x"802efedc",
         10289 => x"38850b81",
         10290 => x"8a1883e4",
         10291 => x"98405d58",
         10292 => x"ffb7398d",
         10293 => x"0b84b8e4",
         10294 => x"0c973d0d",
         10295 => x"04830b80",
         10296 => x"ee1883e4",
         10297 => x"945c5a58",
         10298 => x"78708105",
         10299 => x"5a337a70",
         10300 => x"81055c33",
         10301 => x"717131ff",
         10302 => x"1b5b575f",
         10303 => x"5f77802e",
         10304 => x"83d13874",
         10305 => x"802ee138",
         10306 => x"850b818a",
         10307 => x"1883e498",
         10308 => x"5c5a5878",
         10309 => x"7081055a",
         10310 => x"337a7081",
         10311 => x"055c3371",
         10312 => x"7131ff1b",
         10313 => x"5b584240",
         10314 => x"77802e84",
         10315 => x"91387580",
         10316 => x"2ee13893",
         10317 => x"3d77575a",
         10318 => x"8359fc83",
         10319 => x"398158fd",
         10320 => x"c63980e9",
         10321 => x"173380e8",
         10322 => x"18337188",
         10323 => x"2b075755",
         10324 => x"75812e09",
         10325 => x"8106f9d5",
         10326 => x"38811b58",
         10327 => x"805ab417",
         10328 => x"08782eb1",
         10329 => x"38831733",
         10330 => x"5b7a7a2e",
         10331 => x"09810682",
         10332 => x"9b388154",
         10333 => x"7753b817",
         10334 => x"52811733",
         10335 => x"51ffb0d2",
         10336 => x"3f84b8e4",
         10337 => x"08802e85",
         10338 => x"38ff5881",
         10339 => x"5a77b418",
         10340 => x"0c79f999",
         10341 => x"38798418",
         10342 => x"3484b717",
         10343 => x"3384b618",
         10344 => x"3371882b",
         10345 => x"07575e75",
         10346 => x"82d4d52e",
         10347 => x"098106f8",
         10348 => x"fc38b817",
         10349 => x"83113382",
         10350 => x"12337190",
         10351 => x"2b71882b",
         10352 => x"07811433",
         10353 => x"70720788",
         10354 => x"2b753371",
         10355 => x"075e4159",
         10356 => x"45425c59",
         10357 => x"77848b85",
         10358 => x"a4d22e09",
         10359 => x"8106f8cd",
         10360 => x"38849c17",
         10361 => x"83113382",
         10362 => x"12337190",
         10363 => x"2b71882b",
         10364 => x"07811433",
         10365 => x"70720788",
         10366 => x"2b753371",
         10367 => x"07474440",
         10368 => x"5b5c5a5e",
         10369 => x"60868a85",
         10370 => x"e4f22e09",
         10371 => x"8106f89d",
         10372 => x"3884a017",
         10373 => x"83113382",
         10374 => x"12337190",
         10375 => x"2b71882b",
         10376 => x"07811433",
         10377 => x"70720788",
         10378 => x"2b753371",
         10379 => x"07941e0c",
         10380 => x"5d84a41c",
         10381 => x"83113382",
         10382 => x"12337190",
         10383 => x"2b71882b",
         10384 => x"07811433",
         10385 => x"70720788",
         10386 => x"2b753371",
         10387 => x"07629005",
         10388 => x"0c594449",
         10389 => x"465c4540",
         10390 => x"455b565a",
         10391 => x"7c773484",
         10392 => x"d0bc2281",
         10393 => x"055d7c84",
         10394 => x"d0bc237c",
         10395 => x"86182384",
         10396 => x"d0c40b8c",
         10397 => x"180c800b",
         10398 => x"98180cf7",
         10399 => x"cf397b83",
         10400 => x"24f8f038",
         10401 => x"7b7a7f0c",
         10402 => x"56f29539",
         10403 => x"7554b417",
         10404 => x"0853b817",
         10405 => x"70538118",
         10406 => x"335259ff",
         10407 => x"afb33f84",
         10408 => x"b8e4087a",
         10409 => x"2e098106",
         10410 => x"81a43884",
         10411 => x"b8e40883",
         10412 => x"1834b417",
         10413 => x"08a81808",
         10414 => x"31407fa0",
         10415 => x"1808278b",
         10416 => x"38821733",
         10417 => x"4160822e",
         10418 => x"818d3884",
         10419 => x"b8e4085a",
         10420 => x"fda03974",
         10421 => x"5674802e",
         10422 => x"f3913885",
         10423 => x"0b818a18",
         10424 => x"83e4985c",
         10425 => x"5a58fcab",
         10426 => x"3980e317",
         10427 => x"3380e218",
         10428 => x"3371882b",
         10429 => x"075f5a8d",
         10430 => x"587df6d2",
         10431 => x"38881722",
         10432 => x"4261f6ca",
         10433 => x"3880e417",
         10434 => x"83113382",
         10435 => x"12337190",
         10436 => x"2b71882b",
         10437 => x"07811433",
         10438 => x"70720788",
         10439 => x"2b753371",
         10440 => x"07ac1e0c",
         10441 => x"5a7d822b",
         10442 => x"5a434440",
         10443 => x"5940f5d8",
         10444 => x"39755875",
         10445 => x"802ef9e8",
         10446 => x"388258f9",
         10447 => x"e3397580",
         10448 => x"2ef2a838",
         10449 => x"933d7757",
         10450 => x"5a8359f7",
         10451 => x"f239755a",
         10452 => x"79f5da38",
         10453 => x"fcbf3975",
         10454 => x"54b41708",
         10455 => x"a0180805",
         10456 => x"53785281",
         10457 => x"173351ff",
         10458 => x"ade73ffc",
         10459 => x"8539f03d",
         10460 => x"0d0280d3",
         10461 => x"05336470",
         10462 => x"43933d41",
         10463 => x"575dff76",
         10464 => x"5a407580",
         10465 => x"2e80e938",
         10466 => x"78708105",
         10467 => x"5a33709f",
         10468 => x"26555574",
         10469 => x"ba2e80e2",
         10470 => x"3873ed38",
         10471 => x"74ba2e80",
         10472 => x"d93884d0",
         10473 => x"c0335480",
         10474 => x"742480c4",
         10475 => x"38731010",
         10476 => x"84d0ac05",
         10477 => x"70085555",
         10478 => x"73802e84",
         10479 => x"38807434",
         10480 => x"62547380",
         10481 => x"2e863880",
         10482 => x"74346254",
         10483 => x"73750c7c",
         10484 => x"547c802e",
         10485 => x"92388053",
         10486 => x"933d7053",
         10487 => x"840551ef",
         10488 => x"813f84b8",
         10489 => x"e4085473",
         10490 => x"84b8e40c",
         10491 => x"923d0d04",
         10492 => x"8b0b84b8",
         10493 => x"e40c923d",
         10494 => x"0d047533",
         10495 => x"d0117081",
         10496 => x"ff065656",
         10497 => x"57738926",
         10498 => x"91388216",
         10499 => x"7781ff06",
         10500 => x"d0055c58",
         10501 => x"77792e80",
         10502 => x"f738807f",
         10503 => x"0883e4d4",
         10504 => x"5e5f5b7b",
         10505 => x"087e595a",
         10506 => x"79708105",
         10507 => x"5b337870",
         10508 => x"81055a33",
         10509 => x"ff9f1259",
         10510 => x"57557699",
         10511 => x"268938e0",
         10512 => x"157081ff",
         10513 => x"065654ff",
         10514 => x"9f165776",
         10515 => x"99268938",
         10516 => x"e0167081",
         10517 => x"ff065754",
         10518 => x"7430709f",
         10519 => x"2a585474",
         10520 => x"762e0981",
         10521 => x"06853876",
         10522 => x"ffbe3877",
         10523 => x"79327030",
         10524 => x"7072079f",
         10525 => x"2a79075c",
         10526 => x"57547980",
         10527 => x"2e923881",
         10528 => x"1b841d5d",
         10529 => x"5b837b25",
         10530 => x"ff99387f",
         10531 => x"54fe9839",
         10532 => x"7a8324f7",
         10533 => x"387a7960",
         10534 => x"0c54fe8b",
         10535 => x"39e63d0d",
         10536 => x"6c028405",
         10537 => x"80fb0533",
         10538 => x"56598956",
         10539 => x"78802ea6",
         10540 => x"3874bf06",
         10541 => x"70549d3d",
         10542 => x"cc05539e",
         10543 => x"3d840552",
         10544 => x"58ed9f3f",
         10545 => x"84b8e408",
         10546 => x"5784b8e4",
         10547 => x"08802e8f",
         10548 => x"3880790c",
         10549 => x"76567584",
         10550 => x"b8e40c9c",
         10551 => x"3d0d047e",
         10552 => x"406d5290",
         10553 => x"3d70525a",
         10554 => x"e19a3f84",
         10555 => x"b8e40857",
         10556 => x"84b8e408",
         10557 => x"802e81ba",
         10558 => x"38779c06",
         10559 => x"5d7c802e",
         10560 => x"81ca3876",
         10561 => x"802e83c1",
         10562 => x"3876842e",
         10563 => x"83ea3877",
         10564 => x"88075876",
         10565 => x"ffbb3877",
         10566 => x"832a8106",
         10567 => x"5b7a802e",
         10568 => x"81d13866",
         10569 => x"9b11339a",
         10570 => x"12337188",
         10571 => x"2b076170",
         10572 => x"3342585e",
         10573 => x"5e567d83",
         10574 => x"2e84e938",
         10575 => x"800b8e17",
         10576 => x"34800b8f",
         10577 => x"1734a10b",
         10578 => x"90173480",
         10579 => x"cc0b9117",
         10580 => x"346656a0",
         10581 => x"0b8b1734",
         10582 => x"7e67575e",
         10583 => x"800b9a17",
         10584 => x"34800b9b",
         10585 => x"17347d33",
         10586 => x"5d7c832e",
         10587 => x"84a93866",
         10588 => x"5b800b9c",
         10589 => x"1c34800b",
         10590 => x"9d1c3480",
         10591 => x"0b9e1c34",
         10592 => x"800b9f1c",
         10593 => x"347e5581",
         10594 => x"0b831634",
         10595 => x"7b802e80",
         10596 => x"e2387eb4",
         10597 => x"11087d7c",
         10598 => x"0853575f",
         10599 => x"57817c27",
         10600 => x"89389c17",
         10601 => x"087c2683",
         10602 => x"8a388257",
         10603 => x"80790cfe",
         10604 => x"a3390280",
         10605 => x"e7053370",
         10606 => x"982b5d5b",
         10607 => x"7b8025fe",
         10608 => x"b8388678",
         10609 => x"9c065e57",
         10610 => x"7cfeb838",
         10611 => x"76fe8238",
         10612 => x"0280c205",
         10613 => x"3370842a",
         10614 => x"81065d56",
         10615 => x"7b829138",
         10616 => x"77812a81",
         10617 => x"065e7d80",
         10618 => x"2e893875",
         10619 => x"81065a79",
         10620 => x"81f63877",
         10621 => x"832a8106",
         10622 => x"5675802e",
         10623 => x"86387780",
         10624 => x"c007587e",
         10625 => x"b41108a0",
         10626 => x"1b0c67a4",
         10627 => x"1b0c679b",
         10628 => x"11339a12",
         10629 => x"3371882b",
         10630 => x"07733340",
         10631 => x"5e40575a",
         10632 => x"7b832e81",
         10633 => x"f1387a88",
         10634 => x"1a0c9c16",
         10635 => x"83113382",
         10636 => x"12337190",
         10637 => x"2b71882b",
         10638 => x"07811433",
         10639 => x"70720788",
         10640 => x"2b753371",
         10641 => x"0770608c",
         10642 => x"050c6060",
         10643 => x"0c515241",
         10644 => x"59575d5e",
         10645 => x"861a2284",
         10646 => x"1a237790",
         10647 => x"1a34800b",
         10648 => x"911a3480",
         10649 => x"0b9c1a0c",
         10650 => x"77852a81",
         10651 => x"06557480",
         10652 => x"2e84ac38",
         10653 => x"75802e84",
         10654 => x"f1387594",
         10655 => x"1a0c8a1a",
         10656 => x"2270892b",
         10657 => x"7c525b58",
         10658 => x"76307078",
         10659 => x"07802556",
         10660 => x"5b797627",
         10661 => x"84923881",
         10662 => x"7076065f",
         10663 => x"5b7d802e",
         10664 => x"84863877",
         10665 => x"527851ff",
         10666 => x"acdb3f84",
         10667 => x"b8e40858",
         10668 => x"84b8e408",
         10669 => x"81268338",
         10670 => x"825784b8",
         10671 => x"e408ff2e",
         10672 => x"80cb3875",
         10673 => x"7a3156c0",
         10674 => x"390280c2",
         10675 => x"05339106",
         10676 => x"5e7d9538",
         10677 => x"77822a81",
         10678 => x"06557480",
         10679 => x"2efcb838",
         10680 => x"88578079",
         10681 => x"0cfbed39",
         10682 => x"87578079",
         10683 => x"0cfbe539",
         10684 => x"84578079",
         10685 => x"0cfbdd39",
         10686 => x"7951cdca",
         10687 => x"3f84b8e4",
         10688 => x"08788807",
         10689 => x"595776fb",
         10690 => x"c838fc8b",
         10691 => x"397a767b",
         10692 => x"315757fe",
         10693 => x"f3399516",
         10694 => x"33941733",
         10695 => x"71982b71",
         10696 => x"902b077d",
         10697 => x"075d5e5c",
         10698 => x"fdfc397c",
         10699 => x"557c7b27",
         10700 => x"81bd3874",
         10701 => x"527951ff",
         10702 => x"abcb3f84",
         10703 => x"b8e4085d",
         10704 => x"84b8e408",
         10705 => x"802e81a7",
         10706 => x"3884b8e4",
         10707 => x"08812efc",
         10708 => x"d93884b8",
         10709 => x"e408ff2e",
         10710 => x"83993880",
         10711 => x"53745276",
         10712 => x"51ffb282",
         10713 => x"3f84b8e4",
         10714 => x"08839038",
         10715 => x"9c1708fe",
         10716 => x"11941908",
         10717 => x"58565b75",
         10718 => x"7527ffaf",
         10719 => x"38811694",
         10720 => x"180c8417",
         10721 => x"33810755",
         10722 => x"74841834",
         10723 => x"7c557a7d",
         10724 => x"26ffa038",
         10725 => x"80d93980",
         10726 => x"0b941734",
         10727 => x"800b9517",
         10728 => x"34fbcc39",
         10729 => x"95163394",
         10730 => x"17337198",
         10731 => x"2b71902b",
         10732 => x"077e075e",
         10733 => x"565b800b",
         10734 => x"8e173480",
         10735 => x"0b8f1734",
         10736 => x"a10b9017",
         10737 => x"3480cc0b",
         10738 => x"91173466",
         10739 => x"56a00b8b",
         10740 => x"17347e67",
         10741 => x"575e800b",
         10742 => x"9a173480",
         10743 => x"0b9b1734",
         10744 => x"7d335d7c",
         10745 => x"832e0981",
         10746 => x"06fb8438",
         10747 => x"ffa93980",
         10748 => x"7f7f725e",
         10749 => x"59575db4",
         10750 => x"16087e2e",
         10751 => x"ae388316",
         10752 => x"335a797d",
         10753 => x"2e098106",
         10754 => x"b5388154",
         10755 => x"7d53b816",
         10756 => x"52811633",
         10757 => x"51ffa3ba",
         10758 => x"3f84b8e4",
         10759 => x"08802e85",
         10760 => x"38ff5781",
         10761 => x"5b76b417",
         10762 => x"0c7e567a",
         10763 => x"ff1d9018",
         10764 => x"0c577a80",
         10765 => x"2efbbc38",
         10766 => x"80790cf9",
         10767 => x"97398154",
         10768 => x"b4160853",
         10769 => x"b8167053",
         10770 => x"81173352",
         10771 => x"5affa481",
         10772 => x"3f84b8e4",
         10773 => x"087d2e09",
         10774 => x"810681aa",
         10775 => x"3884b8e4",
         10776 => x"08831734",
         10777 => x"b41608a8",
         10778 => x"17083184",
         10779 => x"b8e4085c",
         10780 => x"5574a017",
         10781 => x"0827ff92",
         10782 => x"38821633",
         10783 => x"5574822e",
         10784 => x"098106ff",
         10785 => x"85388154",
         10786 => x"b41608a0",
         10787 => x"17080553",
         10788 => x"79528116",
         10789 => x"3351ffa3",
         10790 => x"b83f7c5b",
         10791 => x"feec3974",
         10792 => x"941a0c76",
         10793 => x"56f8af39",
         10794 => x"77981a0c",
         10795 => x"76f8a238",
         10796 => x"7583ff06",
         10797 => x"5a79802e",
         10798 => x"f89a387e",
         10799 => x"fe199c12",
         10800 => x"08fe055f",
         10801 => x"595a777d",
         10802 => x"27f9df38",
         10803 => x"8a1a2278",
         10804 => x"7129b01c",
         10805 => x"0805565c",
         10806 => x"74802ef9",
         10807 => x"cd387589",
         10808 => x"2a159c1a",
         10809 => x"0c7656f7",
         10810 => x"ed397594",
         10811 => x"1a0c7656",
         10812 => x"f7e43981",
         10813 => x"5780790c",
         10814 => x"f7da3984",
         10815 => x"b8e40857",
         10816 => x"80790cf7",
         10817 => x"cf39817f",
         10818 => x"575bfe9f",
         10819 => x"39f03d0d",
         10820 => x"62656766",
         10821 => x"40405d5a",
         10822 => x"807e0c89",
         10823 => x"5779802e",
         10824 => x"9f387908",
         10825 => x"5675802e",
         10826 => x"97387533",
         10827 => x"5574802e",
         10828 => x"8f388616",
         10829 => x"22841b22",
         10830 => x"59597878",
         10831 => x"2e84b738",
         10832 => x"80557441",
         10833 => x"76557682",
         10834 => x"8c38911a",
         10835 => x"33557482",
         10836 => x"8438901a",
         10837 => x"33810657",
         10838 => x"87567680",
         10839 => x"2e81ed38",
         10840 => x"941a088c",
         10841 => x"1b087131",
         10842 => x"56567b75",
         10843 => x"2681ef38",
         10844 => x"7b802e81",
         10845 => x"d5386059",
         10846 => x"7583ff06",
         10847 => x"5b7a81e3",
         10848 => x"388a1922",
         10849 => x"ff057689",
         10850 => x"2a065b7a",
         10851 => x"9b387583",
         10852 => x"d338881a",
         10853 => x"08558175",
         10854 => x"27848538",
         10855 => x"74ff2e83",
         10856 => x"f0387498",
         10857 => x"1b0c6059",
         10858 => x"981a08fe",
         10859 => x"059c1a08",
         10860 => x"fe054157",
         10861 => x"76602783",
         10862 => x"e7388a19",
         10863 => x"22707829",
         10864 => x"b01b0805",
         10865 => x"56567480",
         10866 => x"2e83d538",
         10867 => x"7a157c89",
         10868 => x"2a595777",
         10869 => x"802e8381",
         10870 => x"38771b55",
         10871 => x"75752785",
         10872 => x"38757b31",
         10873 => x"58775476",
         10874 => x"537c5281",
         10875 => x"193351ff",
         10876 => x"9fe03f84",
         10877 => x"b8e40883",
         10878 => x"98386083",
         10879 => x"11335759",
         10880 => x"75802ea9",
         10881 => x"38b41908",
         10882 => x"77315675",
         10883 => x"78279e38",
         10884 => x"84807671",
         10885 => x"291eb81b",
         10886 => x"58585575",
         10887 => x"70810557",
         10888 => x"33777081",
         10889 => x"055934ff",
         10890 => x"155574ef",
         10891 => x"3877892b",
         10892 => x"587b7831",
         10893 => x"7e08197f",
         10894 => x"0c781e94",
         10895 => x"1c081a70",
         10896 => x"59941d0c",
         10897 => x"5e5c7bfe",
         10898 => x"af388056",
         10899 => x"7584b8e4",
         10900 => x"0c923d0d",
         10901 => x"047484b8",
         10902 => x"e40c923d",
         10903 => x"0d04745c",
         10904 => x"fe8e399c",
         10905 => x"1a085775",
         10906 => x"83ff0684",
         10907 => x"80713159",
         10908 => x"5b7b7827",
         10909 => x"83387b58",
         10910 => x"7656b419",
         10911 => x"08772eb6",
         10912 => x"38800b83",
         10913 => x"1a33715d",
         10914 => x"415f7f7f",
         10915 => x"2e098106",
         10916 => x"80e43881",
         10917 => x"547653b8",
         10918 => x"19528119",
         10919 => x"3351ff9e",
         10920 => x"b13f84b8",
         10921 => x"e408802e",
         10922 => x"8538ff56",
         10923 => x"815b75b4",
         10924 => x"1a0c7a81",
         10925 => x"dc386094",
         10926 => x"1b0883ff",
         10927 => x"0611797f",
         10928 => x"5a58b805",
         10929 => x"56597780",
         10930 => x"2efee638",
         10931 => x"74708105",
         10932 => x"56337770",
         10933 => x"81055934",
         10934 => x"ff165675",
         10935 => x"802efed1",
         10936 => x"38747081",
         10937 => x"05563377",
         10938 => x"70810559",
         10939 => x"34ff1656",
         10940 => x"75da38fe",
         10941 => x"bc398154",
         10942 => x"b4190853",
         10943 => x"b8197053",
         10944 => x"811a3352",
         10945 => x"40ff9ec9",
         10946 => x"3f815b84",
         10947 => x"b8e4087f",
         10948 => x"2e098106",
         10949 => x"ff9c3884",
         10950 => x"b8e40883",
         10951 => x"1a34b419",
         10952 => x"08a81a08",
         10953 => x"3184b8e4",
         10954 => x"085c5574",
         10955 => x"a01a0827",
         10956 => x"fee13882",
         10957 => x"19335574",
         10958 => x"822e0981",
         10959 => x"06fed438",
         10960 => x"8154b419",
         10961 => x"08a01a08",
         10962 => x"05537f52",
         10963 => x"81193351",
         10964 => x"ff9dfe3f",
         10965 => x"7e5bfebb",
         10966 => x"39769c1b",
         10967 => x"0c941a08",
         10968 => x"56fe8439",
         10969 => x"981a0852",
         10970 => x"7951ffa3",
         10971 => x"983f84b8",
         10972 => x"e40855fc",
         10973 => x"a1398116",
         10974 => x"3351ff9c",
         10975 => x"833f84b8",
         10976 => x"e4088106",
         10977 => x"5574fbb8",
         10978 => x"38747a08",
         10979 => x"5657fbb2",
         10980 => x"39810b91",
         10981 => x"1b34810b",
         10982 => x"84b8e40c",
         10983 => x"923d0d04",
         10984 => x"820b911b",
         10985 => x"34820b84",
         10986 => x"b8e40c92",
         10987 => x"3d0d04f0",
         10988 => x"3d0d6265",
         10989 => x"67664040",
         10990 => x"5c5a807e",
         10991 => x"0c895779",
         10992 => x"802e9f38",
         10993 => x"79085675",
         10994 => x"802e9738",
         10995 => x"75335574",
         10996 => x"802e8f38",
         10997 => x"86162284",
         10998 => x"1b225959",
         10999 => x"78782e85",
         11000 => x"fd388055",
         11001 => x"74417655",
         11002 => x"7682c438",
         11003 => x"911a3355",
         11004 => x"7482bc38",
         11005 => x"901a3370",
         11006 => x"812a8106",
         11007 => x"58588756",
         11008 => x"76802e82",
         11009 => x"a138941a",
         11010 => x"087b115d",
         11011 => x"577b7727",
         11012 => x"84387609",
         11013 => x"5b7a802e",
         11014 => x"82813876",
         11015 => x"83ff065f",
         11016 => x"7e82a238",
         11017 => x"608a1122",
         11018 => x"ff057889",
         11019 => x"2a065a56",
         11020 => x"78aa3876",
         11021 => x"849e3888",
         11022 => x"1a085574",
         11023 => x"802e84b1",
         11024 => x"3874812e",
         11025 => x"86a13874",
         11026 => x"ff2e868c",
         11027 => x"3874981b",
         11028 => x"0c881a08",
         11029 => x"85387488",
         11030 => x"1b0c6056",
         11031 => x"b416089c",
         11032 => x"1b082e81",
         11033 => x"d338981a",
         11034 => x"08fe059c",
         11035 => x"1708fe05",
         11036 => x"58587777",
         11037 => x"2785f038",
         11038 => x"8a162270",
         11039 => x"7929b018",
         11040 => x"08055657",
         11041 => x"74802e85",
         11042 => x"de387815",
         11043 => x"7b892a59",
         11044 => x"5c77802e",
         11045 => x"83983877",
         11046 => x"195f767f",
         11047 => x"27853876",
         11048 => x"79315877",
         11049 => x"547b537c",
         11050 => x"52811633",
         11051 => x"51ff9ba1",
         11052 => x"3f84b8e4",
         11053 => x"0885a138",
         11054 => x"60b41108",
         11055 => x"7d315657",
         11056 => x"747827a5",
         11057 => x"3884800b",
         11058 => x"b8187672",
         11059 => x"291f5758",
         11060 => x"56747081",
         11061 => x"05563377",
         11062 => x"70810559",
         11063 => x"34ff1656",
         11064 => x"75ef3860",
         11065 => x"5975831a",
         11066 => x"3477892b",
         11067 => x"597a7931",
         11068 => x"7e081a7f",
         11069 => x"0c791e94",
         11070 => x"1c081b70",
         11071 => x"71941f0c",
         11072 => x"8c1e085a",
         11073 => x"5a575e5b",
         11074 => x"75752783",
         11075 => x"38745675",
         11076 => x"8c1b0c7a",
         11077 => x"fe853890",
         11078 => x"1a335877",
         11079 => x"80c0075b",
         11080 => x"7a901b34",
         11081 => x"80567584",
         11082 => x"b8e40c92",
         11083 => x"3d0d0474",
         11084 => x"84b8e40c",
         11085 => x"923d0d04",
         11086 => x"83163355",
         11087 => x"7482c838",
         11088 => x"6056fea2",
         11089 => x"39609c1b",
         11090 => x"08595676",
         11091 => x"83ff0684",
         11092 => x"8071315a",
         11093 => x"5c7a7927",
         11094 => x"83387a59",
         11095 => x"7757b416",
         11096 => x"08782eb6",
         11097 => x"38800b83",
         11098 => x"1733715e",
         11099 => x"415f7f7f",
         11100 => x"2e098106",
         11101 => x"80d53881",
         11102 => x"547753b8",
         11103 => x"16528116",
         11104 => x"3351ff98",
         11105 => x"cd3f84b8",
         11106 => x"e408802e",
         11107 => x"8538ff57",
         11108 => x"815c76b4",
         11109 => x"170c7b83",
         11110 => x"bf386094",
         11111 => x"1b0883ff",
         11112 => x"06117a58",
         11113 => x"b8057e59",
         11114 => x"56587880",
         11115 => x"2e953876",
         11116 => x"70810558",
         11117 => x"33757081",
         11118 => x"055734ff",
         11119 => x"165675ef",
         11120 => x"38605881",
         11121 => x"0b831934",
         11122 => x"fea33981",
         11123 => x"54b41608",
         11124 => x"53b81670",
         11125 => x"53811733",
         11126 => x"5240ff98",
         11127 => x"f43f815c",
         11128 => x"84b8e408",
         11129 => x"7f2e0981",
         11130 => x"06ffab38",
         11131 => x"84b8e408",
         11132 => x"831734b4",
         11133 => x"1608a817",
         11134 => x"083184b8",
         11135 => x"e4085d55",
         11136 => x"74a01708",
         11137 => x"27fef038",
         11138 => x"82163355",
         11139 => x"74822e09",
         11140 => x"8106fee3",
         11141 => x"388154b4",
         11142 => x"1608a017",
         11143 => x"0805537f",
         11144 => x"52811633",
         11145 => x"51ff98a9",
         11146 => x"3f7e5cfe",
         11147 => x"ca39941a",
         11148 => x"08578c1a",
         11149 => x"08772693",
         11150 => x"38831633",
         11151 => x"407f81b9",
         11152 => x"38607cb4",
         11153 => x"120c941b",
         11154 => x"0858567b",
         11155 => x"7c9c1c0c",
         11156 => x"58fdf839",
         11157 => x"981a0852",
         11158 => x"7951ffab",
         11159 => x"e73f84b8",
         11160 => x"e4085584",
         11161 => x"b8e408fb",
         11162 => x"d838901a",
         11163 => x"3358fdab",
         11164 => x"39765279",
         11165 => x"51ffabcc",
         11166 => x"3f84b8e4",
         11167 => x"085584b8",
         11168 => x"e408fbbd",
         11169 => x"38e43981",
         11170 => x"54b41608",
         11171 => x"53b81670",
         11172 => x"53811733",
         11173 => x"5257ff97",
         11174 => x"b83f84b8",
         11175 => x"e40881b8",
         11176 => x"3884b8e4",
         11177 => x"08831734",
         11178 => x"b41608a8",
         11179 => x"17083158",
         11180 => x"77a01708",
         11181 => x"27fd8938",
         11182 => x"8216335c",
         11183 => x"7b822e09",
         11184 => x"8106fcfc",
         11185 => x"388154b4",
         11186 => x"1608a017",
         11187 => x"08055376",
         11188 => x"52811633",
         11189 => x"51ff96f9",
         11190 => x"3f6056fb",
         11191 => x"89398116",
         11192 => x"3351ff95",
         11193 => x"9b3f84b8",
         11194 => x"e4088106",
         11195 => x"5574f9f2",
         11196 => x"38747a08",
         11197 => x"5657f9ec",
         11198 => x"398154b4",
         11199 => x"160853b8",
         11200 => x"16705381",
         11201 => x"17335257",
         11202 => x"ff96c63f",
         11203 => x"84b8e408",
         11204 => x"80c63884",
         11205 => x"b8e40883",
         11206 => x"1734b416",
         11207 => x"08a81708",
         11208 => x"315574a0",
         11209 => x"170827fe",
         11210 => x"98388216",
         11211 => x"33587782",
         11212 => x"2e098106",
         11213 => x"fe8b3881",
         11214 => x"54b41608",
         11215 => x"a0170805",
         11216 => x"53765281",
         11217 => x"163351ff",
         11218 => x"96873f60",
         11219 => x"7cb4120c",
         11220 => x"941b0858",
         11221 => x"56fdf439",
         11222 => x"810b911b",
         11223 => x"34810b84",
         11224 => x"b8e40c92",
         11225 => x"3d0d0482",
         11226 => x"0b911b34",
         11227 => x"820b84b8",
         11228 => x"e40c923d",
         11229 => x"0d04f53d",
         11230 => x"0d7d5889",
         11231 => x"5a77802e",
         11232 => x"9f387708",
         11233 => x"5675802e",
         11234 => x"97387533",
         11235 => x"5574802e",
         11236 => x"8f388616",
         11237 => x"22841922",
         11238 => x"58597877",
         11239 => x"2e83b538",
         11240 => x"8055745c",
         11241 => x"79567981",
         11242 => x"d8389018",
         11243 => x"3370862a",
         11244 => x"81065c57",
         11245 => x"7a802e81",
         11246 => x"c8387ba0",
         11247 => x"19085a57",
         11248 => x"b4170879",
         11249 => x"2eac3883",
         11250 => x"17335b7a",
         11251 => x"81bc3881",
         11252 => x"547853b8",
         11253 => x"17528117",
         11254 => x"3351ff93",
         11255 => x"f53f84b8",
         11256 => x"e408802e",
         11257 => x"8538ff59",
         11258 => x"815678b4",
         11259 => x"180c7581",
         11260 => x"9038a418",
         11261 => x"088b1133",
         11262 => x"a0075a57",
         11263 => x"788b1834",
         11264 => x"77088819",
         11265 => x"087083ff",
         11266 => x"ff065d5a",
         11267 => x"567a9a18",
         11268 => x"347a882a",
         11269 => x"5a799b18",
         11270 => x"349c1776",
         11271 => x"3396195c",
         11272 => x"565b7483",
         11273 => x"2e81c138",
         11274 => x"8c180855",
         11275 => x"747b3474",
         11276 => x"882a5b7a",
         11277 => x"9d183474",
         11278 => x"902a5675",
         11279 => x"9e183474",
         11280 => x"982a5978",
         11281 => x"9f183480",
         11282 => x"7a34800b",
         11283 => x"971834a1",
         11284 => x"0b981834",
         11285 => x"80cc0b99",
         11286 => x"1834800b",
         11287 => x"92183480",
         11288 => x"0b931834",
         11289 => x"7b5b810b",
         11290 => x"831c347b",
         11291 => x"51ff9694",
         11292 => x"3f84b8e4",
         11293 => x"08901933",
         11294 => x"81bf065b",
         11295 => x"56799019",
         11296 => x"347584b8",
         11297 => x"e40c8d3d",
         11298 => x"0d048154",
         11299 => x"b4170853",
         11300 => x"b8177053",
         11301 => x"81183352",
         11302 => x"5bff93b5",
         11303 => x"3f815684",
         11304 => x"b8e408fe",
         11305 => x"c93884b8",
         11306 => x"e4088318",
         11307 => x"34b41708",
         11308 => x"a8180831",
         11309 => x"84b8e408",
         11310 => x"575574a0",
         11311 => x"180827fe",
         11312 => x"8e388217",
         11313 => x"33557482",
         11314 => x"2e098106",
         11315 => x"fe813881",
         11316 => x"54b41708",
         11317 => x"a0180805",
         11318 => x"537a5281",
         11319 => x"173351ff",
         11320 => x"92ef3f79",
         11321 => x"56fde839",
         11322 => x"78902a55",
         11323 => x"74941834",
         11324 => x"74882a56",
         11325 => x"75951834",
         11326 => x"8c180855",
         11327 => x"747b3474",
         11328 => x"882a5b7a",
         11329 => x"9d183474",
         11330 => x"902a5675",
         11331 => x"9e183474",
         11332 => x"982a5978",
         11333 => x"9f183480",
         11334 => x"7a34800b",
         11335 => x"971834a1",
         11336 => x"0b981834",
         11337 => x"80cc0b99",
         11338 => x"1834800b",
         11339 => x"92183480",
         11340 => x"0b931834",
         11341 => x"7b5b810b",
         11342 => x"831c347b",
         11343 => x"51ff94c4",
         11344 => x"3f84b8e4",
         11345 => x"08901933",
         11346 => x"81bf065b",
         11347 => x"56799019",
         11348 => x"34feae39",
         11349 => x"81163351",
         11350 => x"ff90a53f",
         11351 => x"84b8e408",
         11352 => x"81065574",
         11353 => x"fcba3874",
         11354 => x"7808565a",
         11355 => x"fcb439f9",
         11356 => x"3d0d7970",
         11357 => x"5255fbfe",
         11358 => x"3f84b8e4",
         11359 => x"085484b8",
         11360 => x"e408b138",
         11361 => x"89567480",
         11362 => x"2e9e3874",
         11363 => x"08537280",
         11364 => x"2e963872",
         11365 => x"33527180",
         11366 => x"2e8e3886",
         11367 => x"13228416",
         11368 => x"22585271",
         11369 => x"772e9638",
         11370 => x"80527158",
         11371 => x"75547584",
         11372 => x"3875750c",
         11373 => x"7384b8e4",
         11374 => x"0c893d0d",
         11375 => x"04811333",
         11376 => x"51ff8fbc",
         11377 => x"3f84b8e4",
         11378 => x"08810653",
         11379 => x"72da3873",
         11380 => x"75085356",
         11381 => x"d539f63d",
         11382 => x"0dff7d70",
         11383 => x"5b575b75",
         11384 => x"802eb238",
         11385 => x"75708105",
         11386 => x"5733709f",
         11387 => x"26525271",
         11388 => x"ba2eac38",
         11389 => x"70ee3871",
         11390 => x"ba2ea438",
         11391 => x"84d0c033",
         11392 => x"51807124",
         11393 => x"90387084",
         11394 => x"d0c03480",
         11395 => x"0b84b8e4",
         11396 => x"0c8c3d0d",
         11397 => x"048b0b84",
         11398 => x"b8e40c8c",
         11399 => x"3d0d0478",
         11400 => x"33d01170",
         11401 => x"81ff0653",
         11402 => x"53537089",
         11403 => x"26913882",
         11404 => x"197381ff",
         11405 => x"06d00559",
         11406 => x"5473762e",
         11407 => x"80f53880",
         11408 => x"0b83e4d4",
         11409 => x"5b587908",
         11410 => x"79565776",
         11411 => x"70810558",
         11412 => x"33757081",
         11413 => x"055733ff",
         11414 => x"9f125354",
         11415 => x"52709926",
         11416 => x"8938e012",
         11417 => x"7081ff06",
         11418 => x"5354ff9f",
         11419 => x"13517099",
         11420 => x"268938e0",
         11421 => x"137081ff",
         11422 => x"06545471",
         11423 => x"30709f2a",
         11424 => x"55517173",
         11425 => x"2e098106",
         11426 => x"853873ff",
         11427 => x"be387476",
         11428 => x"32703070",
         11429 => x"72079f2a",
         11430 => x"76075952",
         11431 => x"5276802e",
         11432 => x"92388118",
         11433 => x"841b5b58",
         11434 => x"837825ff",
         11435 => x"99387a51",
         11436 => x"fecf3977",
         11437 => x"8324f738",
         11438 => x"77765e51",
         11439 => x"fec339ea",
         11440 => x"3d0d8053",
         11441 => x"983dcc05",
         11442 => x"52993d51",
         11443 => x"d1943f84",
         11444 => x"b8e40855",
         11445 => x"84b8e408",
         11446 => x"802e8a38",
         11447 => x"7484b8e4",
         11448 => x"0c983d0d",
         11449 => x"047a5c68",
         11450 => x"52983dd0",
         11451 => x"0551c594",
         11452 => x"3f84b8e4",
         11453 => x"085584b8",
         11454 => x"e40880c6",
         11455 => x"380280d7",
         11456 => x"05337098",
         11457 => x"2b585a80",
         11458 => x"772480e2",
         11459 => x"3802b205",
         11460 => x"3370842a",
         11461 => x"81065759",
         11462 => x"75802eb2",
         11463 => x"387a639b",
         11464 => x"11339a12",
         11465 => x"3371882b",
         11466 => x"0773335e",
         11467 => x"5a5b5758",
         11468 => x"79832ea4",
         11469 => x"38769819",
         11470 => x"0c7484b8",
         11471 => x"e40c983d",
         11472 => x"0d0484b8",
         11473 => x"e408842e",
         11474 => x"098106ff",
         11475 => x"8f38850b",
         11476 => x"84b8e40c",
         11477 => x"983d0d04",
         11478 => x"95163394",
         11479 => x"17337198",
         11480 => x"2b71902b",
         11481 => x"07790798",
         11482 => x"1b0c5b54",
         11483 => x"cc397a7e",
         11484 => x"98120c58",
         11485 => x"7484b8e4",
         11486 => x"0c983d0d",
         11487 => x"04ff9e3d",
         11488 => x"0d80e63d",
         11489 => x"0880e63d",
         11490 => x"085d4080",
         11491 => x"7c348053",
         11492 => x"80e43dfd",
         11493 => x"b4055280",
         11494 => x"e53d51cf",
         11495 => x"c53f84b8",
         11496 => x"e4085984",
         11497 => x"b8e40883",
         11498 => x"c8386080",
         11499 => x"d93d0c7f",
         11500 => x"61981108",
         11501 => x"80dd3d0c",
         11502 => x"5880db3d",
         11503 => x"085b5879",
         11504 => x"802e82cc",
         11505 => x"3880d83d",
         11506 => x"983d405b",
         11507 => x"a0527a51",
         11508 => x"ffa4aa3f",
         11509 => x"84b8e408",
         11510 => x"5984b8e4",
         11511 => x"08839238",
         11512 => x"6080df3d",
         11513 => x"085856b4",
         11514 => x"1608772e",
         11515 => x"b13884b8",
         11516 => x"e4088317",
         11517 => x"335f5d7d",
         11518 => x"83c73881",
         11519 => x"547653b8",
         11520 => x"16528116",
         11521 => x"3351ff8b",
         11522 => x"c93f84b8",
         11523 => x"e408802e",
         11524 => x"8538ff57",
         11525 => x"815976b4",
         11526 => x"170c7882",
         11527 => x"d43880df",
         11528 => x"3d089b11",
         11529 => x"339a1233",
         11530 => x"71882b07",
         11531 => x"6370335d",
         11532 => x"40595656",
         11533 => x"78832e82",
         11534 => x"da387680",
         11535 => x"db3d0c80",
         11536 => x"527a51ff",
         11537 => x"a3b73f84",
         11538 => x"b8e40859",
         11539 => x"84b8e408",
         11540 => x"829f3880",
         11541 => x"527a51ff",
         11542 => x"a8f53f84",
         11543 => x"b8e40859",
         11544 => x"84b8e408",
         11545 => x"bb3880df",
         11546 => x"3d089b11",
         11547 => x"339a1233",
         11548 => x"71882b07",
         11549 => x"63703342",
         11550 => x"58595e56",
         11551 => x"7d832e81",
         11552 => x"fd38767a",
         11553 => x"2ea43884",
         11554 => x"b8e40852",
         11555 => x"7a51ffa4",
         11556 => x"e23f84b8",
         11557 => x"e4085984",
         11558 => x"b8e40880",
         11559 => x"2effb438",
         11560 => x"78842e83",
         11561 => x"d8387881",
         11562 => x"c83880e4",
         11563 => x"3dfdb805",
         11564 => x"527a51ff",
         11565 => x"bd893f78",
         11566 => x"7f820533",
         11567 => x"5b577980",
         11568 => x"2e903882",
         11569 => x"1f568117",
         11570 => x"81177033",
         11571 => x"5f57577c",
         11572 => x"f5388117",
         11573 => x"56757826",
         11574 => x"81953876",
         11575 => x"802e9c38",
         11576 => x"7e178205",
         11577 => x"56ff1880",
         11578 => x"e63d0811",
         11579 => x"ff19ff19",
         11580 => x"59595658",
         11581 => x"75337534",
         11582 => x"76eb38ff",
         11583 => x"1880e63d",
         11584 => x"08115f58",
         11585 => x"af7e3480",
         11586 => x"da3d085a",
         11587 => x"79fdbd38",
         11588 => x"77602e82",
         11589 => x"8a38800b",
         11590 => x"84d0c033",
         11591 => x"70101083",
         11592 => x"e4d40570",
         11593 => x"08703343",
         11594 => x"59595e5a",
         11595 => x"7e7a2e8d",
         11596 => x"38811a70",
         11597 => x"17703357",
         11598 => x"5f5a74f5",
         11599 => x"38821a5b",
         11600 => x"7a7826ab",
         11601 => x"38805776",
         11602 => x"7a279438",
         11603 => x"76165f7e",
         11604 => x"337c7081",
         11605 => x"055e3481",
         11606 => x"17577977",
         11607 => x"26ee38ba",
         11608 => x"7c708105",
         11609 => x"5e3476ff",
         11610 => x"2e098106",
         11611 => x"81df3891",
         11612 => x"59807c34",
         11613 => x"7884b8e4",
         11614 => x"0c80e43d",
         11615 => x"0d049516",
         11616 => x"33941733",
         11617 => x"71982b71",
         11618 => x"902b0779",
         11619 => x"0759565e",
         11620 => x"fdf03995",
         11621 => x"16339417",
         11622 => x"3371982b",
         11623 => x"71902b07",
         11624 => x"790780dd",
         11625 => x"3d0c5a5d",
         11626 => x"80527a51",
         11627 => x"ffa0ce3f",
         11628 => x"84b8e408",
         11629 => x"5984b8e4",
         11630 => x"08802efd",
         11631 => x"9638ffb1",
         11632 => x"398154b4",
         11633 => x"160853b8",
         11634 => x"16705381",
         11635 => x"1733525e",
         11636 => x"ff88fe3f",
         11637 => x"815984b8",
         11638 => x"e408fcbe",
         11639 => x"3884b8e4",
         11640 => x"08831734",
         11641 => x"b41608a8",
         11642 => x"17083184",
         11643 => x"b8e4085a",
         11644 => x"5574a017",
         11645 => x"0827fc83",
         11646 => x"38821633",
         11647 => x"5574822e",
         11648 => x"098106fb",
         11649 => x"f6388154",
         11650 => x"b41608a0",
         11651 => x"17080553",
         11652 => x"7d528116",
         11653 => x"3351ff88",
         11654 => x"b83f7c59",
         11655 => x"fbdd39ff",
         11656 => x"1880e63d",
         11657 => x"08115c58",
         11658 => x"af7b3480",
         11659 => x"0b84d0c0",
         11660 => x"33701010",
         11661 => x"83e4d405",
         11662 => x"70087033",
         11663 => x"4359595e",
         11664 => x"5a7e7a2e",
         11665 => x"098106fd",
         11666 => x"e838fdf1",
         11667 => x"3980e53d",
         11668 => x"08188119",
         11669 => x"595a7933",
         11670 => x"7c708105",
         11671 => x"5e347760",
         11672 => x"27fe8e38",
         11673 => x"80e53d08",
         11674 => x"18811959",
         11675 => x"5a79337c",
         11676 => x"7081055e",
         11677 => x"347f7826",
         11678 => x"d438fdf5",
         11679 => x"39825980",
         11680 => x"7c347884",
         11681 => x"b8e40c80",
         11682 => x"e43d0d04",
         11683 => x"f73d0d7b",
         11684 => x"7d585589",
         11685 => x"5674802e",
         11686 => x"9f387408",
         11687 => x"5473802e",
         11688 => x"97387333",
         11689 => x"5372802e",
         11690 => x"8f388614",
         11691 => x"22841622",
         11692 => x"59597878",
         11693 => x"2e83a038",
         11694 => x"8053725a",
         11695 => x"75537581",
         11696 => x"c2389115",
         11697 => x"33537281",
         11698 => x"ba388c15",
         11699 => x"08567676",
         11700 => x"2681b938",
         11701 => x"94150854",
         11702 => x"80587678",
         11703 => x"2e81cc38",
         11704 => x"798a1122",
         11705 => x"70892b52",
         11706 => x"5a567378",
         11707 => x"2e81f738",
         11708 => x"7552ff17",
         11709 => x"51fdbbad",
         11710 => x"3f84b8e4",
         11711 => x"08ff1577",
         11712 => x"54705355",
         11713 => x"53fdbb9d",
         11714 => x"3f84b8e4",
         11715 => x"08732681",
         11716 => x"d5387530",
         11717 => x"74067094",
         11718 => x"170c7771",
         11719 => x"31981708",
         11720 => x"56585973",
         11721 => x"802e8298",
         11722 => x"38757727",
         11723 => x"81d93876",
         11724 => x"76319416",
         11725 => x"08179417",
         11726 => x"0c901633",
         11727 => x"70812a81",
         11728 => x"06515a57",
         11729 => x"78802e81",
         11730 => x"fe387352",
         11731 => x"7451ff99",
         11732 => x"f33f84b8",
         11733 => x"e4085484",
         11734 => x"b8e40880",
         11735 => x"2e81a338",
         11736 => x"73ff2e98",
         11737 => x"38817427",
         11738 => x"82b43879",
         11739 => x"53739c14",
         11740 => x"082782aa",
         11741 => x"38739816",
         11742 => x"0cffae39",
         11743 => x"810b9116",
         11744 => x"34815372",
         11745 => x"84b8e40c",
         11746 => x"8b3d0d04",
         11747 => x"90153370",
         11748 => x"812a8106",
         11749 => x"555873fe",
         11750 => x"bb387594",
         11751 => x"16085557",
         11752 => x"80587678",
         11753 => x"2e098106",
         11754 => x"feb63877",
         11755 => x"94160c94",
         11756 => x"15085475",
         11757 => x"74279038",
         11758 => x"738c160c",
         11759 => x"90153380",
         11760 => x"c0075776",
         11761 => x"90163473",
         11762 => x"83ff0659",
         11763 => x"78802e8c",
         11764 => x"389c1508",
         11765 => x"782e8538",
         11766 => x"779c160c",
         11767 => x"800b84b8",
         11768 => x"e40c8b3d",
         11769 => x"0d04800b",
         11770 => x"94160c88",
         11771 => x"15085473",
         11772 => x"802e80fe",
         11773 => x"38739816",
         11774 => x"0c73802e",
         11775 => x"80c238fe",
         11776 => x"a83984b8",
         11777 => x"e4085794",
         11778 => x"15081794",
         11779 => x"160c7683",
         11780 => x"ff065675",
         11781 => x"802ea938",
         11782 => x"79fe159c",
         11783 => x"1208fe05",
         11784 => x"5a555673",
         11785 => x"782780f6",
         11786 => x"388a1622",
         11787 => x"747129b0",
         11788 => x"18080578",
         11789 => x"892a115a",
         11790 => x"5a537880",
         11791 => x"2e80df38",
         11792 => x"8c150856",
         11793 => x"fee93973",
         11794 => x"527451ff",
         11795 => x"89b73f84",
         11796 => x"b8e40854",
         11797 => x"fe8a3981",
         11798 => x"143351ff",
         11799 => x"82a23f84",
         11800 => x"b8e40881",
         11801 => x"065372fc",
         11802 => x"cf387275",
         11803 => x"085456fc",
         11804 => x"c9397352",
         11805 => x"7451ff97",
         11806 => x"cb3f84b8",
         11807 => x"e4085484",
         11808 => x"b8e40881",
         11809 => x"2e983884",
         11810 => x"b8e408ff",
         11811 => x"2efded38",
         11812 => x"84b8e408",
         11813 => x"88160c73",
         11814 => x"98160cfe",
         11815 => x"dc39820b",
         11816 => x"91163482",
         11817 => x"0b84b8e4",
         11818 => x"0c8b3d0d",
         11819 => x"04f63d0d",
         11820 => x"7c568954",
         11821 => x"75802ea2",
         11822 => x"3880538c",
         11823 => x"3dfc0552",
         11824 => x"8d3d8405",
         11825 => x"51c59b3f",
         11826 => x"84b8e408",
         11827 => x"5584b8e4",
         11828 => x"08802e8f",
         11829 => x"3880760c",
         11830 => x"74547384",
         11831 => x"b8e40c8c",
         11832 => x"3d0d047a",
         11833 => x"760c7d52",
         11834 => x"7551ffb9",
         11835 => x"973f84b8",
         11836 => x"e4085584",
         11837 => x"b8e40880",
         11838 => x"d138ab16",
         11839 => x"3370982b",
         11840 => x"59598078",
         11841 => x"24af3886",
         11842 => x"16337084",
         11843 => x"2a81065b",
         11844 => x"5479802e",
         11845 => x"80c5389c",
         11846 => x"16089b11",
         11847 => x"339a1233",
         11848 => x"71882b07",
         11849 => x"7d70335d",
         11850 => x"5d5a5557",
         11851 => x"78832eb3",
         11852 => x"38778817",
         11853 => x"0c7a5886",
         11854 => x"18228417",
         11855 => x"23745275",
         11856 => x"51ff99b9",
         11857 => x"3f84b8e4",
         11858 => x"08557484",
         11859 => x"2e8d3874",
         11860 => x"802eff84",
         11861 => x"3880760c",
         11862 => x"fefe3985",
         11863 => x"5580760c",
         11864 => x"fef63995",
         11865 => x"17339418",
         11866 => x"3371982b",
         11867 => x"71902b07",
         11868 => x"7a078819",
         11869 => x"0c5a5aff",
         11870 => x"bc39fa3d",
         11871 => x"0d785589",
         11872 => x"5474802e",
         11873 => x"9e387408",
         11874 => x"5372802e",
         11875 => x"96387233",
         11876 => x"5271802e",
         11877 => x"8e388613",
         11878 => x"22841622",
         11879 => x"57527176",
         11880 => x"2e943880",
         11881 => x"52715773",
         11882 => x"84387375",
         11883 => x"0c7384b8",
         11884 => x"e40c883d",
         11885 => x"0d048113",
         11886 => x"3351feff",
         11887 => x"c33f84b8",
         11888 => x"e4088106",
         11889 => x"5271dc38",
         11890 => x"71750853",
         11891 => x"54d739f8",
         11892 => x"3d0d7a7c",
         11893 => x"58558956",
         11894 => x"74802e9f",
         11895 => x"38740854",
         11896 => x"73802e97",
         11897 => x"38733353",
         11898 => x"72802e8f",
         11899 => x"38861422",
         11900 => x"84162259",
         11901 => x"5372782e",
         11902 => x"81973880",
         11903 => x"53725975",
         11904 => x"537580c7",
         11905 => x"3876802e",
         11906 => x"80f33875",
         11907 => x"527451ff",
         11908 => x"9dbd3f84",
         11909 => x"b8e40853",
         11910 => x"84b8e408",
         11911 => x"842eb538",
         11912 => x"84b8e408",
         11913 => x"a6387652",
         11914 => x"7451ffb2",
         11915 => x"923f7252",
         11916 => x"7451ff99",
         11917 => x"be3f84b8",
         11918 => x"e4088432",
         11919 => x"70307072",
         11920 => x"079f2c84",
         11921 => x"b8e40806",
         11922 => x"55575472",
         11923 => x"84b8e40c",
         11924 => x"8a3d0d04",
         11925 => x"75775375",
         11926 => x"5253ffb1",
         11927 => x"e23f7252",
         11928 => x"7451ff99",
         11929 => x"8e3f84b8",
         11930 => x"e4088432",
         11931 => x"70307072",
         11932 => x"079f2c84",
         11933 => x"b8e40806",
         11934 => x"555754cf",
         11935 => x"39755274",
         11936 => x"51ff96f9",
         11937 => x"3f84b8e4",
         11938 => x"0884b8e4",
         11939 => x"0c8a3d0d",
         11940 => x"04811433",
         11941 => x"51fefde8",
         11942 => x"3f84b8e4",
         11943 => x"08810653",
         11944 => x"72fed838",
         11945 => x"72750854",
         11946 => x"56fed239",
         11947 => x"ed3d0d66",
         11948 => x"57805389",
         11949 => x"3d705397",
         11950 => x"3d5256c1",
         11951 => x"a53f84b8",
         11952 => x"e4085584",
         11953 => x"b8e40880",
         11954 => x"2e8a3874",
         11955 => x"84b8e40c",
         11956 => x"953d0d04",
         11957 => x"65527551",
         11958 => x"ffb5a93f",
         11959 => x"84b8e408",
         11960 => x"5584b8e4",
         11961 => x"08e53802",
         11962 => x"80cb0533",
         11963 => x"70982b55",
         11964 => x"58807424",
         11965 => x"97387680",
         11966 => x"2ed13876",
         11967 => x"527551ff",
         11968 => x"b0bd3f74",
         11969 => x"84b8e40c",
         11970 => x"953d0d04",
         11971 => x"860b84b8",
         11972 => x"e40c953d",
         11973 => x"0d04ed3d",
         11974 => x"0d666856",
         11975 => x"5f805395",
         11976 => x"3dec0552",
         11977 => x"963d51c0",
         11978 => x"b93f84b8",
         11979 => x"e4085a84",
         11980 => x"b8e4089a",
         11981 => x"387f750c",
         11982 => x"74089c11",
         11983 => x"08fe1194",
         11984 => x"13085957",
         11985 => x"59577575",
         11986 => x"268d3875",
         11987 => x"7f0c7984",
         11988 => x"b8e40c95",
         11989 => x"3d0d0484",
         11990 => x"b8e40877",
         11991 => x"335a5b78",
         11992 => x"812e8293",
         11993 => x"3877a818",
         11994 => x"0884b8e4",
         11995 => x"085a5d59",
         11996 => x"7780c138",
         11997 => x"7b811d71",
         11998 => x"5c5d56b4",
         11999 => x"1708762e",
         12000 => x"82ef3883",
         12001 => x"1733785f",
         12002 => x"5d7c818d",
         12003 => x"38815475",
         12004 => x"53b81752",
         12005 => x"81173351",
         12006 => x"fefcb73f",
         12007 => x"84b8e408",
         12008 => x"802e8538",
         12009 => x"ff5a815e",
         12010 => x"79b4180c",
         12011 => x"7f7e5b57",
         12012 => x"7d80cc38",
         12013 => x"76335e7d",
         12014 => x"822e828d",
         12015 => x"387717b8",
         12016 => x"05831133",
         12017 => x"82123371",
         12018 => x"902b7188",
         12019 => x"2b078114",
         12020 => x"33707207",
         12021 => x"882b7533",
         12022 => x"7180ffff",
         12023 => x"fe800607",
         12024 => x"70307080",
         12025 => x"25630560",
         12026 => x"840583ff",
         12027 => x"0662ff05",
         12028 => x"43414353",
         12029 => x"54525358",
         12030 => x"405e5678",
         12031 => x"fef2387a",
         12032 => x"7f0c7a94",
         12033 => x"180c8417",
         12034 => x"33810758",
         12035 => x"77841834",
         12036 => x"7984b8e4",
         12037 => x"0c953d0d",
         12038 => x"048154b4",
         12039 => x"170853b8",
         12040 => x"17705381",
         12041 => x"1833525d",
         12042 => x"fefca63f",
         12043 => x"815e84b8",
         12044 => x"e408fef8",
         12045 => x"3884b8e4",
         12046 => x"08831834",
         12047 => x"b41708a8",
         12048 => x"18083184",
         12049 => x"b8e4085f",
         12050 => x"5574a018",
         12051 => x"0827febd",
         12052 => x"38821733",
         12053 => x"5574822e",
         12054 => x"098106fe",
         12055 => x"b0388154",
         12056 => x"b41708a0",
         12057 => x"18080553",
         12058 => x"7c528117",
         12059 => x"3351fefb",
         12060 => x"e03f775e",
         12061 => x"fe973982",
         12062 => x"7742923d",
         12063 => x"59567552",
         12064 => x"7751ff81",
         12065 => x"803f84b8",
         12066 => x"e408ff2e",
         12067 => x"80e83884",
         12068 => x"b8e40881",
         12069 => x"2e80f738",
         12070 => x"84b8e408",
         12071 => x"307084b8",
         12072 => x"e4080780",
         12073 => x"257c0581",
         12074 => x"18625a58",
         12075 => x"5c5c9c17",
         12076 => x"087626ca",
         12077 => x"387a7f0c",
         12078 => x"7a94180c",
         12079 => x"84173381",
         12080 => x"07587784",
         12081 => x"1834fec8",
         12082 => x"397717b8",
         12083 => x"05811133",
         12084 => x"71337188",
         12085 => x"2b077030",
         12086 => x"7080251f",
         12087 => x"821d83ff",
         12088 => x"06ff1f5f",
         12089 => x"5d5f595f",
         12090 => x"5f5578fd",
         12091 => x"8338fe8f",
         12092 => x"39775afd",
         12093 => x"bf398160",
         12094 => x"585a7a7f",
         12095 => x"0c7a9418",
         12096 => x"0c841733",
         12097 => x"81075877",
         12098 => x"841834fe",
         12099 => x"83398260",
         12100 => x"585ae739",
         12101 => x"f73d0d7b",
         12102 => x"57895676",
         12103 => x"802e9f38",
         12104 => x"76085574",
         12105 => x"802e9738",
         12106 => x"74335473",
         12107 => x"802e8f38",
         12108 => x"86152284",
         12109 => x"18225959",
         12110 => x"78782e81",
         12111 => x"da388054",
         12112 => x"735a7580",
         12113 => x"dc389117",
         12114 => x"33567580",
         12115 => x"d4389017",
         12116 => x"3370812a",
         12117 => x"81065558",
         12118 => x"87557380",
         12119 => x"2e80c438",
         12120 => x"94170854",
         12121 => x"738c1808",
         12122 => x"27b73873",
         12123 => x"81d53888",
         12124 => x"17087708",
         12125 => x"57548174",
         12126 => x"2788389c",
         12127 => x"16087426",
         12128 => x"b3388256",
         12129 => x"800b8818",
         12130 => x"0c941708",
         12131 => x"8c180c77",
         12132 => x"80c00759",
         12133 => x"78901834",
         12134 => x"75802e85",
         12135 => x"38759118",
         12136 => x"34755574",
         12137 => x"84b8e40c",
         12138 => x"8b3d0d04",
         12139 => x"78547878",
         12140 => x"2780ff38",
         12141 => x"73527651",
         12142 => x"fefeca3f",
         12143 => x"84b8e408",
         12144 => x"5984b8e4",
         12145 => x"08802e80",
         12146 => x"e93884b8",
         12147 => x"e408812e",
         12148 => x"82d83884",
         12149 => x"b8e408ff",
         12150 => x"2e82e538",
         12151 => x"80537352",
         12152 => x"7551ff85",
         12153 => x"813f84b8",
         12154 => x"e40882c8",
         12155 => x"389c1608",
         12156 => x"fe119418",
         12157 => x"08575558",
         12158 => x"747427ff",
         12159 => x"af388115",
         12160 => x"94170c84",
         12161 => x"16338107",
         12162 => x"54738417",
         12163 => x"34785477",
         12164 => x"7926ffa0",
         12165 => x"389c3981",
         12166 => x"153351fe",
         12167 => x"f6e23f84",
         12168 => x"b8e40881",
         12169 => x"065473fe",
         12170 => x"95387377",
         12171 => x"085556fe",
         12172 => x"8f39800b",
         12173 => x"90183359",
         12174 => x"54735680",
         12175 => x"0b88180c",
         12176 => x"fec73998",
         12177 => x"17085276",
         12178 => x"51fefdb9",
         12179 => x"3f84b8e4",
         12180 => x"08ff2e81",
         12181 => x"c23884b8",
         12182 => x"e408812e",
         12183 => x"81be3875",
         12184 => x"81ae3879",
         12185 => x"5884b8e4",
         12186 => x"089c1908",
         12187 => x"2781a138",
         12188 => x"84b8e408",
         12189 => x"98180878",
         12190 => x"08585654",
         12191 => x"810b84b8",
         12192 => x"e4082781",
         12193 => x"a13884b8",
         12194 => x"e4089c17",
         12195 => x"08278196",
         12196 => x"3874802e",
         12197 => x"9738ff53",
         12198 => x"74527551",
         12199 => x"ff83c73f",
         12200 => x"84b8e408",
         12201 => x"5584b8e4",
         12202 => x"0880e338",
         12203 => x"73527651",
         12204 => x"fefcd23f",
         12205 => x"84b8e408",
         12206 => x"5984b8e4",
         12207 => x"08802e80",
         12208 => x"cb3884b8",
         12209 => x"e408812e",
         12210 => x"80dc3884",
         12211 => x"b8e408ff",
         12212 => x"2e80fe38",
         12213 => x"80537352",
         12214 => x"7551ff83",
         12215 => x"893f84b8",
         12216 => x"e40880e6",
         12217 => x"389c1608",
         12218 => x"fe119418",
         12219 => x"08575558",
         12220 => x"74742790",
         12221 => x"38811594",
         12222 => x"170c8416",
         12223 => x"33810754",
         12224 => x"73841734",
         12225 => x"78547779",
         12226 => x"26ffa138",
         12227 => x"80557456",
         12228 => x"90173358",
         12229 => x"fcf33981",
         12230 => x"56febb39",
         12231 => x"820b9018",
         12232 => x"335956fc",
         12233 => x"e4398256",
         12234 => x"e739820b",
         12235 => x"90183359",
         12236 => x"54fe8639",
         12237 => x"84b8e408",
         12238 => x"90183359",
         12239 => x"54fdfa39",
         12240 => x"810b9018",
         12241 => x"335954fd",
         12242 => x"f03984b8",
         12243 => x"e40856c0",
         12244 => x"398156ff",
         12245 => x"bb39db3d",
         12246 => x"0d8253a7",
         12247 => x"3dff9c05",
         12248 => x"52a83d51",
         12249 => x"ffb7fb3f",
         12250 => x"84b8e408",
         12251 => x"5684b8e4",
         12252 => x"08802e8a",
         12253 => x"387584b8",
         12254 => x"e40ca73d",
         12255 => x"0d047d4b",
         12256 => x"a83d0852",
         12257 => x"9b3d7052",
         12258 => x"59ffabf8",
         12259 => x"3f84b8e4",
         12260 => x"085684b8",
         12261 => x"e408de38",
         12262 => x"02819305",
         12263 => x"3370852a",
         12264 => x"81065957",
         12265 => x"865677cd",
         12266 => x"3876982b",
         12267 => x"5b807b24",
         12268 => x"c4380280",
         12269 => x"ee053370",
         12270 => x"81065d57",
         12271 => x"87567bff",
         12272 => x"b4387da3",
         12273 => x"3d089b11",
         12274 => x"339a1233",
         12275 => x"71882b07",
         12276 => x"7333415e",
         12277 => x"5c57587c",
         12278 => x"832e80d5",
         12279 => x"3876842a",
         12280 => x"81065776",
         12281 => x"802e80ed",
         12282 => x"38875698",
         12283 => x"18087b2e",
         12284 => x"ff833877",
         12285 => x"5f7a4184",
         12286 => x"b8e40852",
         12287 => x"8f3d7052",
         12288 => x"55ff8bf9",
         12289 => x"3f84b8e4",
         12290 => x"085684b8",
         12291 => x"e408fee5",
         12292 => x"3884b8e4",
         12293 => x"08527451",
         12294 => x"ff91b43f",
         12295 => x"84b8e408",
         12296 => x"5684b8e4",
         12297 => x"08a03887",
         12298 => x"0b84b8e4",
         12299 => x"0ca73d0d",
         12300 => x"04951633",
         12301 => x"94173371",
         12302 => x"982b7190",
         12303 => x"2b077d07",
         12304 => x"5d5d5dff",
         12305 => x"983984b8",
         12306 => x"e408842e",
         12307 => x"883884b8",
         12308 => x"e408fea1",
         12309 => x"3878086f",
         12310 => x"a83d0857",
         12311 => x"5d5774ff",
         12312 => x"2e80d338",
         12313 => x"74527851",
         12314 => x"ff8b923f",
         12315 => x"84b8e408",
         12316 => x"5684b8e4",
         12317 => x"08802ebe",
         12318 => x"38753070",
         12319 => x"77078025",
         12320 => x"565a7a80",
         12321 => x"2e9a3874",
         12322 => x"802e9538",
         12323 => x"7a790858",
         12324 => x"55817b27",
         12325 => x"89389c17",
         12326 => x"087b2681",
         12327 => x"fd388256",
         12328 => x"75fdd238",
         12329 => x"7d51fef5",
         12330 => x"db3f84b8",
         12331 => x"e40884b8",
         12332 => x"e40ca73d",
         12333 => x"0d04b817",
         12334 => x"5d981908",
         12335 => x"56805ab4",
         12336 => x"1708762e",
         12337 => x"82b93883",
         12338 => x"17337a59",
         12339 => x"55747a2e",
         12340 => x"09810680",
         12341 => x"dd388154",
         12342 => x"7553b817",
         12343 => x"52811733",
         12344 => x"51fef1ee",
         12345 => x"3f84b8e4",
         12346 => x"08802e85",
         12347 => x"38ff5681",
         12348 => x"5875b418",
         12349 => x"0c775677",
         12350 => x"ab389c19",
         12351 => x"0858e578",
         12352 => x"34810b83",
         12353 => x"18349019",
         12354 => x"087c27fe",
         12355 => x"ec388052",
         12356 => x"7851ff8b",
         12357 => x"de3f84b8",
         12358 => x"e4085684",
         12359 => x"b8e40880",
         12360 => x"2eff9638",
         12361 => x"75842e09",
         12362 => x"8106fecd",
         12363 => x"388256fe",
         12364 => x"c8398154",
         12365 => x"b4170853",
         12366 => x"7c528117",
         12367 => x"3351fef2",
         12368 => x"903f8158",
         12369 => x"84b8e408",
         12370 => x"7a2e0981",
         12371 => x"06ffa638",
         12372 => x"84b8e408",
         12373 => x"831834b4",
         12374 => x"1708a818",
         12375 => x"083184b8",
         12376 => x"e4085955",
         12377 => x"74a01808",
         12378 => x"27feeb38",
         12379 => x"82173355",
         12380 => x"74822e09",
         12381 => x"8106fede",
         12382 => x"388154b4",
         12383 => x"1708a018",
         12384 => x"0805537c",
         12385 => x"52811733",
         12386 => x"51fef1c5",
         12387 => x"3f7958fe",
         12388 => x"c5397955",
         12389 => x"79782780",
         12390 => x"e1387452",
         12391 => x"7851fef6",
         12392 => x"e43f84b8",
         12393 => x"e4085a84",
         12394 => x"b8e40880",
         12395 => x"2e80cb38",
         12396 => x"84b8e408",
         12397 => x"812efde6",
         12398 => x"3884b8e4",
         12399 => x"08ff2e80",
         12400 => x"cb388053",
         12401 => x"74527651",
         12402 => x"fefd9b3f",
         12403 => x"84b8e408",
         12404 => x"b3389c17",
         12405 => x"08fe1194",
         12406 => x"1908585c",
         12407 => x"58757b27",
         12408 => x"ffb03881",
         12409 => x"1694180c",
         12410 => x"84173381",
         12411 => x"075c7b84",
         12412 => x"18347955",
         12413 => x"777a26ff",
         12414 => x"a1388056",
         12415 => x"fda23979",
         12416 => x"56fdf739",
         12417 => x"84b8e408",
         12418 => x"56fd9539",
         12419 => x"8156fd90",
         12420 => x"39e33d0d",
         12421 => x"82539f3d",
         12422 => x"ffbc0552",
         12423 => x"a03d51ff",
         12424 => x"b2c03f84",
         12425 => x"b8e40856",
         12426 => x"84b8e408",
         12427 => x"802e8a38",
         12428 => x"7584b8e4",
         12429 => x"0c9f3d0d",
         12430 => x"047d436f",
         12431 => x"52933d70",
         12432 => x"525affa6",
         12433 => x"bf3f84b8",
         12434 => x"e4085684",
         12435 => x"b8e4088b",
         12436 => x"38880b84",
         12437 => x"b8e40c9f",
         12438 => x"3d0d0484",
         12439 => x"b8e40884",
         12440 => x"2e098106",
         12441 => x"cb380280",
         12442 => x"f3053370",
         12443 => x"852a8106",
         12444 => x"56588656",
         12445 => x"74ffb938",
         12446 => x"7d5f7452",
         12447 => x"8f3d7052",
         12448 => x"5dff83c0",
         12449 => x"3f84b8e4",
         12450 => x"0875575c",
         12451 => x"84b8e408",
         12452 => x"83388756",
         12453 => x"84b8e408",
         12454 => x"812e80f9",
         12455 => x"3884b8e4",
         12456 => x"08ff2e81",
         12457 => x"cb387581",
         12458 => x"c9387d84",
         12459 => x"b8e40883",
         12460 => x"12335d5a",
         12461 => x"577a80e2",
         12462 => x"38fe199c",
         12463 => x"1808fe05",
         12464 => x"5a56805b",
         12465 => x"7579278d",
         12466 => x"388a1722",
         12467 => x"767129b0",
         12468 => x"1908055c",
         12469 => x"587ab418",
         12470 => x"0cb81759",
         12471 => x"84807957",
         12472 => x"55807670",
         12473 => x"81055834",
         12474 => x"ff155574",
         12475 => x"f4387458",
         12476 => x"8a172255",
         12477 => x"77752781",
         12478 => x"f9388154",
         12479 => x"771b5378",
         12480 => x"52811733",
         12481 => x"51feeec9",
         12482 => x"3f84b8e4",
         12483 => x"0881df38",
         12484 => x"811858dc",
         12485 => x"398256ff",
         12486 => x"84398154",
         12487 => x"b4170853",
         12488 => x"b8177053",
         12489 => x"81183352",
         12490 => x"58feeea5",
         12491 => x"3f815684",
         12492 => x"b8e408be",
         12493 => x"3884b8e4",
         12494 => x"08831834",
         12495 => x"b41708a8",
         12496 => x"18083155",
         12497 => x"74a01808",
         12498 => x"27feee38",
         12499 => x"8217335b",
         12500 => x"7a822e09",
         12501 => x"8106fee1",
         12502 => x"387554b4",
         12503 => x"1708a018",
         12504 => x"08055377",
         12505 => x"52811733",
         12506 => x"51feede5",
         12507 => x"3ffeca39",
         12508 => x"81567b7d",
         12509 => x"08585581",
         12510 => x"7c27fdb4",
         12511 => x"387b9c18",
         12512 => x"0827fdac",
         12513 => x"3874527c",
         12514 => x"51fef2f9",
         12515 => x"3f84b8e4",
         12516 => x"085a84b8",
         12517 => x"e408802e",
         12518 => x"fd963884",
         12519 => x"b8e40881",
         12520 => x"2efd8d38",
         12521 => x"84b8e408",
         12522 => x"ff2efd84",
         12523 => x"38805374",
         12524 => x"527651fe",
         12525 => x"f9b03f84",
         12526 => x"b8e408fc",
         12527 => x"f3389c17",
         12528 => x"08fe1194",
         12529 => x"19085a5c",
         12530 => x"59777b27",
         12531 => x"90388118",
         12532 => x"94180c84",
         12533 => x"17338107",
         12534 => x"5c7b8418",
         12535 => x"34795578",
         12536 => x"7a26ffa1",
         12537 => x"387584b8",
         12538 => x"e40c9f3d",
         12539 => x"0d048a17",
         12540 => x"22557483",
         12541 => x"ffff0657",
         12542 => x"81567678",
         12543 => x"2e098106",
         12544 => x"fef0388b",
         12545 => x"0bb81f56",
         12546 => x"56a07570",
         12547 => x"81055734",
         12548 => x"ff165675",
         12549 => x"f4387d57",
         12550 => x"ae0bb818",
         12551 => x"347d5890",
         12552 => x"0b80c319",
         12553 => x"347d5975",
         12554 => x"80ce1a34",
         12555 => x"7580cf1a",
         12556 => x"34a10b80",
         12557 => x"d01a3480",
         12558 => x"cc0b80d1",
         12559 => x"1a347d7c",
         12560 => x"83ffff06",
         12561 => x"59567780",
         12562 => x"d2173477",
         12563 => x"882a5b7a",
         12564 => x"80d31734",
         12565 => x"75335574",
         12566 => x"832e81cc",
         12567 => x"387d59a0",
         12568 => x"0b80d81a",
         12569 => x"b81b5758",
         12570 => x"56747081",
         12571 => x"05563377",
         12572 => x"70810559",
         12573 => x"34ff1656",
         12574 => x"75ef387d",
         12575 => x"56ae0b80",
         12576 => x"d9173464",
         12577 => x"7e7183ff",
         12578 => x"ff065b57",
         12579 => x"577880f2",
         12580 => x"17347888",
         12581 => x"2a5b7a80",
         12582 => x"f3173475",
         12583 => x"33557483",
         12584 => x"2e80f038",
         12585 => x"7d5b810b",
         12586 => x"831c3479",
         12587 => x"51ff9296",
         12588 => x"3f84b8e4",
         12589 => x"085684b8",
         12590 => x"e408fdb6",
         12591 => x"38695684",
         12592 => x"b8e40896",
         12593 => x"173484b8",
         12594 => x"e4089717",
         12595 => x"34a10b98",
         12596 => x"173480cc",
         12597 => x"0b991734",
         12598 => x"7d6a585d",
         12599 => x"779a1834",
         12600 => x"77882a59",
         12601 => x"789b1834",
         12602 => x"7c335a79",
         12603 => x"832e80d9",
         12604 => x"38695590",
         12605 => x"0b8b1634",
         12606 => x"7d57810b",
         12607 => x"8318347d",
         12608 => x"51feed80",
         12609 => x"3f84b8e4",
         12610 => x"08567584",
         12611 => x"b8e40c9f",
         12612 => x"3d0d0476",
         12613 => x"902a5574",
         12614 => x"80ec1734",
         12615 => x"74882a57",
         12616 => x"7680ed17",
         12617 => x"34fefd39",
         12618 => x"7b902a5b",
         12619 => x"7a80cc17",
         12620 => x"347a882a",
         12621 => x"557480cd",
         12622 => x"17347d59",
         12623 => x"a00b80d8",
         12624 => x"1ab81b57",
         12625 => x"5856fea1",
         12626 => x"397b902a",
         12627 => x"58779418",
         12628 => x"3477882a",
         12629 => x"5c7b9518",
         12630 => x"34695590",
         12631 => x"0b8b1634",
         12632 => x"7d57810b",
         12633 => x"8318347d",
         12634 => x"51feec98",
         12635 => x"3f84b8e4",
         12636 => x"0856ff96",
         12637 => x"39d13d0d",
         12638 => x"b33db43d",
         12639 => x"0870595b",
         12640 => x"5f79802e",
         12641 => x"9b387970",
         12642 => x"81055b33",
         12643 => x"709f2656",
         12644 => x"5675ba2e",
         12645 => x"81b83874",
         12646 => x"ed3875ba",
         12647 => x"2e81af38",
         12648 => x"8253b13d",
         12649 => x"fefc0552",
         12650 => x"b23d51ff",
         12651 => x"abb43f84",
         12652 => x"b8e40856",
         12653 => x"84b8e408",
         12654 => x"802e8a38",
         12655 => x"7584b8e4",
         12656 => x"0cb13d0d",
         12657 => x"047fa63d",
         12658 => x"0cb23d08",
         12659 => x"52a53d70",
         12660 => x"5259ff9f",
         12661 => x"af3f84b8",
         12662 => x"e4085684",
         12663 => x"b8e408dc",
         12664 => x"380281bb",
         12665 => x"053381a0",
         12666 => x"065d8656",
         12667 => x"7cce38a0",
         12668 => x"0b923dae",
         12669 => x"3d085858",
         12670 => x"55757081",
         12671 => x"05573377",
         12672 => x"70810559",
         12673 => x"34ff1555",
         12674 => x"74ef3899",
         12675 => x"3d58b078",
         12676 => x"7a585855",
         12677 => x"75708105",
         12678 => x"57337770",
         12679 => x"81055934",
         12680 => x"ff155574",
         12681 => x"ef38b33d",
         12682 => x"08527751",
         12683 => x"ff9ed53f",
         12684 => x"84b8e408",
         12685 => x"5684b8e4",
         12686 => x"0885d838",
         12687 => x"6aa83d08",
         12688 => x"2e81cb38",
         12689 => x"880b84b8",
         12690 => x"e40cb13d",
         12691 => x"0d047633",
         12692 => x"d0117081",
         12693 => x"ff065757",
         12694 => x"58748926",
         12695 => x"91388217",
         12696 => x"7881ff06",
         12697 => x"d0055d59",
         12698 => x"787a2e80",
         12699 => x"fa38807f",
         12700 => x"0883e4d4",
         12701 => x"7008725d",
         12702 => x"5e5f5f5c",
         12703 => x"7a708105",
         12704 => x"5c337970",
         12705 => x"81055b33",
         12706 => x"ff9f125a",
         12707 => x"58567799",
         12708 => x"268938e0",
         12709 => x"167081ff",
         12710 => x"065755ff",
         12711 => x"9f175877",
         12712 => x"99268938",
         12713 => x"e0177081",
         12714 => x"ff065855",
         12715 => x"7530709f",
         12716 => x"2a595575",
         12717 => x"772e0981",
         12718 => x"06853877",
         12719 => x"ffbe3878",
         12720 => x"7a327030",
         12721 => x"7072079f",
         12722 => x"2a7a075d",
         12723 => x"58557a80",
         12724 => x"2e953881",
         12725 => x"1c841e5e",
         12726 => x"5c7b8324",
         12727 => x"fdc2387c",
         12728 => x"087e5a5b",
         12729 => x"ff96397b",
         12730 => x"8324fdb4",
         12731 => x"38797f0c",
         12732 => x"8253b13d",
         12733 => x"fefc0552",
         12734 => x"b23d51ff",
         12735 => x"a8e43f84",
         12736 => x"b8e40856",
         12737 => x"84b8e408",
         12738 => x"fdb238fd",
         12739 => x"b8396caa",
         12740 => x"3d082e09",
         12741 => x"8106feac",
         12742 => x"387751ff",
         12743 => x"8da83f84",
         12744 => x"b8e40856",
         12745 => x"84b8e408",
         12746 => x"fd92386f",
         12747 => x"58930b8d",
         12748 => x"19028805",
         12749 => x"80cd0558",
         12750 => x"565a7570",
         12751 => x"81055733",
         12752 => x"75708105",
         12753 => x"5734ff1a",
         12754 => x"5a79ef38",
         12755 => x"0280cb05",
         12756 => x"338b1934",
         12757 => x"8b183370",
         12758 => x"842a8106",
         12759 => x"40567e89",
         12760 => x"3875a007",
         12761 => x"57768b19",
         12762 => x"347f5d81",
         12763 => x"0b831e34",
         12764 => x"8b183370",
         12765 => x"842a8106",
         12766 => x"575c7580",
         12767 => x"2e81c538",
         12768 => x"a73d086b",
         12769 => x"2e81bd38",
         12770 => x"7f9b1933",
         12771 => x"9a1a3371",
         12772 => x"882b0772",
         12773 => x"3341585c",
         12774 => x"577d832e",
         12775 => x"82e038fe",
         12776 => x"169c1808",
         12777 => x"fe055e56",
         12778 => x"757d2782",
         12779 => x"c7388a17",
         12780 => x"22767129",
         12781 => x"b0190805",
         12782 => x"575e7580",
         12783 => x"2e82b538",
         12784 => x"757a5d58",
         12785 => x"b4170876",
         12786 => x"2eaa3883",
         12787 => x"17335f7e",
         12788 => x"83bc3881",
         12789 => x"547553b8",
         12790 => x"17528117",
         12791 => x"3351fee3",
         12792 => x"f13f84b8",
         12793 => x"e408802e",
         12794 => x"8538ff58",
         12795 => x"815c77b4",
         12796 => x"180c7f57",
         12797 => x"7b80d818",
         12798 => x"56567bfb",
         12799 => x"bf388115",
         12800 => x"335a79ae",
         12801 => x"2e098106",
         12802 => x"bb386a70",
         12803 => x"83ffff06",
         12804 => x"5d567b80",
         12805 => x"f218347b",
         12806 => x"882a5877",
         12807 => x"80f31834",
         12808 => x"76335b7a",
         12809 => x"832e0981",
         12810 => x"06933875",
         12811 => x"902a5e7d",
         12812 => x"80ec1834",
         12813 => x"7d882a56",
         12814 => x"7580ed18",
         12815 => x"347f5781",
         12816 => x"0b831834",
         12817 => x"7808aa3d",
         12818 => x"08b23d08",
         12819 => x"575c5674",
         12820 => x"ff2e9538",
         12821 => x"74527851",
         12822 => x"fefba23f",
         12823 => x"84b8e408",
         12824 => x"5584b8e4",
         12825 => x"0880f538",
         12826 => x"b8165c98",
         12827 => x"19085780",
         12828 => x"5ab41608",
         12829 => x"772eb438",
         12830 => x"8316337a",
         12831 => x"595f7e7a",
         12832 => x"2e098106",
         12833 => x"81a83881",
         12834 => x"547653b8",
         12835 => x"16528116",
         12836 => x"3351fee2",
         12837 => x"bd3f84b8",
         12838 => x"e408802e",
         12839 => x"8538ff57",
         12840 => x"815876b4",
         12841 => x"170c7755",
         12842 => x"77aa389c",
         12843 => x"19085ae5",
         12844 => x"7a34810b",
         12845 => x"83173490",
         12846 => x"19087b27",
         12847 => x"a5388052",
         12848 => x"7851fefc",
         12849 => x"ae3f84b8",
         12850 => x"e4085584",
         12851 => x"b8e40880",
         12852 => x"2eff9838",
         12853 => x"82567484",
         12854 => x"2ef9e138",
         12855 => x"745674f9",
         12856 => x"db387f51",
         12857 => x"fee59d3f",
         12858 => x"84b8e408",
         12859 => x"84b8e40c",
         12860 => x"b13d0d04",
         12861 => x"820b84b8",
         12862 => x"e40cb13d",
         12863 => x"0d049518",
         12864 => x"33941933",
         12865 => x"71982b71",
         12866 => x"902b0778",
         12867 => x"0758565c",
         12868 => x"fd8d3984",
         12869 => x"b8e40884",
         12870 => x"2efbfe38",
         12871 => x"84b8e408",
         12872 => x"802efea0",
         12873 => x"387584b8",
         12874 => x"e40cb13d",
         12875 => x"0d048154",
         12876 => x"b4160853",
         12877 => x"7b528116",
         12878 => x"3351fee2",
         12879 => x"943f8158",
         12880 => x"84b8e408",
         12881 => x"7a2e0981",
         12882 => x"06fedb38",
         12883 => x"84b8e408",
         12884 => x"831734b4",
         12885 => x"1608a817",
         12886 => x"083184b8",
         12887 => x"e4085955",
         12888 => x"74a01708",
         12889 => x"27fea038",
         12890 => x"8216335d",
         12891 => x"7c822e09",
         12892 => x"8106fe93",
         12893 => x"388154b4",
         12894 => x"1608a017",
         12895 => x"0805537b",
         12896 => x"52811633",
         12897 => x"51fee1c9",
         12898 => x"3f7958fd",
         12899 => x"fa398154",
         12900 => x"b4170853",
         12901 => x"b8177053",
         12902 => x"81183352",
         12903 => x"5bfee1b1",
         12904 => x"3f815c84",
         12905 => x"b8e408fc",
         12906 => x"c93884b8",
         12907 => x"e4088318",
         12908 => x"34b41708",
         12909 => x"a8180831",
         12910 => x"84b8e408",
         12911 => x"5d5574a0",
         12912 => x"180827fc",
         12913 => x"8e388217",
         12914 => x"335d7c82",
         12915 => x"2e098106",
         12916 => x"fc813881",
         12917 => x"54b41708",
         12918 => x"a0180805",
         12919 => x"537a5281",
         12920 => x"173351fe",
         12921 => x"e0eb3f79",
         12922 => x"5cfbe839",
         12923 => x"ec3d0d02",
         12924 => x"80df0533",
         12925 => x"02840580",
         12926 => x"e3053356",
         12927 => x"57825396",
         12928 => x"3dcc0552",
         12929 => x"973d51ff",
         12930 => x"a2d83f84",
         12931 => x"b8e40856",
         12932 => x"84b8e408",
         12933 => x"802e8a38",
         12934 => x"7584b8e4",
         12935 => x"0c963d0d",
         12936 => x"04785a66",
         12937 => x"52963dd0",
         12938 => x"0551ff96",
         12939 => x"d73f84b8",
         12940 => x"e4085684",
         12941 => x"b8e408e0",
         12942 => x"380280cf",
         12943 => x"053381a0",
         12944 => x"06548656",
         12945 => x"73d23874",
         12946 => x"a7066171",
         12947 => x"098b1233",
         12948 => x"71067a74",
         12949 => x"06075156",
         12950 => x"5755738b",
         12951 => x"17347855",
         12952 => x"810b8316",
         12953 => x"347851fe",
         12954 => x"e29a3f84",
         12955 => x"b8e40884",
         12956 => x"b8e40c96",
         12957 => x"3d0d04ec",
         12958 => x"3d0d6757",
         12959 => x"8253963d",
         12960 => x"cc055297",
         12961 => x"3d51ffa1",
         12962 => x"d93f84b8",
         12963 => x"e4085584",
         12964 => x"b8e40880",
         12965 => x"2e8a3874",
         12966 => x"84b8e40c",
         12967 => x"963d0d04",
         12968 => x"785a6652",
         12969 => x"963dd005",
         12970 => x"51ff95d8",
         12971 => x"3f84b8e4",
         12972 => x"085584b8",
         12973 => x"e408e038",
         12974 => x"0280cf05",
         12975 => x"3381a006",
         12976 => x"56865575",
         12977 => x"d2386084",
         12978 => x"18228619",
         12979 => x"2271902b",
         12980 => x"07595956",
         12981 => x"76961734",
         12982 => x"76882a55",
         12983 => x"74971734",
         12984 => x"76902a58",
         12985 => x"77981734",
         12986 => x"76982a54",
         12987 => x"73991734",
         12988 => x"7857810b",
         12989 => x"83183478",
         12990 => x"51fee188",
         12991 => x"3f84b8e4",
         12992 => x"0884b8e4",
         12993 => x"0c963d0d",
         12994 => x"04e83d0d",
         12995 => x"6b6d5d5b",
         12996 => x"80539a3d",
         12997 => x"cc05529b",
         12998 => x"3d51ffa0",
         12999 => x"c53f84b8",
         13000 => x"e40884b8",
         13001 => x"e4083070",
         13002 => x"84b8e408",
         13003 => x"07802551",
         13004 => x"56577a80",
         13005 => x"2e8b3881",
         13006 => x"7076065a",
         13007 => x"567881a4",
         13008 => x"38763070",
         13009 => x"78078025",
         13010 => x"565b7b80",
         13011 => x"2e818c38",
         13012 => x"81707606",
         13013 => x"5a587880",
         13014 => x"2e818038",
         13015 => x"7ca41108",
         13016 => x"5856805a",
         13017 => x"b4160877",
         13018 => x"2e82f638",
         13019 => x"8316337a",
         13020 => x"5a55747a",
         13021 => x"2e098106",
         13022 => x"81983881",
         13023 => x"547653b8",
         13024 => x"16528116",
         13025 => x"3351fedc",
         13026 => x"c93f84b8",
         13027 => x"e408802e",
         13028 => x"8538ff57",
         13029 => x"815976b4",
         13030 => x"170c7857",
         13031 => x"78bd387c",
         13032 => x"70335658",
         13033 => x"80c35674",
         13034 => x"832e8b38",
         13035 => x"80e45674",
         13036 => x"842e8338",
         13037 => x"a7567518",
         13038 => x"b8058311",
         13039 => x"33821233",
         13040 => x"71902b71",
         13041 => x"882b0781",
         13042 => x"14337072",
         13043 => x"07882b75",
         13044 => x"33710762",
         13045 => x"0c5f5d5e",
         13046 => x"57595676",
         13047 => x"84b8e40c",
         13048 => x"9a3d0d04",
         13049 => x"7c5e8040",
         13050 => x"80528e3d",
         13051 => x"705255fe",
         13052 => x"f48b3f84",
         13053 => x"b8e40857",
         13054 => x"84b8e408",
         13055 => x"802e818d",
         13056 => x"3876842e",
         13057 => x"098106fe",
         13058 => x"b838807b",
         13059 => x"348057fe",
         13060 => x"b0397754",
         13061 => x"b4160853",
         13062 => x"b8167053",
         13063 => x"81173352",
         13064 => x"5bfedcad",
         13065 => x"3f775984",
         13066 => x"b8e4087a",
         13067 => x"2e098106",
         13068 => x"fee83884",
         13069 => x"b8e40883",
         13070 => x"1734b416",
         13071 => x"08a81708",
         13072 => x"3184b8e4",
         13073 => x"085a5574",
         13074 => x"a0170827",
         13075 => x"fead3882",
         13076 => x"16335574",
         13077 => x"822e0981",
         13078 => x"06fea038",
         13079 => x"7754b416",
         13080 => x"08a01708",
         13081 => x"05537a52",
         13082 => x"81163351",
         13083 => x"fedbe23f",
         13084 => x"79598154",
         13085 => x"7653b816",
         13086 => x"52811633",
         13087 => x"51fedad2",
         13088 => x"3f84b8e4",
         13089 => x"08802efe",
         13090 => x"8d38fe86",
         13091 => x"39755274",
         13092 => x"51fef8bb",
         13093 => x"3f84b8e4",
         13094 => x"085784b8",
         13095 => x"e408fee1",
         13096 => x"3884b8e4",
         13097 => x"0884b8e4",
         13098 => x"08665c59",
         13099 => x"59791881",
         13100 => x"197c1b57",
         13101 => x"59567533",
         13102 => x"75348119",
         13103 => x"598a7827",
         13104 => x"ec388b70",
         13105 => x"1c575880",
         13106 => x"76347780",
         13107 => x"2efcf238",
         13108 => x"ff187b11",
         13109 => x"70335c57",
         13110 => x"5879a02e",
         13111 => x"ea38fce1",
         13112 => x"397957fd",
         13113 => x"ba39e13d",
         13114 => x"0d8253a1",
         13115 => x"3dffb405",
         13116 => x"52a23d51",
         13117 => x"ff9ceb3f",
         13118 => x"84b8e408",
         13119 => x"5684b8e4",
         13120 => x"0882a638",
         13121 => x"8f3d5d8b",
         13122 => x"7d5755a0",
         13123 => x"76708105",
         13124 => x"5834ff15",
         13125 => x"5574f438",
         13126 => x"74a33d08",
         13127 => x"70337081",
         13128 => x"ff065b58",
         13129 => x"585a9f78",
         13130 => x"2781b738",
         13131 => x"a23d903d",
         13132 => x"5c5c7581",
         13133 => x"ff068118",
         13134 => x"57557481",
         13135 => x"f538757c",
         13136 => x"0c7483ff",
         13137 => x"ff2681ff",
         13138 => x"387451a1",
         13139 => x"953f83b5",
         13140 => x"5284b8e4",
         13141 => x"08519fdc",
         13142 => x"3f84b8e4",
         13143 => x"0883ffff",
         13144 => x"06577680",
         13145 => x"2e81e038",
         13146 => x"83e5f40b",
         13147 => x"83e5f433",
         13148 => x"7081ff06",
         13149 => x"5b565878",
         13150 => x"802e81d6",
         13151 => x"38745678",
         13152 => x"772e9938",
         13153 => x"81187033",
         13154 => x"7081ff06",
         13155 => x"57575874",
         13156 => x"802e8938",
         13157 => x"74772e09",
         13158 => x"8106e938",
         13159 => x"7581ff06",
         13160 => x"597881a3",
         13161 => x"3881ff77",
         13162 => x"2781f838",
         13163 => x"79892681",
         13164 => x"963881ff",
         13165 => x"77278f38",
         13166 => x"76882a55",
         13167 => x"747b7081",
         13168 => x"055d3481",
         13169 => x"1a5a767b",
         13170 => x"7081055d",
         13171 => x"34811aa3",
         13172 => x"3d087033",
         13173 => x"7081ff06",
         13174 => x"5b58585a",
         13175 => x"779f26fe",
         13176 => x"d1388f3d",
         13177 => x"33578656",
         13178 => x"7681e52e",
         13179 => x"bc387980",
         13180 => x"2e993802",
         13181 => x"b7055679",
         13182 => x"1670335c",
         13183 => x"5c7aa02e",
         13184 => x"09810687",
         13185 => x"38ff1a5a",
         13186 => x"79ed387d",
         13187 => x"45804780",
         13188 => x"52953d70",
         13189 => x"5256feef",
         13190 => x"e43f84b8",
         13191 => x"e4085584",
         13192 => x"b8e40880",
         13193 => x"2eb43874",
         13194 => x"567584b8",
         13195 => x"e40ca13d",
         13196 => x"0d0483b5",
         13197 => x"5274519e",
         13198 => x"e73f84b8",
         13199 => x"e40883ff",
         13200 => x"ff065574",
         13201 => x"fdf83886",
         13202 => x"567584b8",
         13203 => x"e40ca13d",
         13204 => x"0d0483e5",
         13205 => x"f43356fe",
         13206 => x"c3398152",
         13207 => x"7551fef4",
         13208 => x"ee3f84b8",
         13209 => x"e4085584",
         13210 => x"b8e40880",
         13211 => x"c1387980",
         13212 => x"2e82c438",
         13213 => x"8b6c7e59",
         13214 => x"57557670",
         13215 => x"81055833",
         13216 => x"76708105",
         13217 => x"5834ff15",
         13218 => x"5574ef38",
         13219 => x"7d5d810b",
         13220 => x"831e347d",
         13221 => x"51fed9ec",
         13222 => x"3f84b8e4",
         13223 => x"08557456",
         13224 => x"ff87398a",
         13225 => x"7a27fe8a",
         13226 => x"388656ff",
         13227 => x"9c3984b8",
         13228 => x"e408842e",
         13229 => x"098106fe",
         13230 => x"ee388055",
         13231 => x"79752efe",
         13232 => x"e6387508",
         13233 => x"75537652",
         13234 => x"58feeeb1",
         13235 => x"3f84b8e4",
         13236 => x"085784b8",
         13237 => x"e408752e",
         13238 => x"09810681",
         13239 => x"843884b8",
         13240 => x"e408b819",
         13241 => x"5c5a9816",
         13242 => x"08578059",
         13243 => x"b4180877",
         13244 => x"2eb23883",
         13245 => x"18335574",
         13246 => x"792e0981",
         13247 => x"0681d738",
         13248 => x"81547653",
         13249 => x"b8185281",
         13250 => x"183351fe",
         13251 => x"d5c43f84",
         13252 => x"b8e40880",
         13253 => x"2e8538ff",
         13254 => x"57815976",
         13255 => x"b4190c78",
         13256 => x"5778be38",
         13257 => x"789c1708",
         13258 => x"7033575a",
         13259 => x"577481e5",
         13260 => x"2e819e38",
         13261 => x"74307080",
         13262 => x"25780756",
         13263 => x"5c74802e",
         13264 => x"81d73881",
         13265 => x"1a5a7981",
         13266 => x"2ea53881",
         13267 => x"527551fe",
         13268 => x"efa13f84",
         13269 => x"b8e40857",
         13270 => x"84b8e408",
         13271 => x"802eff86",
         13272 => x"38875576",
         13273 => x"842efdbf",
         13274 => x"38765576",
         13275 => x"fdb938a0",
         13276 => x"6c575580",
         13277 => x"76708105",
         13278 => x"5834ff15",
         13279 => x"5574f438",
         13280 => x"6b56880b",
         13281 => x"8b17348b",
         13282 => x"6c7e5957",
         13283 => x"55767081",
         13284 => x"05583376",
         13285 => x"70810558",
         13286 => x"34ff1555",
         13287 => x"74802efd",
         13288 => x"eb387670",
         13289 => x"81055833",
         13290 => x"76708105",
         13291 => x"5834ff15",
         13292 => x"5574da38",
         13293 => x"fdd6396b",
         13294 => x"5ae57a34",
         13295 => x"7d5d810b",
         13296 => x"831e347d",
         13297 => x"51fed7bc",
         13298 => x"3f84b8e4",
         13299 => x"0855fdce",
         13300 => x"398157fe",
         13301 => x"df398154",
         13302 => x"b4180853",
         13303 => x"7a528118",
         13304 => x"3351fed4",
         13305 => x"ec3f84b8",
         13306 => x"e408792e",
         13307 => x"09810680",
         13308 => x"c33884b8",
         13309 => x"e4088319",
         13310 => x"34b41808",
         13311 => x"a8190831",
         13312 => x"5c7ba019",
         13313 => x"08278a38",
         13314 => x"82183355",
         13315 => x"74822eb1",
         13316 => x"3884b8e4",
         13317 => x"0859fde8",
         13318 => x"39745a81",
         13319 => x"527551fe",
         13320 => x"edd13f84",
         13321 => x"b8e40857",
         13322 => x"84b8e408",
         13323 => x"802efdb6",
         13324 => x"38feae39",
         13325 => x"81705859",
         13326 => x"78802efd",
         13327 => x"e738fea1",
         13328 => x"398154b4",
         13329 => x"1808a019",
         13330 => x"0805537a",
         13331 => x"52811833",
         13332 => x"51fed3fd",
         13333 => x"3ffda939",
         13334 => x"f23d0d60",
         13335 => x"62028805",
         13336 => x"80cb0533",
         13337 => x"5e5b5789",
         13338 => x"5676802e",
         13339 => x"9f387608",
         13340 => x"5574802e",
         13341 => x"97387433",
         13342 => x"5473802e",
         13343 => x"8f388615",
         13344 => x"22841822",
         13345 => x"59597878",
         13346 => x"2e81c238",
         13347 => x"8054735f",
         13348 => x"7581a538",
         13349 => x"91173356",
         13350 => x"75819d38",
         13351 => x"79802e81",
         13352 => x"a2388c17",
         13353 => x"08819c38",
         13354 => x"90173370",
         13355 => x"812a8106",
         13356 => x"565d7480",
         13357 => x"2e818c38",
         13358 => x"7e8a1122",
         13359 => x"70892b70",
         13360 => x"557c5457",
         13361 => x"5c59fd87",
         13362 => x"dc3fff15",
         13363 => x"7a067030",
         13364 => x"7072079f",
         13365 => x"2a84b8e4",
         13366 => x"0805901c",
         13367 => x"08794253",
         13368 => x"5f555881",
         13369 => x"78278838",
         13370 => x"9c190878",
         13371 => x"26833882",
         13372 => x"58777856",
         13373 => x"5b805974",
         13374 => x"527651fe",
         13375 => x"d8873f81",
         13376 => x"157f5555",
         13377 => x"9c140875",
         13378 => x"26833882",
         13379 => x"5584b8e4",
         13380 => x"08812e81",
         13381 => x"dc3884b8",
         13382 => x"e408ff2e",
         13383 => x"81d83884",
         13384 => x"b8e40881",
         13385 => x"c5388119",
         13386 => x"59787d2e",
         13387 => x"bb387478",
         13388 => x"2e098106",
         13389 => x"c2388756",
         13390 => x"75547384",
         13391 => x"b8e40c90",
         13392 => x"3d0d0487",
         13393 => x"0b84b8e4",
         13394 => x"0c903d0d",
         13395 => x"04811533",
         13396 => x"51fed0ac",
         13397 => x"3f84b8e4",
         13398 => x"08810654",
         13399 => x"73fead38",
         13400 => x"73770855",
         13401 => x"56fea739",
         13402 => x"7b802e81",
         13403 => x"8e387a7d",
         13404 => x"56587c80",
         13405 => x"2eab3881",
         13406 => x"18547481",
         13407 => x"2e80e638",
         13408 => x"73537752",
         13409 => x"7e51fedd",
         13410 => x"dd3f84b8",
         13411 => x"e4085684",
         13412 => x"b8e408ff",
         13413 => x"a3387781",
         13414 => x"19ff1757",
         13415 => x"595e74d7",
         13416 => x"387e7e90",
         13417 => x"120c557b",
         13418 => x"802eff8c",
         13419 => x"387a8818",
         13420 => x"0c798c18",
         13421 => x"0c901733",
         13422 => x"80c0075c",
         13423 => x"7b901834",
         13424 => x"9c1508fe",
         13425 => x"05941608",
         13426 => x"585a767a",
         13427 => x"26fee938",
         13428 => x"767d3194",
         13429 => x"160c8415",
         13430 => x"3381075d",
         13431 => x"7c841634",
         13432 => x"7554fed6",
         13433 => x"39ff54ff",
         13434 => x"9739745b",
         13435 => x"8059febe",
         13436 => x"398254fe",
         13437 => x"c5398154",
         13438 => x"fec039ff",
         13439 => x"1b5effa1",
         13440 => x"3984b8f0",
         13441 => x"08e33d0d",
         13442 => x"a33d08a5",
         13443 => x"3d080288",
         13444 => x"05818705",
         13445 => x"3344425f",
         13446 => x"ff0ba23d",
         13447 => x"08705f5b",
         13448 => x"4079802e",
         13449 => x"858a3879",
         13450 => x"7081055b",
         13451 => x"33709f26",
         13452 => x"565675ba",
         13453 => x"2e859b38",
         13454 => x"74ed3875",
         13455 => x"ba2e8592",
         13456 => x"3884d0c0",
         13457 => x"33568076",
         13458 => x"2484e538",
         13459 => x"75101084",
         13460 => x"d0ac0570",
         13461 => x"08565a74",
         13462 => x"802e8438",
         13463 => x"80753475",
         13464 => x"1684b8d8",
         13465 => x"113384b8",
         13466 => x"d9123340",
         13467 => x"5b5d8152",
         13468 => x"7951fece",
         13469 => x"a93f84b8",
         13470 => x"e40881ff",
         13471 => x"06708106",
         13472 => x"5d568357",
         13473 => x"7b84ab38",
         13474 => x"75822a81",
         13475 => x"06408a57",
         13476 => x"7f849f38",
         13477 => x"9f3dfc05",
         13478 => x"53835279",
         13479 => x"51fed0b0",
         13480 => x"3f84b8e4",
         13481 => x"08849838",
         13482 => x"6d557480",
         13483 => x"2e849038",
         13484 => x"74828080",
         13485 => x"26848838",
         13486 => x"ff157506",
         13487 => x"557483ff",
         13488 => x"387e802e",
         13489 => x"88388480",
         13490 => x"7f2683f8",
         13491 => x"387e8180",
         13492 => x"0a2683f0",
         13493 => x"38ff1f7f",
         13494 => x"06557483",
         13495 => x"e7387e89",
         13496 => x"2aa63d08",
         13497 => x"892a7089",
         13498 => x"2b77594c",
         13499 => x"475b6080",
         13500 => x"2e85ab38",
         13501 => x"65307080",
         13502 => x"25770756",
         13503 => x"5f915774",
         13504 => x"83b0387d",
         13505 => x"802e84df",
         13506 => x"38815474",
         13507 => x"53605279",
         13508 => x"51fecdbe",
         13509 => x"3f815784",
         13510 => x"b8e40883",
         13511 => x"95386083",
         13512 => x"ff053361",
         13513 => x"83fe0533",
         13514 => x"71882b07",
         13515 => x"59568e57",
         13516 => x"7782d4d5",
         13517 => x"2e098106",
         13518 => x"82f8387d",
         13519 => x"90296105",
         13520 => x"83b21133",
         13521 => x"44586280",
         13522 => x"2e82e738",
         13523 => x"83b61883",
         13524 => x"11338212",
         13525 => x"3371902b",
         13526 => x"71882b07",
         13527 => x"81143370",
         13528 => x"7207882b",
         13529 => x"75337107",
         13530 => x"83ba1f83",
         13531 => x"11338212",
         13532 => x"3371902b",
         13533 => x"71882b07",
         13534 => x"81143370",
         13535 => x"7207882b",
         13536 => x"75337107",
         13537 => x"5ca23d0c",
         13538 => x"42a33d0c",
         13539 => x"a33d0c44",
         13540 => x"4e544559",
         13541 => x"4f415a4b",
         13542 => x"784d8e57",
         13543 => x"80ff7927",
         13544 => x"82903893",
         13545 => x"577a8180",
         13546 => x"26828738",
         13547 => x"61812a70",
         13548 => x"81064549",
         13549 => x"63802e83",
         13550 => x"f9386187",
         13551 => x"06456482",
         13552 => x"2e893861",
         13553 => x"81064766",
         13554 => x"83f43883",
         13555 => x"6e70304a",
         13556 => x"46437a58",
         13557 => x"62832e8a",
         13558 => x"c2387aae",
         13559 => x"38788c2a",
         13560 => x"57810b83",
         13561 => x"e6882256",
         13562 => x"5874802e",
         13563 => x"9d387477",
         13564 => x"26983883",
         13565 => x"e6885677",
         13566 => x"10821770",
         13567 => x"22575758",
         13568 => x"74802e86",
         13569 => x"38767527",
         13570 => x"ee387752",
         13571 => x"7851fd81",
         13572 => x"943f84b8",
         13573 => x"e4081084",
         13574 => x"055584b8",
         13575 => x"e4089ff5",
         13576 => x"26963881",
         13577 => x"0b84b8e4",
         13578 => x"081084b8",
         13579 => x"e4080571",
         13580 => x"11722a83",
         13581 => x"05574c43",
         13582 => x"83ff1589",
         13583 => x"2a5d815c",
         13584 => x"a0477b1f",
         13585 => x"7d116805",
         13586 => x"6611ff05",
         13587 => x"706b0672",
         13588 => x"31584e57",
         13589 => x"4462832e",
         13590 => x"89b83874",
         13591 => x"1d5d7790",
         13592 => x"29167060",
         13593 => x"31565774",
         13594 => x"792682f2",
         13595 => x"38787c31",
         13596 => x"7d317853",
         13597 => x"70683152",
         13598 => x"56fd80a9",
         13599 => x"3f84b8e4",
         13600 => x"08406283",
         13601 => x"2e89f638",
         13602 => x"62822e09",
         13603 => x"810682dd",
         13604 => x"3883fff5",
         13605 => x"0b84b8e4",
         13606 => x"082782ac",
         13607 => x"387a89f9",
         13608 => x"38771855",
         13609 => x"7480c026",
         13610 => x"89ef3874",
         13611 => x"5bfea339",
         13612 => x"8b577684",
         13613 => x"b8e40c9f",
         13614 => x"3d0d84b8",
         13615 => x"f00c0481",
         13616 => x"4efbfe39",
         13617 => x"930b84b8",
         13618 => x"e40c9f3d",
         13619 => x"0d84b8f0",
         13620 => x"0c047c33",
         13621 => x"d0117081",
         13622 => x"ff065757",
         13623 => x"57748926",
         13624 => x"9138821d",
         13625 => x"7781ff06",
         13626 => x"d0055d58",
         13627 => x"777a2e81",
         13628 => x"b238800b",
         13629 => x"83e4d45f",
         13630 => x"5c7d087d",
         13631 => x"575b7a70",
         13632 => x"81055c33",
         13633 => x"76708105",
         13634 => x"5833ff9f",
         13635 => x"12455957",
         13636 => x"62992689",
         13637 => x"38e01770",
         13638 => x"81ff0658",
         13639 => x"44ff9f18",
         13640 => x"45649926",
         13641 => x"8938e018",
         13642 => x"7081ff06",
         13643 => x"59467630",
         13644 => x"709f2a5a",
         13645 => x"4776782e",
         13646 => x"09810685",
         13647 => x"3878ffbe",
         13648 => x"38757a32",
         13649 => x"70307072",
         13650 => x"079f2a7b",
         13651 => x"075d4a4a",
         13652 => x"7a802e80",
         13653 => x"ce38811c",
         13654 => x"841f5f5c",
         13655 => x"837c25ff",
         13656 => x"98387f56",
         13657 => x"f9e0399f",
         13658 => x"3df80553",
         13659 => x"81527951",
         13660 => x"fecadd3f",
         13661 => x"815784b8",
         13662 => x"e408feb6",
         13663 => x"3861832a",
         13664 => x"770684b8",
         13665 => x"e4084056",
         13666 => x"758338bf",
         13667 => x"5f6c558e",
         13668 => x"577e7526",
         13669 => x"fe9c3874",
         13670 => x"7f3159fb",
         13671 => x"fb398156",
         13672 => x"fad2397b",
         13673 => x"8324ffba",
         13674 => x"387b7aa3",
         13675 => x"3d0c56f9",
         13676 => x"95396181",
         13677 => x"06489357",
         13678 => x"67802efd",
         13679 => x"f538826e",
         13680 => x"70304a46",
         13681 => x"43fc8b39",
         13682 => x"84b8e408",
         13683 => x"9ff5269d",
         13684 => x"387a8b38",
         13685 => x"77185b81",
         13686 => x"807b27fb",
         13687 => x"f5388e57",
         13688 => x"7684b8e4",
         13689 => x"0c9f3d0d",
         13690 => x"84b8f00c",
         13691 => x"04805562",
         13692 => x"812e8699",
         13693 => x"389ff560",
         13694 => x"278b3874",
         13695 => x"81065b8e",
         13696 => x"577afdae",
         13697 => x"38848061",
         13698 => x"57558076",
         13699 => x"70810558",
         13700 => x"34ff1555",
         13701 => x"74f4388b",
         13702 => x"6183e4a0",
         13703 => x"59575576",
         13704 => x"70810558",
         13705 => x"33767081",
         13706 => x"055834ff",
         13707 => x"155574ef",
         13708 => x"38608b05",
         13709 => x"45746534",
         13710 => x"82618c05",
         13711 => x"3477618d",
         13712 => x"05347b83",
         13713 => x"ffff064b",
         13714 => x"6a618e05",
         13715 => x"346a882a",
         13716 => x"5c7b618f",
         13717 => x"05348161",
         13718 => x"90053462",
         13719 => x"83327030",
         13720 => x"5a488061",
         13721 => x"91053478",
         13722 => x"9e2a8206",
         13723 => x"49686192",
         13724 => x"05346c56",
         13725 => x"7583ffff",
         13726 => x"2686ad38",
         13727 => x"7583ffff",
         13728 => x"06557461",
         13729 => x"93053474",
         13730 => x"882a4c6b",
         13731 => x"61940534",
         13732 => x"f8619505",
         13733 => x"34bf6198",
         13734 => x"05348061",
         13735 => x"990534ff",
         13736 => x"619a0534",
         13737 => x"80619b05",
         13738 => x"347e619c",
         13739 => x"05347e88",
         13740 => x"2a486761",
         13741 => x"9d05347e",
         13742 => x"902a4c6b",
         13743 => x"619e0534",
         13744 => x"7e982a84",
         13745 => x"b8f00c84",
         13746 => x"b8f00861",
         13747 => x"9f053462",
         13748 => x"832e85f7",
         13749 => x"388061a7",
         13750 => x"05348061",
         13751 => x"a80534a1",
         13752 => x"61a90534",
         13753 => x"80cc61aa",
         13754 => x"05347c83",
         13755 => x"ffff0655",
         13756 => x"74619605",
         13757 => x"3474882a",
         13758 => x"4b6a6197",
         13759 => x"0534ff80",
         13760 => x"61a40534",
         13761 => x"a961a605",
         13762 => x"349361ab",
         13763 => x"0583e4ac",
         13764 => x"59575576",
         13765 => x"70810558",
         13766 => x"33767081",
         13767 => x"055834ff",
         13768 => x"155574ef",
         13769 => x"386083fe",
         13770 => x"054980d5",
         13771 => x"69346083",
         13772 => x"ff054bff",
         13773 => x"aa6b3481",
         13774 => x"547e5360",
         13775 => x"527951fe",
         13776 => x"c68f3f81",
         13777 => x"5784b8e4",
         13778 => x"08fae738",
         13779 => x"60175c62",
         13780 => x"832e879c",
         13781 => x"38696157",
         13782 => x"55807670",
         13783 => x"81055834",
         13784 => x"ff155574",
         13785 => x"f4386375",
         13786 => x"415b6283",
         13787 => x"2e86c038",
         13788 => x"87fffff8",
         13789 => x"5762812e",
         13790 => x"8338f857",
         13791 => x"76613476",
         13792 => x"882a7c45",
         13793 => x"55746470",
         13794 => x"81054634",
         13795 => x"76902a59",
         13796 => x"78647081",
         13797 => x"05463476",
         13798 => x"982a5675",
         13799 => x"64347c57",
         13800 => x"65597666",
         13801 => x"26833876",
         13802 => x"5978547a",
         13803 => x"53605279",
         13804 => x"51fec59d",
         13805 => x"3f84b8e4",
         13806 => x"0885e638",
         13807 => x"84806157",
         13808 => x"55807670",
         13809 => x"81055834",
         13810 => x"ff155574",
         13811 => x"f438781b",
         13812 => x"777a3158",
         13813 => x"5b76c938",
         13814 => x"7f810540",
         13815 => x"7f802eff",
         13816 => x"89387756",
         13817 => x"62832e83",
         13818 => x"38665665",
         13819 => x"55756626",
         13820 => x"83387555",
         13821 => x"74547a53",
         13822 => x"60527951",
         13823 => x"fec4d23f",
         13824 => x"84b8e408",
         13825 => x"859b3874",
         13826 => x"1b767631",
         13827 => x"575b75db",
         13828 => x"388c5862",
         13829 => x"832e9338",
         13830 => x"86586c83",
         13831 => x"ffff268a",
         13832 => x"38845862",
         13833 => x"822e8338",
         13834 => x"81587d84",
         13835 => x"c1386183",
         13836 => x"2a81065e",
         13837 => x"7d81b338",
         13838 => x"84806156",
         13839 => x"59807570",
         13840 => x"81055734",
         13841 => x"ff195978",
         13842 => x"f43880d5",
         13843 => x"6934ffaa",
         13844 => x"6b346083",
         13845 => x"be054778",
         13846 => x"67348167",
         13847 => x"81053481",
         13848 => x"67820534",
         13849 => x"78678305",
         13850 => x"34776784",
         13851 => x"05346c43",
         13852 => x"80fdc152",
         13853 => x"621f51fc",
         13854 => x"f8ab3ffe",
         13855 => x"67850534",
         13856 => x"84b8e408",
         13857 => x"822abf07",
         13858 => x"57766786",
         13859 => x"053484b8",
         13860 => x"e4086787",
         13861 => x"05347e61",
         13862 => x"83c60534",
         13863 => x"676183c7",
         13864 => x"05346b61",
         13865 => x"83c80534",
         13866 => x"84b8f008",
         13867 => x"6183c905",
         13868 => x"34626183",
         13869 => x"ca053462",
         13870 => x"882a4564",
         13871 => x"6183cb05",
         13872 => x"3462902a",
         13873 => x"58776183",
         13874 => x"cc053462",
         13875 => x"982a5f7e",
         13876 => x"6183cd05",
         13877 => x"34815478",
         13878 => x"53605279",
         13879 => x"51fec2f1",
         13880 => x"3f815784",
         13881 => x"b8e408f7",
         13882 => x"c9388053",
         13883 => x"80527951",
         13884 => x"fec3dd3f",
         13885 => x"815784b8",
         13886 => x"e408f7b6",
         13887 => x"3884b8e4",
         13888 => x"0884b8e4",
         13889 => x"0c9f3d0d",
         13890 => x"84b8f00c",
         13891 => x"046255f9",
         13892 => x"e439741c",
         13893 => x"6416455c",
         13894 => x"f6c4397a",
         13895 => x"ae387891",
         13896 => x"2a57810b",
         13897 => x"83e69822",
         13898 => x"56587480",
         13899 => x"2e9d3874",
         13900 => x"77269838",
         13901 => x"83e69856",
         13902 => x"77108217",
         13903 => x"70225757",
         13904 => x"5874802e",
         13905 => x"86387675",
         13906 => x"27ee3877",
         13907 => x"527851fc",
         13908 => x"f6d33f84",
         13909 => x"b8e40810",
         13910 => x"10848705",
         13911 => x"70892a5e",
         13912 => x"5ca05c80",
         13913 => x"0b84b8e4",
         13914 => x"08fc808a",
         13915 => x"055847fd",
         13916 => x"fff00a77",
         13917 => x"27f5cb38",
         13918 => x"8e57f8e4",
         13919 => x"3984b8e4",
         13920 => x"0883fff5",
         13921 => x"26f8e638",
         13922 => x"7af8d338",
         13923 => x"77812a5b",
         13924 => x"7af4bf38",
         13925 => x"8e57f8c8",
         13926 => x"39688106",
         13927 => x"4463802e",
         13928 => x"f8af3883",
         13929 => x"43f4ab39",
         13930 => x"7561a005",
         13931 => x"3475882a",
         13932 => x"496861a1",
         13933 => x"05347590",
         13934 => x"2a5b7a61",
         13935 => x"a2053475",
         13936 => x"982a5776",
         13937 => x"61a30534",
         13938 => x"f9c63980",
         13939 => x"6180c305",
         13940 => x"34806180",
         13941 => x"c40534a1",
         13942 => x"6180c505",
         13943 => x"3480cc61",
         13944 => x"80c60534",
         13945 => x"7c61a405",
         13946 => x"347c882a",
         13947 => x"5c7b61a5",
         13948 => x"05347c90",
         13949 => x"2a597861",
         13950 => x"a605347c",
         13951 => x"982a5675",
         13952 => x"61a70534",
         13953 => x"8261ac05",
         13954 => x"348061ad",
         13955 => x"05348061",
         13956 => x"ae053480",
         13957 => x"61af0534",
         13958 => x"8161b005",
         13959 => x"348061b1",
         13960 => x"05348661",
         13961 => x"b2053480",
         13962 => x"61b30534",
         13963 => x"ff806180",
         13964 => x"c00534a9",
         13965 => x"6180c205",
         13966 => x"34936180",
         13967 => x"c70583e4",
         13968 => x"c0595755",
         13969 => x"76708105",
         13970 => x"58337670",
         13971 => x"81055834",
         13972 => x"ff155574",
         13973 => x"802ef9cd",
         13974 => x"38767081",
         13975 => x"05583376",
         13976 => x"70810558",
         13977 => x"34ff1555",
         13978 => x"74da38f9",
         13979 => x"b8398154",
         13980 => x"80536052",
         13981 => x"7951febe",
         13982 => x"d93f8157",
         13983 => x"84b8e408",
         13984 => x"f4b0387d",
         13985 => x"90296105",
         13986 => x"42776283",
         13987 => x"b2053476",
         13988 => x"5484b8e4",
         13989 => x"08536052",
         13990 => x"7951febf",
         13991 => x"b43ffcc3",
         13992 => x"39810b84",
         13993 => x"b8e40c9f",
         13994 => x"3d0d84b8",
         13995 => x"f00c04f8",
         13996 => x"61347b4a",
         13997 => x"ff6a7081",
         13998 => x"054c34ff",
         13999 => x"6a708105",
         14000 => x"4c34ff6a",
         14001 => x"34ff6184",
         14002 => x"0534ff61",
         14003 => x"850534ff",
         14004 => x"61860534",
         14005 => x"ff618705",
         14006 => x"34ff6188",
         14007 => x"0534ff61",
         14008 => x"890534ff",
         14009 => x"618a0534",
         14010 => x"8f65347c",
         14011 => x"57f9b139",
         14012 => x"7654861f",
         14013 => x"53605279",
         14014 => x"51febed5",
         14015 => x"3f848061",
         14016 => x"56578075",
         14017 => x"70810557",
         14018 => x"34ff1757",
         14019 => x"76f43860",
         14020 => x"5c80d27c",
         14021 => x"7081055e",
         14022 => x"347b5580",
         14023 => x"d2757081",
         14024 => x"05573480",
         14025 => x"e1757081",
         14026 => x"05573480",
         14027 => x"c1753480",
         14028 => x"f26183e4",
         14029 => x"053480f2",
         14030 => x"6183e505",
         14031 => x"3480c161",
         14032 => x"83e60534",
         14033 => x"80e16183",
         14034 => x"e705347f",
         14035 => x"ff055b7a",
         14036 => x"6183e805",
         14037 => x"347a882a",
         14038 => x"59786183",
         14039 => x"e905347a",
         14040 => x"902a5675",
         14041 => x"6183ea05",
         14042 => x"347a982a",
         14043 => x"407f6183",
         14044 => x"eb053482",
         14045 => x"6183ec05",
         14046 => x"34766183",
         14047 => x"ed053476",
         14048 => x"6183ee05",
         14049 => x"34766183",
         14050 => x"ef053480",
         14051 => x"d56934ff",
         14052 => x"aa6b3481",
         14053 => x"54871f53",
         14054 => x"60527951",
         14055 => x"febdb23f",
         14056 => x"8154811f",
         14057 => x"53605279",
         14058 => x"51febda5",
         14059 => x"3f696157",
         14060 => x"55f7a639",
         14061 => x"f43d0d7e",
         14062 => x"615b5b80",
         14063 => x"7b61ff05",
         14064 => x"5a575776",
         14065 => x"7825b838",
         14066 => x"8d3d598e",
         14067 => x"3df80554",
         14068 => x"81537852",
         14069 => x"7951ff9a",
         14070 => x"b43f7b81",
         14071 => x"2e098106",
         14072 => x"9e388d3d",
         14073 => x"3355748d",
         14074 => x"2e903874",
         14075 => x"76708105",
         14076 => x"58348117",
         14077 => x"57748a2e",
         14078 => x"86387777",
         14079 => x"24cd3880",
         14080 => x"76347a55",
         14081 => x"76833876",
         14082 => x"557484b8",
         14083 => x"e40c8e3d",
         14084 => x"0d04f73d",
         14085 => x"0d7b0284",
         14086 => x"05b30533",
         14087 => x"5957778a",
         14088 => x"2e80d538",
         14089 => x"84170856",
         14090 => x"8076249e",
         14091 => x"38881708",
         14092 => x"77178c05",
         14093 => x"56597775",
         14094 => x"34811655",
         14095 => x"74bb248e",
         14096 => x"38748418",
         14097 => x"0c811988",
         14098 => x"180c8b3d",
         14099 => x"0d048b3d",
         14100 => x"fc055474",
         14101 => x"538c1752",
         14102 => x"760851ff",
         14103 => x"9ed13f74",
         14104 => x"7a327030",
         14105 => x"7072079f",
         14106 => x"2a703084",
         14107 => x"1b0c811c",
         14108 => x"881b0c5a",
         14109 => x"5656d339",
         14110 => x"8d527651",
         14111 => x"ff943fff",
         14112 => x"a339e33d",
         14113 => x"0d0280ff",
         14114 => x"05338d3d",
         14115 => x"585880cc",
         14116 => x"77575580",
         14117 => x"76708105",
         14118 => x"5834ff15",
         14119 => x"5574f438",
         14120 => x"a13d0877",
         14121 => x"0c778a2e",
         14122 => x"80f7387c",
         14123 => x"56807624",
         14124 => x"80c0387d",
         14125 => x"77178c05",
         14126 => x"56597775",
         14127 => x"34811655",
         14128 => x"74bb24b8",
         14129 => x"38748418",
         14130 => x"0c811988",
         14131 => x"180c7c55",
         14132 => x"8075249e",
         14133 => x"389f3dff",
         14134 => x"ac115575",
         14135 => x"54c00552",
         14136 => x"760851ff",
         14137 => x"9dc93f84",
         14138 => x"b8e40886",
         14139 => x"387c7a2e",
         14140 => x"ba38ff0b",
         14141 => x"84b8e40c",
         14142 => x"9f3d0d04",
         14143 => x"9f3dffb0",
         14144 => x"11557554",
         14145 => x"c0055276",
         14146 => x"0851ff9d",
         14147 => x"a23f747b",
         14148 => x"32703070",
         14149 => x"72079f2a",
         14150 => x"7030525a",
         14151 => x"5656ffa5",
         14152 => x"398d5276",
         14153 => x"51fdeb3f",
         14154 => x"ff81397d",
         14155 => x"84b8e40c",
         14156 => x"9f3d0d04",
         14157 => x"fd3d0d75",
         14158 => x"0284059a",
         14159 => x"05225253",
         14160 => x"80527280",
         14161 => x"ff269038",
         14162 => x"7283ffff",
         14163 => x"06527184",
         14164 => x"b8e40c85",
         14165 => x"3d0d0483",
         14166 => x"ffff7327",
         14167 => x"547083b5",
         14168 => x"2e098106",
         14169 => x"e9387380",
         14170 => x"2ee43883",
         14171 => x"e6a82251",
         14172 => x"72712e9c",
         14173 => x"38811270",
         14174 => x"83ffff06",
         14175 => x"53547180",
         14176 => x"ff268d38",
         14177 => x"711083e6",
         14178 => x"a8057022",
         14179 => x"5151e139",
         14180 => x"81801270",
         14181 => x"81ff0684",
         14182 => x"b8e40c53",
         14183 => x"853d0d04",
         14184 => x"fe3d0d02",
         14185 => x"92052202",
         14186 => x"84059605",
         14187 => x"22535180",
         14188 => x"537080ff",
         14189 => x"268c3870",
         14190 => x"537284b8",
         14191 => x"e40c843d",
         14192 => x"0d047183",
         14193 => x"b52e0981",
         14194 => x"06ef3870",
         14195 => x"81ff26e9",
         14196 => x"38701083",
         14197 => x"e4a80570",
         14198 => x"2284b8e4",
         14199 => x"0c51843d",
         14200 => x"0d04fb3d",
         14201 => x"0d775170",
         14202 => x"83ffff26",
         14203 => x"80e13870",
         14204 => x"83ffff06",
         14205 => x"83e8a856",
         14206 => x"56759fff",
         14207 => x"2680d938",
         14208 => x"74708205",
         14209 => x"56227571",
         14210 => x"30708025",
         14211 => x"737a2607",
         14212 => x"54565353",
         14213 => x"70b73871",
         14214 => x"70820553",
         14215 => x"22727188",
         14216 => x"2a545681",
         14217 => x"ff067014",
         14218 => x"52547076",
         14219 => x"24b13871",
         14220 => x"cf387310",
         14221 => x"15707082",
         14222 => x"05522254",
         14223 => x"73307080",
         14224 => x"25757926",
         14225 => x"07535552",
         14226 => x"70802ecb",
         14227 => x"38755170",
         14228 => x"84b8e40c",
         14229 => x"873d0d04",
         14230 => x"83ec9c55",
         14231 => x"ffa23971",
         14232 => x"8826ea38",
         14233 => x"71101083",
         14234 => x"c9d00554",
         14235 => x"730804c7",
         14236 => x"a0167083",
         14237 => x"ffff0657",
         14238 => x"517551d3",
         14239 => x"39ffb016",
         14240 => x"7083ffff",
         14241 => x"065751f1",
         14242 => x"39881670",
         14243 => x"83ffff06",
         14244 => x"5751e639",
         14245 => x"e6167083",
         14246 => x"ffff0657",
         14247 => x"51db39d0",
         14248 => x"167083ff",
         14249 => x"ff065751",
         14250 => x"d039e016",
         14251 => x"7083ffff",
         14252 => x"065751c5",
         14253 => x"39f01670",
         14254 => x"83ffff06",
         14255 => x"5751ffb9",
         14256 => x"39757331",
         14257 => x"81067671",
         14258 => x"317083ff",
         14259 => x"ff065852",
         14260 => x"55ffa639",
         14261 => x"75733110",
         14262 => x"75057022",
         14263 => x"5252feef",
         14264 => x"39000000",
         14265 => x"00ffffff",
         14266 => x"ff00ffff",
         14267 => x"ffff00ff",
         14268 => x"ffffff00",
         14269 => x"0000198b",
         14270 => x"00001980",
         14271 => x"00001975",
         14272 => x"0000196a",
         14273 => x"0000195f",
         14274 => x"00001954",
         14275 => x"00001949",
         14276 => x"0000193e",
         14277 => x"00001933",
         14278 => x"00001928",
         14279 => x"0000191d",
         14280 => x"00001912",
         14281 => x"00001907",
         14282 => x"000018fc",
         14283 => x"000018f1",
         14284 => x"000018e6",
         14285 => x"000018db",
         14286 => x"000018d0",
         14287 => x"000018c5",
         14288 => x"000018ba",
         14289 => x"00001ebf",
         14290 => x"00001f59",
         14291 => x"00001f59",
         14292 => x"00001f59",
         14293 => x"00001f59",
         14294 => x"00001f59",
         14295 => x"00001f59",
         14296 => x"00001f59",
         14297 => x"00001f59",
         14298 => x"00001f59",
         14299 => x"00001f59",
         14300 => x"00001f59",
         14301 => x"00001f59",
         14302 => x"00001f59",
         14303 => x"00001f59",
         14304 => x"00001f59",
         14305 => x"00001f59",
         14306 => x"00001f59",
         14307 => x"00001f59",
         14308 => x"00001f59",
         14309 => x"00001f59",
         14310 => x"00001f59",
         14311 => x"00001f59",
         14312 => x"00001f59",
         14313 => x"00001f59",
         14314 => x"00001f59",
         14315 => x"00001f59",
         14316 => x"00001f59",
         14317 => x"00001f59",
         14318 => x"00001f59",
         14319 => x"00001f59",
         14320 => x"00001f59",
         14321 => x"00001f59",
         14322 => x"00001f59",
         14323 => x"00001f59",
         14324 => x"00001f59",
         14325 => x"00001f59",
         14326 => x"00001f59",
         14327 => x"00001f59",
         14328 => x"00001f59",
         14329 => x"00001f59",
         14330 => x"00001f59",
         14331 => x"00001f59",
         14332 => x"00002471",
         14333 => x"00001f59",
         14334 => x"00001f59",
         14335 => x"00001f59",
         14336 => x"00001f59",
         14337 => x"00001f59",
         14338 => x"00001f59",
         14339 => x"00001f59",
         14340 => x"00001f59",
         14341 => x"00001f59",
         14342 => x"00001f59",
         14343 => x"00001f59",
         14344 => x"00001f59",
         14345 => x"00001f59",
         14346 => x"00001f59",
         14347 => x"00001f59",
         14348 => x"00001f59",
         14349 => x"00002407",
         14350 => x"00002306",
         14351 => x"00001f59",
         14352 => x"0000228a",
         14353 => x"000024a8",
         14354 => x"00002367",
         14355 => x"0000222c",
         14356 => x"000021ce",
         14357 => x"00001f59",
         14358 => x"00001f59",
         14359 => x"00001f59",
         14360 => x"00001f59",
         14361 => x"00001f59",
         14362 => x"00001f59",
         14363 => x"00001f59",
         14364 => x"00001f59",
         14365 => x"00001f59",
         14366 => x"00001f59",
         14367 => x"00001f59",
         14368 => x"00001f59",
         14369 => x"00001f59",
         14370 => x"00001f59",
         14371 => x"00001f59",
         14372 => x"00001f59",
         14373 => x"00001f59",
         14374 => x"00001f59",
         14375 => x"00001f59",
         14376 => x"00001f59",
         14377 => x"00001f59",
         14378 => x"00001f59",
         14379 => x"00001f59",
         14380 => x"00001f59",
         14381 => x"00001f59",
         14382 => x"00001f59",
         14383 => x"00001f59",
         14384 => x"00001f59",
         14385 => x"00001f59",
         14386 => x"00001f59",
         14387 => x"00001f59",
         14388 => x"00001f59",
         14389 => x"00001f59",
         14390 => x"00001f59",
         14391 => x"00001f59",
         14392 => x"00001f59",
         14393 => x"00001f59",
         14394 => x"00001f59",
         14395 => x"00001f59",
         14396 => x"00001f59",
         14397 => x"00001f59",
         14398 => x"00001f59",
         14399 => x"00001f59",
         14400 => x"00001f59",
         14401 => x"00001f59",
         14402 => x"00001f59",
         14403 => x"00001f59",
         14404 => x"00001f59",
         14405 => x"00001f59",
         14406 => x"00001f59",
         14407 => x"00001f59",
         14408 => x"00001f59",
         14409 => x"000021ab",
         14410 => x"00002170",
         14411 => x"00001f59",
         14412 => x"00001f59",
         14413 => x"00001f59",
         14414 => x"00001f59",
         14415 => x"00001f59",
         14416 => x"00001f59",
         14417 => x"00001f59",
         14418 => x"00001f59",
         14419 => x"00002163",
         14420 => x"00002158",
         14421 => x"00001f59",
         14422 => x"00002141",
         14423 => x"00001f59",
         14424 => x"00002151",
         14425 => x"00002147",
         14426 => x"0000213a",
         14427 => x"00003212",
         14428 => x"0000322a",
         14429 => x"00003236",
         14430 => x"00003242",
         14431 => x"0000324e",
         14432 => x"0000321e",
         14433 => x"00003b86",
         14434 => x"00003a74",
         14435 => x"000038f0",
         14436 => x"0000363e",
         14437 => x"00003a10",
         14438 => x"000034cd",
         14439 => x"0000378a",
         14440 => x"00003663",
         14441 => x"000039ba",
         14442 => x"00003692",
         14443 => x"00003701",
         14444 => x"00003919",
         14445 => x"000034cd",
         14446 => x"000038f0",
         14447 => x"000037fa",
         14448 => x"0000378a",
         14449 => x"000034cd",
         14450 => x"000034cd",
         14451 => x"00003701",
         14452 => x"00003692",
         14453 => x"00003663",
         14454 => x"0000363e",
         14455 => x"0000466b",
         14456 => x"00004684",
         14457 => x"000046a9",
         14458 => x"000046ca",
         14459 => x"0000462b",
         14460 => x"000046ef",
         14461 => x"00004644",
         14462 => x"00004794",
         14463 => x"00004751",
         14464 => x"00004751",
         14465 => x"00004751",
         14466 => x"00004751",
         14467 => x"00004751",
         14468 => x"00004751",
         14469 => x"0000472a",
         14470 => x"00004751",
         14471 => x"00004751",
         14472 => x"00004751",
         14473 => x"00004751",
         14474 => x"00004751",
         14475 => x"00004751",
         14476 => x"00004751",
         14477 => x"00004751",
         14478 => x"00004751",
         14479 => x"00004751",
         14480 => x"00004751",
         14481 => x"00004751",
         14482 => x"00004751",
         14483 => x"00004751",
         14484 => x"00004751",
         14485 => x"00004751",
         14486 => x"00004751",
         14487 => x"00004751",
         14488 => x"00004751",
         14489 => x"00004751",
         14490 => x"00004751",
         14491 => x"00004751",
         14492 => x"00004869",
         14493 => x"00004857",
         14494 => x"00004844",
         14495 => x"00004831",
         14496 => x"0000475b",
         14497 => x"0000481f",
         14498 => x"0000480c",
         14499 => x"00004774",
         14500 => x"00004751",
         14501 => x"00004774",
         14502 => x"000047fc",
         14503 => x"00004879",
         14504 => x"000047a5",
         14505 => x"00004783",
         14506 => x"000047ea",
         14507 => x"000047d8",
         14508 => x"000047c6",
         14509 => x"000047b7",
         14510 => x"00004751",
         14511 => x"0000475b",
         14512 => x"000053f7",
         14513 => x"00005566",
         14514 => x"00005538",
         14515 => x"0000548f",
         14516 => x"0000546c",
         14517 => x"0000544b",
         14518 => x"00005421",
         14519 => x"000055f1",
         14520 => x"00005278",
         14521 => x"000055cb",
         14522 => x"000057ba",
         14523 => x"00005278",
         14524 => x"00005278",
         14525 => x"00005278",
         14526 => x"00005278",
         14527 => x"00005278",
         14528 => x"00005278",
         14529 => x"00005594",
         14530 => x"000057a2",
         14531 => x"00005659",
         14532 => x"00005278",
         14533 => x"00005278",
         14534 => x"00005278",
         14535 => x"00005278",
         14536 => x"00005278",
         14537 => x"00005278",
         14538 => x"00005278",
         14539 => x"00005278",
         14540 => x"00005278",
         14541 => x"00005278",
         14542 => x"00005278",
         14543 => x"00005278",
         14544 => x"00005278",
         14545 => x"00005278",
         14546 => x"00005278",
         14547 => x"00005278",
         14548 => x"00005278",
         14549 => x"00005278",
         14550 => x"00005278",
         14551 => x"00005516",
         14552 => x"00005278",
         14553 => x"00005278",
         14554 => x"00005278",
         14555 => x"000054b9",
         14556 => x"000053c8",
         14557 => x"0000536a",
         14558 => x"00005278",
         14559 => x"00005278",
         14560 => x"00005278",
         14561 => x"00005278",
         14562 => x"0000534f",
         14563 => x"00005278",
         14564 => x"00005332",
         14565 => x"0000599b",
         14566 => x"00005910",
         14567 => x"00005910",
         14568 => x"00005910",
         14569 => x"00005910",
         14570 => x"00005910",
         14571 => x"00005910",
         14572 => x"000058eb",
         14573 => x"00005910",
         14574 => x"00005910",
         14575 => x"00005910",
         14576 => x"00005910",
         14577 => x"00005910",
         14578 => x"00005910",
         14579 => x"00005910",
         14580 => x"00005910",
         14581 => x"00005910",
         14582 => x"00005910",
         14583 => x"00005910",
         14584 => x"00005910",
         14585 => x"00005910",
         14586 => x"00005910",
         14587 => x"00005910",
         14588 => x"00005910",
         14589 => x"00005910",
         14590 => x"00005910",
         14591 => x"00005910",
         14592 => x"00005910",
         14593 => x"00005910",
         14594 => x"00005910",
         14595 => x"000059ad",
         14596 => x"000059f5",
         14597 => x"000059e2",
         14598 => x"000059cf",
         14599 => x"000059bd",
         14600 => x"00005a80",
         14601 => x"00005a6d",
         14602 => x"00005a5d",
         14603 => x"00005910",
         14604 => x"00005a4d",
         14605 => x"00005a3d",
         14606 => x"00005a2b",
         14607 => x"00005a19",
         14608 => x"00005a07",
         14609 => x"00005978",
         14610 => x"00005967",
         14611 => x"00005956",
         14612 => x"0000593f",
         14613 => x"00005910",
         14614 => x"00005989",
         14615 => x"0000636a",
         14616 => x"000061c6",
         14617 => x"000061c6",
         14618 => x"000061c6",
         14619 => x"000061c6",
         14620 => x"000061c6",
         14621 => x"000061c6",
         14622 => x"000061c6",
         14623 => x"000061c6",
         14624 => x"000061c6",
         14625 => x"000061c6",
         14626 => x"000061c6",
         14627 => x"000061c6",
         14628 => x"000061c6",
         14629 => x"00005ee8",
         14630 => x"000061c6",
         14631 => x"000061c6",
         14632 => x"000061c6",
         14633 => x"000061c6",
         14634 => x"000061c6",
         14635 => x"000061c6",
         14636 => x"000063b4",
         14637 => x"000061c6",
         14638 => x"000061c6",
         14639 => x"0000633f",
         14640 => x"000061c6",
         14641 => x"00006356",
         14642 => x"00005ec7",
         14643 => x"00006328",
         14644 => x"0000ded4",
         14645 => x"0000dec1",
         14646 => x"0000deb5",
         14647 => x"0000deaa",
         14648 => x"0000de9f",
         14649 => x"0000de94",
         14650 => x"0000de89",
         14651 => x"0000de7d",
         14652 => x"0000de6f",
         14653 => x"00000e01",
         14654 => x"00000bfd",
         14655 => x"00000bfd",
         14656 => x"00000f49",
         14657 => x"00000bfd",
         14658 => x"00000bfd",
         14659 => x"00000bfd",
         14660 => x"00000bfd",
         14661 => x"00000bfd",
         14662 => x"00000bfd",
         14663 => x"00000bfd",
         14664 => x"00000dfd",
         14665 => x"00000bfd",
         14666 => x"00000f7f",
         14667 => x"00000f0d",
         14668 => x"00000bfd",
         14669 => x"00000bfd",
         14670 => x"00000bfd",
         14671 => x"00000bfd",
         14672 => x"00000bfd",
         14673 => x"00000bfd",
         14674 => x"00000bfd",
         14675 => x"00000bfd",
         14676 => x"00000bfd",
         14677 => x"00000bfd",
         14678 => x"00000bfd",
         14679 => x"00000bfd",
         14680 => x"00000bfd",
         14681 => x"00000bfd",
         14682 => x"00000bfd",
         14683 => x"00000bfd",
         14684 => x"00000bfd",
         14685 => x"00000bfd",
         14686 => x"00000bfd",
         14687 => x"00000bfd",
         14688 => x"00000bfd",
         14689 => x"00000bfd",
         14690 => x"00000bfd",
         14691 => x"00000bfd",
         14692 => x"00000bfd",
         14693 => x"00000bfd",
         14694 => x"00000bfd",
         14695 => x"00000bfd",
         14696 => x"00000bfd",
         14697 => x"00000bfd",
         14698 => x"00000bfd",
         14699 => x"00000bfd",
         14700 => x"00000bfd",
         14701 => x"00000bfd",
         14702 => x"00000bfd",
         14703 => x"00000bfd",
         14704 => x"00000f1d",
         14705 => x"00000bfd",
         14706 => x"00000bfd",
         14707 => x"00000bfd",
         14708 => x"00000bfd",
         14709 => x"00000e17",
         14710 => x"00000bfd",
         14711 => x"00000bfd",
         14712 => x"00000bfd",
         14713 => x"00000bfd",
         14714 => x"00000bfd",
         14715 => x"00000bfd",
         14716 => x"00000bfd",
         14717 => x"00000bfd",
         14718 => x"00000bfd",
         14719 => x"00000bfd",
         14720 => x"00000e2b",
         14721 => x"00000ee1",
         14722 => x"00000eb8",
         14723 => x"00000eb8",
         14724 => x"00000eb8",
         14725 => x"00000bfd",
         14726 => x"00000ee1",
         14727 => x"00000bfd",
         14728 => x"00000bfd",
         14729 => x"00000eff",
         14730 => x"00000bfd",
         14731 => x"00000bfd",
         14732 => x"00000c16",
         14733 => x"00000e0f",
         14734 => x"00000bfd",
         14735 => x"00000bfd",
         14736 => x"00000f58",
         14737 => x"00000bfd",
         14738 => x"00000c18",
         14739 => x"00000bfd",
         14740 => x"00000bfd",
         14741 => x"00000e17",
         14742 => x"64696e69",
         14743 => x"74000000",
         14744 => x"64696f63",
         14745 => x"746c0000",
         14746 => x"66696e69",
         14747 => x"74000000",
         14748 => x"666c6f61",
         14749 => x"64000000",
         14750 => x"66657865",
         14751 => x"63000000",
         14752 => x"6d636c65",
         14753 => x"61720000",
         14754 => x"6d636f70",
         14755 => x"79000000",
         14756 => x"6d646966",
         14757 => x"66000000",
         14758 => x"6d64756d",
         14759 => x"70000000",
         14760 => x"6d656200",
         14761 => x"6d656800",
         14762 => x"6d657700",
         14763 => x"68696400",
         14764 => x"68696500",
         14765 => x"68666400",
         14766 => x"68666500",
         14767 => x"63616c6c",
         14768 => x"00000000",
         14769 => x"6a6d7000",
         14770 => x"72657374",
         14771 => x"61727400",
         14772 => x"72657365",
         14773 => x"74000000",
         14774 => x"696e666f",
         14775 => x"00000000",
         14776 => x"74657374",
         14777 => x"00000000",
         14778 => x"636c7300",
         14779 => x"7a383000",
         14780 => x"74626173",
         14781 => x"69630000",
         14782 => x"6d626173",
         14783 => x"69630000",
         14784 => x"6b696c6f",
         14785 => x"00000000",
         14786 => x"65640000",
         14787 => x"556e6b6e",
         14788 => x"6f776e20",
         14789 => x"6572726f",
         14790 => x"722e0000",
         14791 => x"50617261",
         14792 => x"6d657465",
         14793 => x"72732069",
         14794 => x"6e636f72",
         14795 => x"72656374",
         14796 => x"2e000000",
         14797 => x"546f6f20",
         14798 => x"6d616e79",
         14799 => x"206f7065",
         14800 => x"6e206669",
         14801 => x"6c65732e",
         14802 => x"00000000",
         14803 => x"496e7375",
         14804 => x"66666963",
         14805 => x"69656e74",
         14806 => x"206d656d",
         14807 => x"6f72792e",
         14808 => x"00000000",
         14809 => x"46696c65",
         14810 => x"20697320",
         14811 => x"6c6f636b",
         14812 => x"65642e00",
         14813 => x"54696d65",
         14814 => x"6f75742c",
         14815 => x"206f7065",
         14816 => x"72617469",
         14817 => x"6f6e2063",
         14818 => x"616e6365",
         14819 => x"6c6c6564",
         14820 => x"2e000000",
         14821 => x"466f726d",
         14822 => x"61742061",
         14823 => x"626f7274",
         14824 => x"65642e00",
         14825 => x"4e6f2063",
         14826 => x"6f6d7061",
         14827 => x"7469626c",
         14828 => x"65206669",
         14829 => x"6c657379",
         14830 => x"7374656d",
         14831 => x"20666f75",
         14832 => x"6e64206f",
         14833 => x"6e206469",
         14834 => x"736b2e00",
         14835 => x"4469736b",
         14836 => x"206e6f74",
         14837 => x"20656e61",
         14838 => x"626c6564",
         14839 => x"2e000000",
         14840 => x"44726976",
         14841 => x"65206e75",
         14842 => x"6d626572",
         14843 => x"20697320",
         14844 => x"696e7661",
         14845 => x"6c69642e",
         14846 => x"00000000",
         14847 => x"53442069",
         14848 => x"73207772",
         14849 => x"69746520",
         14850 => x"70726f74",
         14851 => x"65637465",
         14852 => x"642e0000",
         14853 => x"46696c65",
         14854 => x"2068616e",
         14855 => x"646c6520",
         14856 => x"696e7661",
         14857 => x"6c69642e",
         14858 => x"00000000",
         14859 => x"46696c65",
         14860 => x"20616c72",
         14861 => x"65616479",
         14862 => x"20657869",
         14863 => x"7374732e",
         14864 => x"00000000",
         14865 => x"41636365",
         14866 => x"73732064",
         14867 => x"656e6965",
         14868 => x"642e0000",
         14869 => x"496e7661",
         14870 => x"6c696420",
         14871 => x"66696c65",
         14872 => x"6e616d65",
         14873 => x"2e000000",
         14874 => x"4e6f2070",
         14875 => x"61746820",
         14876 => x"666f756e",
         14877 => x"642e0000",
         14878 => x"4e6f2066",
         14879 => x"696c6520",
         14880 => x"666f756e",
         14881 => x"642e0000",
         14882 => x"4469736b",
         14883 => x"206e6f74",
         14884 => x"20726561",
         14885 => x"64792e00",
         14886 => x"496e7465",
         14887 => x"726e616c",
         14888 => x"20657272",
         14889 => x"6f722e00",
         14890 => x"4469736b",
         14891 => x"20457272",
         14892 => x"6f720000",
         14893 => x"53756363",
         14894 => x"6573732e",
         14895 => x"00000000",
         14896 => x"0a256c75",
         14897 => x"20627974",
         14898 => x"65732025",
         14899 => x"73206174",
         14900 => x"20256c75",
         14901 => x"20627974",
         14902 => x"65732f73",
         14903 => x"65632e0a",
         14904 => x"00000000",
         14905 => x"72656164",
         14906 => x"00000000",
         14907 => x"2530386c",
         14908 => x"58000000",
         14909 => x"3a202000",
         14910 => x"25303258",
         14911 => x"00000000",
         14912 => x"207c0000",
         14913 => x"7c000000",
         14914 => x"20200000",
         14915 => x"25303458",
         14916 => x"00000000",
         14917 => x"20202020",
         14918 => x"20202020",
         14919 => x"00000000",
         14920 => x"7a4f5300",
         14921 => x"2a2a2025",
         14922 => x"73202800",
         14923 => x"30362f30",
         14924 => x"332f3230",
         14925 => x"32310000",
         14926 => x"76312e31",
         14927 => x"66000000",
         14928 => x"205a5055",
         14929 => x"2c207265",
         14930 => x"76202530",
         14931 => x"32782920",
         14932 => x"25732025",
         14933 => x"73202a2a",
         14934 => x"0a0a0000",
         14935 => x"5a505520",
         14936 => x"496e7465",
         14937 => x"72727570",
         14938 => x"74204861",
         14939 => x"6e646c65",
         14940 => x"72000000",
         14941 => x"55415254",
         14942 => x"31205458",
         14943 => x"20696e74",
         14944 => x"65727275",
         14945 => x"70740000",
         14946 => x"55415254",
         14947 => x"31205258",
         14948 => x"20696e74",
         14949 => x"65727275",
         14950 => x"70740000",
         14951 => x"55415254",
         14952 => x"30205458",
         14953 => x"20696e74",
         14954 => x"65727275",
         14955 => x"70740000",
         14956 => x"55415254",
         14957 => x"30205258",
         14958 => x"20696e74",
         14959 => x"65727275",
         14960 => x"70740000",
         14961 => x"494f4354",
         14962 => x"4c205752",
         14963 => x"20696e74",
         14964 => x"65727275",
         14965 => x"70740000",
         14966 => x"494f4354",
         14967 => x"4c205244",
         14968 => x"20696e74",
         14969 => x"65727275",
         14970 => x"70740000",
         14971 => x"50533220",
         14972 => x"696e7465",
         14973 => x"72727570",
         14974 => x"74000000",
         14975 => x"54696d65",
         14976 => x"7220696e",
         14977 => x"74657272",
         14978 => x"75707400",
         14979 => x"53657474",
         14980 => x"696e6720",
         14981 => x"75702074",
         14982 => x"696d6572",
         14983 => x"2e2e2e00",
         14984 => x"456e6162",
         14985 => x"6c696e67",
         14986 => x"2074696d",
         14987 => x"65722e2e",
         14988 => x"2e000000",
         14989 => x"6175746f",
         14990 => x"65786563",
         14991 => x"2e626174",
         14992 => x"00000000",
         14993 => x"7a4f535f",
         14994 => x"7a70752e",
         14995 => x"68737400",
         14996 => x"4661696c",
         14997 => x"65642074",
         14998 => x"6f20696e",
         14999 => x"69746961",
         15000 => x"6c697365",
         15001 => x"20736420",
         15002 => x"63617264",
         15003 => x"20302c20",
         15004 => x"706c6561",
         15005 => x"73652069",
         15006 => x"6e697420",
         15007 => x"6d616e75",
         15008 => x"616c6c79",
         15009 => x"2e000000",
         15010 => x"2a200000",
         15011 => x"25643a5c",
         15012 => x"25730000",
         15013 => x"303a0000",
         15014 => x"42616420",
         15015 => x"636f6d6d",
         15016 => x"616e642e",
         15017 => x"00000000",
         15018 => x"5a505500",
         15019 => x"62696e00",
         15020 => x"25643a5c",
         15021 => x"25735c25",
         15022 => x"732e2573",
         15023 => x"00000000",
         15024 => x"436f6c64",
         15025 => x"20726562",
         15026 => x"6f6f7469",
         15027 => x"6e672e2e",
         15028 => x"2e000000",
         15029 => x"52657374",
         15030 => x"61727469",
         15031 => x"6e672061",
         15032 => x"70706c69",
         15033 => x"63617469",
         15034 => x"6f6e2e2e",
         15035 => x"2e000000",
         15036 => x"43616c6c",
         15037 => x"696e6720",
         15038 => x"636f6465",
         15039 => x"20402025",
         15040 => x"30386c78",
         15041 => x"202e2e2e",
         15042 => x"0a000000",
         15043 => x"43616c6c",
         15044 => x"20726574",
         15045 => x"75726e65",
         15046 => x"6420636f",
         15047 => x"64652028",
         15048 => x"2564292e",
         15049 => x"0a000000",
         15050 => x"45786563",
         15051 => x"7574696e",
         15052 => x"6720636f",
         15053 => x"64652040",
         15054 => x"20253038",
         15055 => x"6c78202e",
         15056 => x"2e2e0a00",
         15057 => x"2530386c",
         15058 => x"58202530",
         15059 => x"386c582d",
         15060 => x"00000000",
         15061 => x"2530386c",
         15062 => x"58202530",
         15063 => x"34582d00",
         15064 => x"436f6d70",
         15065 => x"6172696e",
         15066 => x"672e2e2e",
         15067 => x"00000000",
         15068 => x"2530386c",
         15069 => x"78282530",
         15070 => x"3878292d",
         15071 => x"3e253038",
         15072 => x"6c782825",
         15073 => x"30387829",
         15074 => x"0a000000",
         15075 => x"436f7079",
         15076 => x"696e672e",
         15077 => x"2e2e0000",
         15078 => x"2530386c",
         15079 => x"58202530",
         15080 => x"32582d00",
         15081 => x"436c6561",
         15082 => x"72696e67",
         15083 => x"2e2e2e2e",
         15084 => x"00000000",
         15085 => x"44756d70",
         15086 => x"204d656d",
         15087 => x"6f727900",
         15088 => x"0a436f6d",
         15089 => x"706c6574",
         15090 => x"652e0000",
         15091 => x"25643a5c",
         15092 => x"25735c25",
         15093 => x"73000000",
         15094 => x"4d656d6f",
         15095 => x"72792065",
         15096 => x"78686175",
         15097 => x"73746564",
         15098 => x"2c206361",
         15099 => x"6e6e6f74",
         15100 => x"2070726f",
         15101 => x"63657373",
         15102 => x"20636f6d",
         15103 => x"6d616e64",
         15104 => x"2e000000",
         15105 => x"3f3f3f00",
         15106 => x"25642f25",
         15107 => x"642f2564",
         15108 => x"2025643a",
         15109 => x"25643a25",
         15110 => x"642e2564",
         15111 => x"25640a00",
         15112 => x"536f4320",
         15113 => x"436f6e66",
         15114 => x"69677572",
         15115 => x"6174696f",
         15116 => x"6e000000",
         15117 => x"3a0a4465",
         15118 => x"76696365",
         15119 => x"7320696d",
         15120 => x"706c656d",
         15121 => x"656e7465",
         15122 => x"643a0000",
         15123 => x"41646472",
         15124 => x"65737365",
         15125 => x"733a0000",
         15126 => x"20202020",
         15127 => x"43505520",
         15128 => x"52657365",
         15129 => x"74205665",
         15130 => x"63746f72",
         15131 => x"20416464",
         15132 => x"72657373",
         15133 => x"203d2025",
         15134 => x"3038580a",
         15135 => x"00000000",
         15136 => x"20202020",
         15137 => x"43505520",
         15138 => x"4d656d6f",
         15139 => x"72792053",
         15140 => x"74617274",
         15141 => x"20416464",
         15142 => x"72657373",
         15143 => x"203d2025",
         15144 => x"3038580a",
         15145 => x"00000000",
         15146 => x"20202020",
         15147 => x"53746163",
         15148 => x"6b205374",
         15149 => x"61727420",
         15150 => x"41646472",
         15151 => x"65737320",
         15152 => x"20202020",
         15153 => x"203d2025",
         15154 => x"3038580a",
         15155 => x"00000000",
         15156 => x"4d697363",
         15157 => x"3a000000",
         15158 => x"20202020",
         15159 => x"5a505520",
         15160 => x"49642020",
         15161 => x"20202020",
         15162 => x"20202020",
         15163 => x"20202020",
         15164 => x"20202020",
         15165 => x"203d2025",
         15166 => x"3034580a",
         15167 => x"00000000",
         15168 => x"20202020",
         15169 => x"53797374",
         15170 => x"656d2043",
         15171 => x"6c6f636b",
         15172 => x"20467265",
         15173 => x"71202020",
         15174 => x"20202020",
         15175 => x"203d2025",
         15176 => x"642e2530",
         15177 => x"34644d48",
         15178 => x"7a0a0000",
         15179 => x"20202020",
         15180 => x"57697368",
         15181 => x"626f6e65",
         15182 => x"20534452",
         15183 => x"414d2043",
         15184 => x"6c6f636b",
         15185 => x"20467265",
         15186 => x"713d2025",
         15187 => x"642e2530",
         15188 => x"34644d48",
         15189 => x"7a0a0000",
         15190 => x"20202020",
         15191 => x"53445241",
         15192 => x"4d20436c",
         15193 => x"6f636b20",
         15194 => x"46726571",
         15195 => x"20202020",
         15196 => x"20202020",
         15197 => x"203d2025",
         15198 => x"642e2530",
         15199 => x"34644d48",
         15200 => x"7a0a0000",
         15201 => x"20202020",
         15202 => x"53504900",
         15203 => x"20202020",
         15204 => x"50533200",
         15205 => x"20202020",
         15206 => x"494f4354",
         15207 => x"4c000000",
         15208 => x"20202020",
         15209 => x"57422049",
         15210 => x"32430000",
         15211 => x"20202020",
         15212 => x"57495348",
         15213 => x"424f4e45",
         15214 => x"20425553",
         15215 => x"00000000",
         15216 => x"20202020",
         15217 => x"494e5452",
         15218 => x"20435452",
         15219 => x"4c202843",
         15220 => x"68616e6e",
         15221 => x"656c733d",
         15222 => x"25303264",
         15223 => x"292e0a00",
         15224 => x"20202020",
         15225 => x"54494d45",
         15226 => x"52312020",
         15227 => x"20202854",
         15228 => x"696d6572",
         15229 => x"7320203d",
         15230 => x"25303264",
         15231 => x"292e0a00",
         15232 => x"20202020",
         15233 => x"53442043",
         15234 => x"41524420",
         15235 => x"20202844",
         15236 => x"65766963",
         15237 => x"6573203d",
         15238 => x"25303264",
         15239 => x"292e0a00",
         15240 => x"20202020",
         15241 => x"52414d20",
         15242 => x"20202020",
         15243 => x"20202825",
         15244 => x"3038583a",
         15245 => x"25303858",
         15246 => x"292e0a00",
         15247 => x"20202020",
         15248 => x"4252414d",
         15249 => x"20202020",
         15250 => x"20202825",
         15251 => x"3038583a",
         15252 => x"25303858",
         15253 => x"292e0a00",
         15254 => x"20202020",
         15255 => x"494e534e",
         15256 => x"20425241",
         15257 => x"4d202825",
         15258 => x"3038583a",
         15259 => x"25303858",
         15260 => x"292e0a00",
         15261 => x"20202020",
         15262 => x"53445241",
         15263 => x"4d202020",
         15264 => x"20202825",
         15265 => x"3038583a",
         15266 => x"25303858",
         15267 => x"292e0a00",
         15268 => x"20202020",
         15269 => x"57422053",
         15270 => x"4452414d",
         15271 => x"20202825",
         15272 => x"3038583a",
         15273 => x"25303858",
         15274 => x"292e0a00",
         15275 => x"20286672",
         15276 => x"6f6d2053",
         15277 => x"6f432063",
         15278 => x"6f6e6669",
         15279 => x"67290000",
         15280 => x"556e6b6e",
         15281 => x"6f776e00",
         15282 => x"45564f6d",
         15283 => x"00000000",
         15284 => x"536d616c",
         15285 => x"6c000000",
         15286 => x"4d656469",
         15287 => x"756d0000",
         15288 => x"466c6578",
         15289 => x"00000000",
         15290 => x"45564f00",
         15291 => x"0000f048",
         15292 => x"01000000",
         15293 => x"00000002",
         15294 => x"0000f044",
         15295 => x"01000000",
         15296 => x"00000003",
         15297 => x"0000f040",
         15298 => x"01000000",
         15299 => x"00000004",
         15300 => x"0000f03c",
         15301 => x"01000000",
         15302 => x"00000005",
         15303 => x"0000f038",
         15304 => x"01000000",
         15305 => x"00000006",
         15306 => x"0000f034",
         15307 => x"01000000",
         15308 => x"00000007",
         15309 => x"0000f030",
         15310 => x"01000000",
         15311 => x"00000001",
         15312 => x"0000f02c",
         15313 => x"01000000",
         15314 => x"00000008",
         15315 => x"0000f028",
         15316 => x"01000000",
         15317 => x"0000000b",
         15318 => x"0000f024",
         15319 => x"01000000",
         15320 => x"00000009",
         15321 => x"0000f020",
         15322 => x"01000000",
         15323 => x"0000000a",
         15324 => x"0000f01c",
         15325 => x"04000000",
         15326 => x"0000000d",
         15327 => x"0000f018",
         15328 => x"04000000",
         15329 => x"0000000c",
         15330 => x"0000f014",
         15331 => x"04000000",
         15332 => x"0000000e",
         15333 => x"0000f010",
         15334 => x"03000000",
         15335 => x"0000000f",
         15336 => x"0000f00c",
         15337 => x"04000000",
         15338 => x"0000000f",
         15339 => x"0000f008",
         15340 => x"04000000",
         15341 => x"00000010",
         15342 => x"0000f004",
         15343 => x"04000000",
         15344 => x"00000011",
         15345 => x"0000f000",
         15346 => x"03000000",
         15347 => x"00000012",
         15348 => x"0000effc",
         15349 => x"03000000",
         15350 => x"00000013",
         15351 => x"0000eff8",
         15352 => x"03000000",
         15353 => x"00000014",
         15354 => x"0000eff4",
         15355 => x"03000000",
         15356 => x"00000015",
         15357 => x"1b5b4400",
         15358 => x"1b5b4300",
         15359 => x"1b5b4200",
         15360 => x"1b5b4100",
         15361 => x"1b5b367e",
         15362 => x"1b5b357e",
         15363 => x"1b5b347e",
         15364 => x"1b304600",
         15365 => x"1b5b337e",
         15366 => x"1b5b327e",
         15367 => x"1b5b317e",
         15368 => x"10000000",
         15369 => x"0e000000",
         15370 => x"0d000000",
         15371 => x"0b000000",
         15372 => x"08000000",
         15373 => x"06000000",
         15374 => x"05000000",
         15375 => x"04000000",
         15376 => x"03000000",
         15377 => x"02000000",
         15378 => x"01000000",
         15379 => x"43616e6e",
         15380 => x"6f74206f",
         15381 => x"70656e2f",
         15382 => x"63726561",
         15383 => x"74652068",
         15384 => x"6973746f",
         15385 => x"72792066",
         15386 => x"696c652c",
         15387 => x"20646973",
         15388 => x"61626c69",
         15389 => x"6e672e00",
         15390 => x"68697374",
         15391 => x"6f727900",
         15392 => x"68697374",
         15393 => x"00000000",
         15394 => x"21000000",
         15395 => x"2530366c",
         15396 => x"75202025",
         15397 => x"730a0000",
         15398 => x"4661696c",
         15399 => x"65642074",
         15400 => x"6f207265",
         15401 => x"73657420",
         15402 => x"74686520",
         15403 => x"68697374",
         15404 => x"6f727920",
         15405 => x"66696c65",
         15406 => x"20746f20",
         15407 => x"454f462e",
         15408 => x"00000000",
         15409 => x"3e25730a",
         15410 => x"00000000",
         15411 => x"1b5b317e",
         15412 => x"00000000",
         15413 => x"1b5b4100",
         15414 => x"1b5b4200",
         15415 => x"1b5b4300",
         15416 => x"1b5b4400",
         15417 => x"1b5b3130",
         15418 => x"7e000000",
         15419 => x"1b5b3131",
         15420 => x"7e000000",
         15421 => x"1b5b3132",
         15422 => x"7e000000",
         15423 => x"1b5b3133",
         15424 => x"7e000000",
         15425 => x"1b5b3134",
         15426 => x"7e000000",
         15427 => x"1b5b3135",
         15428 => x"7e000000",
         15429 => x"1b5b3137",
         15430 => x"7e000000",
         15431 => x"1b5b3138",
         15432 => x"7e000000",
         15433 => x"1b5b3139",
         15434 => x"7e000000",
         15435 => x"1b5b3230",
         15436 => x"7e000000",
         15437 => x"1b5b327e",
         15438 => x"00000000",
         15439 => x"1b5b337e",
         15440 => x"00000000",
         15441 => x"1b5b4600",
         15442 => x"1b5b357e",
         15443 => x"00000000",
         15444 => x"1b5b367e",
         15445 => x"00000000",
         15446 => x"583a2564",
         15447 => x"2c25642c",
         15448 => x"25642c25",
         15449 => x"642c2564",
         15450 => x"2c25643a",
         15451 => x"25303278",
         15452 => x"00000000",
         15453 => x"443a2564",
         15454 => x"2d25642d",
         15455 => x"25643a25",
         15456 => x"633a2564",
         15457 => x"2c25642c",
         15458 => x"25643a00",
         15459 => x"25642c00",
         15460 => x"4b3a2564",
         15461 => x"3a000000",
         15462 => x"25303278",
         15463 => x"2c000000",
         15464 => x"25635b25",
         15465 => x"643b2564",
         15466 => x"52000000",
         15467 => x"5265706f",
         15468 => x"72742043",
         15469 => x"7572736f",
         15470 => x"723a0000",
         15471 => x"55703a25",
         15472 => x"30327820",
         15473 => x"25303278",
         15474 => x"00000000",
         15475 => x"44773a25",
         15476 => x"30327820",
         15477 => x"25303278",
         15478 => x"00000000",
         15479 => x"48643a25",
         15480 => x"30327820",
         15481 => x"00000000",
         15482 => x"4e6f2074",
         15483 => x"65737420",
         15484 => x"64656669",
         15485 => x"6e65642e",
         15486 => x"00000000",
         15487 => x"53440000",
         15488 => x"222a3a3c",
         15489 => x"3e3f7c7f",
         15490 => x"00000000",
         15491 => x"2b2c3b3d",
         15492 => x"5b5d0000",
         15493 => x"46415400",
         15494 => x"46415433",
         15495 => x"32000000",
         15496 => x"ebfe904d",
         15497 => x"53444f53",
         15498 => x"352e3000",
         15499 => x"4e4f204e",
         15500 => x"414d4520",
         15501 => x"20202046",
         15502 => x"41542020",
         15503 => x"20202000",
         15504 => x"4e4f204e",
         15505 => x"414d4520",
         15506 => x"20202046",
         15507 => x"41543332",
         15508 => x"20202000",
         15509 => x"0000f1fc",
         15510 => x"00000000",
         15511 => x"00000000",
         15512 => x"00000000",
         15513 => x"01030507",
         15514 => x"090e1012",
         15515 => x"1416181c",
         15516 => x"1e000000",
         15517 => x"809a4541",
         15518 => x"8e418f80",
         15519 => x"45454549",
         15520 => x"49498e8f",
         15521 => x"9092924f",
         15522 => x"994f5555",
         15523 => x"59999a9b",
         15524 => x"9c9d9e9f",
         15525 => x"41494f55",
         15526 => x"a5a5a6a7",
         15527 => x"a8a9aaab",
         15528 => x"acadaeaf",
         15529 => x"b0b1b2b3",
         15530 => x"b4b5b6b7",
         15531 => x"b8b9babb",
         15532 => x"bcbdbebf",
         15533 => x"c0c1c2c3",
         15534 => x"c4c5c6c7",
         15535 => x"c8c9cacb",
         15536 => x"cccdcecf",
         15537 => x"d0d1d2d3",
         15538 => x"d4d5d6d7",
         15539 => x"d8d9dadb",
         15540 => x"dcdddedf",
         15541 => x"e0e1e2e3",
         15542 => x"e4e5e6e7",
         15543 => x"e8e9eaeb",
         15544 => x"ecedeeef",
         15545 => x"f0f1f2f3",
         15546 => x"f4f5f6f7",
         15547 => x"f8f9fafb",
         15548 => x"fcfdfeff",
         15549 => x"2b2e2c3b",
         15550 => x"3d5b5d2f",
         15551 => x"5c222a3a",
         15552 => x"3c3e3f7c",
         15553 => x"7f000000",
         15554 => x"00010004",
         15555 => x"00100040",
         15556 => x"01000200",
         15557 => x"00000000",
         15558 => x"00010002",
         15559 => x"00040008",
         15560 => x"00100020",
         15561 => x"00000000",
         15562 => x"00c700fc",
         15563 => x"00e900e2",
         15564 => x"00e400e0",
         15565 => x"00e500e7",
         15566 => x"00ea00eb",
         15567 => x"00e800ef",
         15568 => x"00ee00ec",
         15569 => x"00c400c5",
         15570 => x"00c900e6",
         15571 => x"00c600f4",
         15572 => x"00f600f2",
         15573 => x"00fb00f9",
         15574 => x"00ff00d6",
         15575 => x"00dc00a2",
         15576 => x"00a300a5",
         15577 => x"20a70192",
         15578 => x"00e100ed",
         15579 => x"00f300fa",
         15580 => x"00f100d1",
         15581 => x"00aa00ba",
         15582 => x"00bf2310",
         15583 => x"00ac00bd",
         15584 => x"00bc00a1",
         15585 => x"00ab00bb",
         15586 => x"25912592",
         15587 => x"25932502",
         15588 => x"25242561",
         15589 => x"25622556",
         15590 => x"25552563",
         15591 => x"25512557",
         15592 => x"255d255c",
         15593 => x"255b2510",
         15594 => x"25142534",
         15595 => x"252c251c",
         15596 => x"2500253c",
         15597 => x"255e255f",
         15598 => x"255a2554",
         15599 => x"25692566",
         15600 => x"25602550",
         15601 => x"256c2567",
         15602 => x"25682564",
         15603 => x"25652559",
         15604 => x"25582552",
         15605 => x"2553256b",
         15606 => x"256a2518",
         15607 => x"250c2588",
         15608 => x"2584258c",
         15609 => x"25902580",
         15610 => x"03b100df",
         15611 => x"039303c0",
         15612 => x"03a303c3",
         15613 => x"00b503c4",
         15614 => x"03a60398",
         15615 => x"03a903b4",
         15616 => x"221e03c6",
         15617 => x"03b52229",
         15618 => x"226100b1",
         15619 => x"22652264",
         15620 => x"23202321",
         15621 => x"00f72248",
         15622 => x"00b02219",
         15623 => x"00b7221a",
         15624 => x"207f00b2",
         15625 => x"25a000a0",
         15626 => x"0061031a",
         15627 => x"00e00317",
         15628 => x"00f80307",
         15629 => x"00ff0001",
         15630 => x"01780100",
         15631 => x"01300132",
         15632 => x"01060139",
         15633 => x"0110014a",
         15634 => x"012e0179",
         15635 => x"01060180",
         15636 => x"004d0243",
         15637 => x"01810182",
         15638 => x"01820184",
         15639 => x"01840186",
         15640 => x"01870187",
         15641 => x"0189018a",
         15642 => x"018b018b",
         15643 => x"018d018e",
         15644 => x"018f0190",
         15645 => x"01910191",
         15646 => x"01930194",
         15647 => x"01f60196",
         15648 => x"01970198",
         15649 => x"0198023d",
         15650 => x"019b019c",
         15651 => x"019d0220",
         15652 => x"019f01a0",
         15653 => x"01a001a2",
         15654 => x"01a201a4",
         15655 => x"01a401a6",
         15656 => x"01a701a7",
         15657 => x"01a901aa",
         15658 => x"01ab01ac",
         15659 => x"01ac01ae",
         15660 => x"01af01af",
         15661 => x"01b101b2",
         15662 => x"01b301b3",
         15663 => x"01b501b5",
         15664 => x"01b701b8",
         15665 => x"01b801ba",
         15666 => x"01bb01bc",
         15667 => x"01bc01be",
         15668 => x"01f701c0",
         15669 => x"01c101c2",
         15670 => x"01c301c4",
         15671 => x"01c501c4",
         15672 => x"01c701c8",
         15673 => x"01c701ca",
         15674 => x"01cb01ca",
         15675 => x"01cd0110",
         15676 => x"01dd0001",
         15677 => x"018e01de",
         15678 => x"011201f3",
         15679 => x"000301f1",
         15680 => x"01f401f4",
         15681 => x"01f80128",
         15682 => x"02220112",
         15683 => x"023a0009",
         15684 => x"2c65023b",
         15685 => x"023b023d",
         15686 => x"2c66023f",
         15687 => x"02400241",
         15688 => x"02410246",
         15689 => x"010a0253",
         15690 => x"00400181",
         15691 => x"01860255",
         15692 => x"0189018a",
         15693 => x"0258018f",
         15694 => x"025a0190",
         15695 => x"025c025d",
         15696 => x"025e025f",
         15697 => x"01930261",
         15698 => x"02620194",
         15699 => x"02640265",
         15700 => x"02660267",
         15701 => x"01970196",
         15702 => x"026a2c62",
         15703 => x"026c026d",
         15704 => x"026e019c",
         15705 => x"02700271",
         15706 => x"019d0273",
         15707 => x"0274019f",
         15708 => x"02760277",
         15709 => x"02780279",
         15710 => x"027a027b",
         15711 => x"027c2c64",
         15712 => x"027e027f",
         15713 => x"01a60281",
         15714 => x"028201a9",
         15715 => x"02840285",
         15716 => x"02860287",
         15717 => x"01ae0244",
         15718 => x"01b101b2",
         15719 => x"0245028d",
         15720 => x"028e028f",
         15721 => x"02900291",
         15722 => x"01b7037b",
         15723 => x"000303fd",
         15724 => x"03fe03ff",
         15725 => x"03ac0004",
         15726 => x"03860388",
         15727 => x"0389038a",
         15728 => x"03b10311",
         15729 => x"03c20002",
         15730 => x"03a303a3",
         15731 => x"03c40308",
         15732 => x"03cc0003",
         15733 => x"038c038e",
         15734 => x"038f03d8",
         15735 => x"011803f2",
         15736 => x"000a03f9",
         15737 => x"03f303f4",
         15738 => x"03f503f6",
         15739 => x"03f703f7",
         15740 => x"03f903fa",
         15741 => x"03fa0430",
         15742 => x"03200450",
         15743 => x"07100460",
         15744 => x"0122048a",
         15745 => x"013604c1",
         15746 => x"010e04cf",
         15747 => x"000104c0",
         15748 => x"04d00144",
         15749 => x"05610426",
         15750 => x"00000000",
         15751 => x"1d7d0001",
         15752 => x"2c631e00",
         15753 => x"01961ea0",
         15754 => x"015a1f00",
         15755 => x"06081f10",
         15756 => x"06061f20",
         15757 => x"06081f30",
         15758 => x"06081f40",
         15759 => x"06061f51",
         15760 => x"00071f59",
         15761 => x"1f521f5b",
         15762 => x"1f541f5d",
         15763 => x"1f561f5f",
         15764 => x"1f600608",
         15765 => x"1f70000e",
         15766 => x"1fba1fbb",
         15767 => x"1fc81fc9",
         15768 => x"1fca1fcb",
         15769 => x"1fda1fdb",
         15770 => x"1ff81ff9",
         15771 => x"1fea1feb",
         15772 => x"1ffa1ffb",
         15773 => x"1f800608",
         15774 => x"1f900608",
         15775 => x"1fa00608",
         15776 => x"1fb00004",
         15777 => x"1fb81fb9",
         15778 => x"1fb21fbc",
         15779 => x"1fcc0001",
         15780 => x"1fc31fd0",
         15781 => x"06021fe0",
         15782 => x"06021fe5",
         15783 => x"00011fec",
         15784 => x"1ff30001",
         15785 => x"1ffc214e",
         15786 => x"00012132",
         15787 => x"21700210",
         15788 => x"21840001",
         15789 => x"218324d0",
         15790 => x"051a2c30",
         15791 => x"042f2c60",
         15792 => x"01022c67",
         15793 => x"01062c75",
         15794 => x"01022c80",
         15795 => x"01642d00",
         15796 => x"0826ff41",
         15797 => x"031a0000",
         15798 => x"00000000",
         15799 => x"0000e658",
         15800 => x"01020100",
         15801 => x"00000000",
         15802 => x"00000000",
         15803 => x"0000e660",
         15804 => x"01040100",
         15805 => x"00000000",
         15806 => x"00000000",
         15807 => x"0000e668",
         15808 => x"01140300",
         15809 => x"00000000",
         15810 => x"00000000",
         15811 => x"0000e670",
         15812 => x"012b0300",
         15813 => x"00000000",
         15814 => x"00000000",
         15815 => x"0000e678",
         15816 => x"01300300",
         15817 => x"00000000",
         15818 => x"00000000",
         15819 => x"0000e680",
         15820 => x"013c0400",
         15821 => x"00000000",
         15822 => x"00000000",
         15823 => x"0000e688",
         15824 => x"013d0400",
         15825 => x"00000000",
         15826 => x"00000000",
         15827 => x"0000e690",
         15828 => x"013f0400",
         15829 => x"00000000",
         15830 => x"00000000",
         15831 => x"0000e698",
         15832 => x"01400400",
         15833 => x"00000000",
         15834 => x"00000000",
         15835 => x"0000e6a0",
         15836 => x"01410400",
         15837 => x"00000000",
         15838 => x"00000000",
         15839 => x"0000e6a4",
         15840 => x"01420400",
         15841 => x"00000000",
         15842 => x"00000000",
         15843 => x"0000e6a8",
         15844 => x"01430400",
         15845 => x"00000000",
         15846 => x"00000000",
         15847 => x"0000e6ac",
         15848 => x"01500500",
         15849 => x"00000000",
         15850 => x"00000000",
         15851 => x"0000e6b0",
         15852 => x"01510500",
         15853 => x"00000000",
         15854 => x"00000000",
         15855 => x"0000e6b4",
         15856 => x"01540500",
         15857 => x"00000000",
         15858 => x"00000000",
         15859 => x"0000e6b8",
         15860 => x"01550500",
         15861 => x"00000000",
         15862 => x"00000000",
         15863 => x"0000e6bc",
         15864 => x"01790700",
         15865 => x"00000000",
         15866 => x"00000000",
         15867 => x"0000e6c4",
         15868 => x"01780700",
         15869 => x"00000000",
         15870 => x"00000000",
         15871 => x"0000e6c8",
         15872 => x"01820800",
         15873 => x"00000000",
         15874 => x"00000000",
         15875 => x"0000e6d0",
         15876 => x"01830800",
         15877 => x"00000000",
         15878 => x"00000000",
         15879 => x"0000e6d8",
         15880 => x"01850800",
         15881 => x"00000000",
         15882 => x"00000000",
         15883 => x"0000e6e0",
         15884 => x"01870800",
         15885 => x"00000000",
         15886 => x"00000000",
         15887 => x"0000e6e8",
         15888 => x"01880800",
         15889 => x"00000000",
         15890 => x"00000000",
         15891 => x"0000e6ec",
         15892 => x"01890800",
         15893 => x"00000000",
         15894 => x"00000000",
         15895 => x"0000e6f0",
         15896 => x"018c0900",
         15897 => x"00000000",
         15898 => x"00000000",
         15899 => x"0000e6f8",
         15900 => x"018d0900",
         15901 => x"00000000",
         15902 => x"00000000",
         15903 => x"0000e700",
         15904 => x"018e0900",
         15905 => x"00000000",
         15906 => x"00000000",
         15907 => x"0000e708",
         15908 => x"018f0900",
         15909 => x"00000000",
         15910 => x"00000000",
         15911 => x"00000000",
         15912 => x"00000000",
         15913 => x"00007fff",
         15914 => x"00000000",
         15915 => x"00007fff",
         15916 => x"00010000",
         15917 => x"00007fff",
         15918 => x"00010000",
         15919 => x"00810000",
         15920 => x"01000000",
         15921 => x"017fffff",
         15922 => x"00000000",
         15923 => x"00000000",
         15924 => x"00007800",
         15925 => x"00000000",
         15926 => x"05f5e100",
         15927 => x"05f5e100",
         15928 => x"05f5e100",
         15929 => x"00000000",
         15930 => x"01010101",
         15931 => x"01010101",
         15932 => x"01011001",
         15933 => x"01000000",
         15934 => x"00000000",
         15935 => x"00000000",
         15936 => x"00000000",
         15937 => x"00000000",
         15938 => x"00000000",
         15939 => x"00000000",
         15940 => x"00000000",
         15941 => x"00000000",
         15942 => x"00000000",
         15943 => x"00000000",
         15944 => x"00000000",
         15945 => x"00000000",
         15946 => x"00000000",
         15947 => x"00000000",
         15948 => x"00000000",
         15949 => x"00000000",
         15950 => x"00000000",
         15951 => x"00000000",
         15952 => x"00000000",
         15953 => x"00000000",
         15954 => x"00000000",
         15955 => x"00000000",
         15956 => x"00000000",
         15957 => x"00000000",
         15958 => x"0000f078",
         15959 => x"01000000",
         15960 => x"0000f080",
         15961 => x"01000000",
         15962 => x"0000f088",
         15963 => x"02000000",
         15964 => x"0001fd80",
         15965 => x"1bfc5ffd",
         15966 => x"f03b3a0d",
         15967 => x"797a405b",
         15968 => x"5df0f0f0",
         15969 => x"71727374",
         15970 => x"75767778",
         15971 => x"696a6b6c",
         15972 => x"6d6e6f70",
         15973 => x"61626364",
         15974 => x"65666768",
         15975 => x"31323334",
         15976 => x"35363738",
         15977 => x"5cf32d20",
         15978 => x"30392c2e",
         15979 => x"f67ff3f4",
         15980 => x"f1f23f2f",
         15981 => x"08f0f0f0",
         15982 => x"f0f0f0f0",
         15983 => x"80818283",
         15984 => x"84f0f0f0",
         15985 => x"1bfc58fd",
         15986 => x"f03a3b0d",
         15987 => x"595a405b",
         15988 => x"5df0f0f0",
         15989 => x"51525354",
         15990 => x"55565758",
         15991 => x"494a4b4c",
         15992 => x"4d4e4f50",
         15993 => x"41424344",
         15994 => x"45464748",
         15995 => x"31323334",
         15996 => x"35363738",
         15997 => x"5cf32d20",
         15998 => x"30392c2e",
         15999 => x"f67ff3f4",
         16000 => x"f1f23f2f",
         16001 => x"08f0f0f0",
         16002 => x"f0f0f0f0",
         16003 => x"80818283",
         16004 => x"84f0f0f0",
         16005 => x"1bfc58fd",
         16006 => x"f02b2a0d",
         16007 => x"595a607b",
         16008 => x"7df0f0f0",
         16009 => x"51525354",
         16010 => x"55565758",
         16011 => x"494a4b4c",
         16012 => x"4d4e4f50",
         16013 => x"41424344",
         16014 => x"45464748",
         16015 => x"21222324",
         16016 => x"25262728",
         16017 => x"7c7e3d20",
         16018 => x"20293c3e",
         16019 => x"f7e2e0e1",
         16020 => x"f9f83f2f",
         16021 => x"fbf0f0f0",
         16022 => x"f0f0f0f0",
         16023 => x"85868788",
         16024 => x"89f0f0f0",
         16025 => x"1bfe1efa",
         16026 => x"f0f0f0f0",
         16027 => x"191a001b",
         16028 => x"1df0f0f0",
         16029 => x"11121314",
         16030 => x"15161718",
         16031 => x"090a0b0c",
         16032 => x"0d0e0f10",
         16033 => x"01020304",
         16034 => x"05060708",
         16035 => x"f0f0f0f0",
         16036 => x"f0f0f0f0",
         16037 => x"f01ef0f0",
         16038 => x"f01ff0f0",
         16039 => x"f0f0f0f0",
         16040 => x"f0f0f01c",
         16041 => x"f0f0f0f0",
         16042 => x"f0f0f0f0",
         16043 => x"80818283",
         16044 => x"84f0f0f0",
         16045 => x"bff0cfc9",
         16046 => x"f0b54dcd",
         16047 => x"3577d7b3",
         16048 => x"b7f0f0f0",
         16049 => x"7c704131",
         16050 => x"39a678dd",
         16051 => x"3d5d6c56",
         16052 => x"1d33d5b1",
         16053 => x"466ed948",
         16054 => x"74434c73",
         16055 => x"3f367e3b",
         16056 => x"7a1e5fa2",
         16057 => x"d39fd100",
         16058 => x"9da3d0b9",
         16059 => x"c6c5c2c1",
         16060 => x"c3c4bbbe",
         16061 => x"f0f0f0f0",
         16062 => x"f0f0f0f0",
         16063 => x"80818283",
         16064 => x"84f0f0f0",
         16065 => x"00000000",
         16066 => x"00000000",
         16067 => x"00000000",
         16068 => x"00000000",
         16069 => x"00000000",
         16070 => x"00000000",
         16071 => x"00000000",
         16072 => x"00000000",
         16073 => x"00000000",
         16074 => x"00000000",
         16075 => x"00000000",
         16076 => x"00000000",
         16077 => x"00000000",
         16078 => x"00000000",
         16079 => x"00000000",
         16080 => x"00000000",
         16081 => x"00000000",
         16082 => x"00000000",
         16083 => x"00000000",
         16084 => x"00000000",
         16085 => x"00000000",
         16086 => x"00000000",
         16087 => x"00000000",
         16088 => x"00000000",
         16089 => x"00000000",
         16090 => x"00010000",
         16091 => x"00000000",
         16092 => x"f8000000",
         16093 => x"0000f0cc",
         16094 => x"f3000000",
         16095 => x"0000f0d4",
         16096 => x"f4000000",
         16097 => x"0000f0d8",
         16098 => x"f1000000",
         16099 => x"0000f0dc",
         16100 => x"f2000000",
         16101 => x"0000f0e0",
         16102 => x"80000000",
         16103 => x"0000f0e4",
         16104 => x"81000000",
         16105 => x"0000f0ec",
         16106 => x"82000000",
         16107 => x"0000f0f4",
         16108 => x"83000000",
         16109 => x"0000f0fc",
         16110 => x"84000000",
         16111 => x"0000f104",
         16112 => x"85000000",
         16113 => x"0000f10c",
         16114 => x"86000000",
         16115 => x"0000f114",
         16116 => x"87000000",
         16117 => x"0000f11c",
         16118 => x"88000000",
         16119 => x"0000f124",
         16120 => x"89000000",
         16121 => x"0000f12c",
         16122 => x"f6000000",
         16123 => x"0000f134",
         16124 => x"7f000000",
         16125 => x"0000f13c",
         16126 => x"f9000000",
         16127 => x"0000f144",
         16128 => x"e0000000",
         16129 => x"0000f148",
         16130 => x"e1000000",
         16131 => x"0000f150",
         16132 => x"71000000",
         16133 => x"00000000",
         16134 => x"00000000",
         16135 => x"00000000",
         16136 => x"00000000",
         16137 => x"00000000",
         16138 => x"00000000",
         16139 => x"00000000",
         16140 => x"00000000",
         16141 => x"00000000",
         16142 => x"00000000",
         16143 => x"00000000",
         16144 => x"00000000",
         16145 => x"00000000",
         16146 => x"00000000",
         16147 => x"00000000",
         16148 => x"00000000",
         16149 => x"00000000",
         16150 => x"00000000",
         16151 => x"00000000",
         16152 => x"00000000",
         16153 => x"00000000",
         16154 => x"00000000",
         16155 => x"00000000",
         16156 => x"00000000",
         16157 => x"00000000",
         16158 => x"00000000",
         16159 => x"00000000",
         16160 => x"00000000",
         16161 => x"00000000",
         16162 => x"00000000",
         16163 => x"00000000",
         16164 => x"00000000",
         16165 => x"00000000",
         16166 => x"00000000",
         16167 => x"00000000",
         16168 => x"00000000",
         16169 => x"00000000",
         16170 => x"00000000",
         16171 => x"00000000",
         16172 => x"00000000",
         16173 => x"00000000",
         16174 => x"00000000",
         16175 => x"00000000",
         16176 => x"00000000",
         16177 => x"00000000",
         16178 => x"00000000",
         16179 => x"00000000",
         16180 => x"00000000",
         16181 => x"00000000",
         16182 => x"00000000",
         16183 => x"00000000",
         16184 => x"00000000",
         16185 => x"00000000",
         16186 => x"00000000",
         16187 => x"00000000",
         16188 => x"00000000",
         16189 => x"00000000",
         16190 => x"00000000",
         16191 => x"00000000",
         16192 => x"00000000",
         16193 => x"00000000",
         16194 => x"00000000",
         16195 => x"00000000",
         16196 => x"00000000",
         16197 => x"00000000",
         16198 => x"00000000",
         16199 => x"00000000",
         16200 => x"00000000",
         16201 => x"00000000",
         16202 => x"00000000",
         16203 => x"00000000",
         16204 => x"00000000",
         16205 => x"00000000",
         16206 => x"00000000",
         16207 => x"00000000",
         16208 => x"00000000",
         16209 => x"00000000",
         16210 => x"00000000",
         16211 => x"00000000",
         16212 => x"00000000",
         16213 => x"00000000",
         16214 => x"00000000",
         16215 => x"00000000",
         16216 => x"00000000",
         16217 => x"00000000",
         16218 => x"00000000",
         16219 => x"00000000",
         16220 => x"00000000",
         16221 => x"00000000",
         16222 => x"00000000",
         16223 => x"00000000",
         16224 => x"00000000",
         16225 => x"00000000",
         16226 => x"00000000",
         16227 => x"00000000",
         16228 => x"00000000",
         16229 => x"00000000",
         16230 => x"00000000",
         16231 => x"00000000",
         16232 => x"00000000",
         16233 => x"00000000",
         16234 => x"00000000",
         16235 => x"00000000",
         16236 => x"00000000",
         16237 => x"00000000",
         16238 => x"00000000",
         16239 => x"00000000",
         16240 => x"00000000",
         16241 => x"00000000",
         16242 => x"00000000",
         16243 => x"00000000",
         16244 => x"00000000",
         16245 => x"00000000",
         16246 => x"00000000",
         16247 => x"00000000",
         16248 => x"00000000",
         16249 => x"00000000",
         16250 => x"00000000",
         16251 => x"00000000",
         16252 => x"00000000",
         16253 => x"00000000",
         16254 => x"00000000",
         16255 => x"00000000",
         16256 => x"00000000",
         16257 => x"00000000",
         16258 => x"00000000",
         16259 => x"00000000",
         16260 => x"00000000",
         16261 => x"00000000",
         16262 => x"00000000",
         16263 => x"00000000",
         16264 => x"00000000",
         16265 => x"00000000",
         16266 => x"00000000",
         16267 => x"00000000",
         16268 => x"00000000",
         16269 => x"00000000",
         16270 => x"00000000",
         16271 => x"00000000",
         16272 => x"00000000",
         16273 => x"00000000",
         16274 => x"00000000",
         16275 => x"00000000",
         16276 => x"00000000",
         16277 => x"00000000",
         16278 => x"00000000",
         16279 => x"00000000",
         16280 => x"00000000",
         16281 => x"00000000",
         16282 => x"00000000",
         16283 => x"00000000",
         16284 => x"00000000",
         16285 => x"00000000",
         16286 => x"00000000",
         16287 => x"00000000",
         16288 => x"00000000",
         16289 => x"00000000",
         16290 => x"00000000",
         16291 => x"00000000",
         16292 => x"00000000",
         16293 => x"00000000",
         16294 => x"00000000",
         16295 => x"00000000",
         16296 => x"00000000",
         16297 => x"00000000",
         16298 => x"00000000",
         16299 => x"00000000",
         16300 => x"00000000",
         16301 => x"00000000",
         16302 => x"00000000",
         16303 => x"00000000",
         16304 => x"00000000",
         16305 => x"00000000",
         16306 => x"00000000",
         16307 => x"00000000",
         16308 => x"00000000",
         16309 => x"00000000",
         16310 => x"00000000",
         16311 => x"00000000",
         16312 => x"00000000",
         16313 => x"00000000",
         16314 => x"00000000",
         16315 => x"00000000",
         16316 => x"00000000",
         16317 => x"00000000",
         16318 => x"00000000",
         16319 => x"00000000",
         16320 => x"00000000",
         16321 => x"00000000",
         16322 => x"00000000",
         16323 => x"00000000",
         16324 => x"00000000",
         16325 => x"00000000",
         16326 => x"00000000",
         16327 => x"00000000",
         16328 => x"00000000",
         16329 => x"00000000",
         16330 => x"00000000",
         16331 => x"00000000",
         16332 => x"00000000",
         16333 => x"00000000",
         16334 => x"00000000",
         16335 => x"00000000",
         16336 => x"00000000",
         16337 => x"00000000",
         16338 => x"00000000",
         16339 => x"00000000",
         16340 => x"00000000",
         16341 => x"00000000",
         16342 => x"00000000",
         16343 => x"00000000",
         16344 => x"00000000",
         16345 => x"00000000",
         16346 => x"00000000",
         16347 => x"00000000",
         16348 => x"00000000",
         16349 => x"00000000",
         16350 => x"00000000",
         16351 => x"00000000",
         16352 => x"00000000",
         16353 => x"00000000",
         16354 => x"00000000",
         16355 => x"00000000",
         16356 => x"00000000",
         16357 => x"00000000",
         16358 => x"00000000",
         16359 => x"00000000",
         16360 => x"00000000",
         16361 => x"00000000",
         16362 => x"00000000",
         16363 => x"00000000",
         16364 => x"00000000",
         16365 => x"00000000",
         16366 => x"00000000",
         16367 => x"00000000",
         16368 => x"00000000",
         16369 => x"00000000",
         16370 => x"00000000",
         16371 => x"00000000",
         16372 => x"00000000",
         16373 => x"00000000",
         16374 => x"00000000",
         16375 => x"00000000",
         16376 => x"00000000",
         16377 => x"00000000",
         16378 => x"00000000",
         16379 => x"00000000",
         16380 => x"00000000",
         16381 => x"00000000",
         16382 => x"00000000",
         16383 => x"00000000",
         16384 => x"00000000",
         16385 => x"00000000",
         16386 => x"00000000",
         16387 => x"00000000",
         16388 => x"00000000",
         16389 => x"00000000",
         16390 => x"00000000",
         16391 => x"00000000",
         16392 => x"00000000",
         16393 => x"00000000",
         16394 => x"00000000",
         16395 => x"00000000",
         16396 => x"00000000",
         16397 => x"00000000",
         16398 => x"00000000",
         16399 => x"00000000",
         16400 => x"00000000",
         16401 => x"00000000",
         16402 => x"00000000",
         16403 => x"00000000",
         16404 => x"00000000",
         16405 => x"00000000",
         16406 => x"00000000",
         16407 => x"00000000",
         16408 => x"00000000",
         16409 => x"00000000",
         16410 => x"00000000",
         16411 => x"00000000",
         16412 => x"00000000",
         16413 => x"00000000",
         16414 => x"00000000",
         16415 => x"00000000",
         16416 => x"00000000",
         16417 => x"00000000",
         16418 => x"00000000",
         16419 => x"00000000",
         16420 => x"00000000",
         16421 => x"00000000",
         16422 => x"00000000",
         16423 => x"00000000",
         16424 => x"00000000",
         16425 => x"00000000",
         16426 => x"00000000",
         16427 => x"00000000",
         16428 => x"00000000",
         16429 => x"00000000",
         16430 => x"00000000",
         16431 => x"00000000",
         16432 => x"00000000",
         16433 => x"00000000",
         16434 => x"00000000",
         16435 => x"00000000",
         16436 => x"00000000",
         16437 => x"00000000",
         16438 => x"00000000",
         16439 => x"00000000",
         16440 => x"00000000",
         16441 => x"00000000",
         16442 => x"00000000",
         16443 => x"00000000",
         16444 => x"00000000",
         16445 => x"00000000",
         16446 => x"00000000",
         16447 => x"00000000",
         16448 => x"00000000",
         16449 => x"00000000",
         16450 => x"00000000",
         16451 => x"00000000",
         16452 => x"00000000",
         16453 => x"00000000",
         16454 => x"00000000",
         16455 => x"00000000",
         16456 => x"00000000",
         16457 => x"00000000",
         16458 => x"00000000",
         16459 => x"00000000",
         16460 => x"00000000",
         16461 => x"00000000",
         16462 => x"00000000",
         16463 => x"00000000",
         16464 => x"00000000",
         16465 => x"00000000",
         16466 => x"00000000",
         16467 => x"00000000",
         16468 => x"00000000",
         16469 => x"00000000",
         16470 => x"00000000",
         16471 => x"00000000",
         16472 => x"00000000",
         16473 => x"00000000",
         16474 => x"00000000",
         16475 => x"00000000",
         16476 => x"00000000",
         16477 => x"00000000",
         16478 => x"00000000",
         16479 => x"00000000",
         16480 => x"00000000",
         16481 => x"00000000",
         16482 => x"00000000",
         16483 => x"00000000",
         16484 => x"00000000",
         16485 => x"00000000",
         16486 => x"00000000",
         16487 => x"00000000",
         16488 => x"00000000",
         16489 => x"00000000",
         16490 => x"00000000",
         16491 => x"00000000",
         16492 => x"00000000",
         16493 => x"00000000",
         16494 => x"00000000",
         16495 => x"00000000",
         16496 => x"00000000",
         16497 => x"00000000",
         16498 => x"00000000",
         16499 => x"00000000",
         16500 => x"00000000",
         16501 => x"00000000",
         16502 => x"00000000",
         16503 => x"00000000",
         16504 => x"00000000",
         16505 => x"00000000",
         16506 => x"00000000",
         16507 => x"00000000",
         16508 => x"00000000",
         16509 => x"00000000",
         16510 => x"00000000",
         16511 => x"00000000",
         16512 => x"00000000",
         16513 => x"00000000",
         16514 => x"00000000",
         16515 => x"00000000",
         16516 => x"00000000",
         16517 => x"00000000",
         16518 => x"00000000",
         16519 => x"00000000",
         16520 => x"00000000",
         16521 => x"00000000",
         16522 => x"00000000",
         16523 => x"00000000",
         16524 => x"00000000",
         16525 => x"00000000",
         16526 => x"00000000",
         16527 => x"00000000",
         16528 => x"00000000",
         16529 => x"00000000",
         16530 => x"00000000",
         16531 => x"00000000",
         16532 => x"00000000",
         16533 => x"00000000",
         16534 => x"00000000",
         16535 => x"00000000",
         16536 => x"00000000",
         16537 => x"00000000",
         16538 => x"00000000",
         16539 => x"00000000",
         16540 => x"00000000",
         16541 => x"00000000",
         16542 => x"00000000",
         16543 => x"00000000",
         16544 => x"00000000",
         16545 => x"00000000",
         16546 => x"00000000",
         16547 => x"00000000",
         16548 => x"00000000",
         16549 => x"00000000",
         16550 => x"00000000",
         16551 => x"00000000",
         16552 => x"00000000",
         16553 => x"00000000",
         16554 => x"00000000",
         16555 => x"00000000",
         16556 => x"00000000",
         16557 => x"00000000",
         16558 => x"00000000",
         16559 => x"00000000",
         16560 => x"00000000",
         16561 => x"00000000",
         16562 => x"00000000",
         16563 => x"00000000",
         16564 => x"00000000",
         16565 => x"00000000",
         16566 => x"00000000",
         16567 => x"00000000",
         16568 => x"00000000",
         16569 => x"00000000",
         16570 => x"00000000",
         16571 => x"00000000",
         16572 => x"00000000",
         16573 => x"00000000",
         16574 => x"00000000",
         16575 => x"00000000",
         16576 => x"00000000",
         16577 => x"00000000",
         16578 => x"00000000",
         16579 => x"00000000",
         16580 => x"00000000",
         16581 => x"00000000",
         16582 => x"00000000",
         16583 => x"00000000",
         16584 => x"00000000",
         16585 => x"00000000",
         16586 => x"00000000",
         16587 => x"00000000",
         16588 => x"00000000",
         16589 => x"00000000",
         16590 => x"00000000",
         16591 => x"00000000",
         16592 => x"00000000",
         16593 => x"00000000",
         16594 => x"00000000",
         16595 => x"00000000",
         16596 => x"00000000",
         16597 => x"00000000",
         16598 => x"00000000",
         16599 => x"00000000",
         16600 => x"00000000",
         16601 => x"00000000",
         16602 => x"00000000",
         16603 => x"00000000",
         16604 => x"00000000",
         16605 => x"00000000",
         16606 => x"00000000",
         16607 => x"00000000",
         16608 => x"00000000",
         16609 => x"00000000",
         16610 => x"00000000",
         16611 => x"00000000",
         16612 => x"00000000",
         16613 => x"00000000",
         16614 => x"00000000",
         16615 => x"00000000",
         16616 => x"00000000",
         16617 => x"00000000",
         16618 => x"00000000",
         16619 => x"00000000",
         16620 => x"00000000",
         16621 => x"00000000",
         16622 => x"00000000",
         16623 => x"00000000",
         16624 => x"00000000",
         16625 => x"00000000",
         16626 => x"00000000",
         16627 => x"00000000",
         16628 => x"00000000",
         16629 => x"00000000",
         16630 => x"00000000",
         16631 => x"00000000",
         16632 => x"00000000",
         16633 => x"00000000",
         16634 => x"00000000",
         16635 => x"00000000",
         16636 => x"00000000",
         16637 => x"00000000",
         16638 => x"00000000",
         16639 => x"00000000",
         16640 => x"00000000",
         16641 => x"00000000",
         16642 => x"00000000",
         16643 => x"00000000",
         16644 => x"00000000",
         16645 => x"00000000",
         16646 => x"00000000",
         16647 => x"00000000",
         16648 => x"00000000",
         16649 => x"00000000",
         16650 => x"00000000",
         16651 => x"00000000",
         16652 => x"00000000",
         16653 => x"00000000",
         16654 => x"00000000",
         16655 => x"00000000",
         16656 => x"00000000",
         16657 => x"00000000",
         16658 => x"00000000",
         16659 => x"00000000",
         16660 => x"00000000",
         16661 => x"00000000",
         16662 => x"00000000",
         16663 => x"00000000",
         16664 => x"00000000",
         16665 => x"00000000",
         16666 => x"00000000",
         16667 => x"00000000",
         16668 => x"00000000",
         16669 => x"00000000",
         16670 => x"00000000",
         16671 => x"00000000",
         16672 => x"00000000",
         16673 => x"00000000",
         16674 => x"00000000",
         16675 => x"00000000",
         16676 => x"00000000",
         16677 => x"00000000",
         16678 => x"00000000",
         16679 => x"00000000",
         16680 => x"00000000",
         16681 => x"00000000",
         16682 => x"00000000",
         16683 => x"00000000",
         16684 => x"00000000",
         16685 => x"00000000",
         16686 => x"00000000",
         16687 => x"00000000",
         16688 => x"00000000",
         16689 => x"00000000",
         16690 => x"00000000",
         16691 => x"00000000",
         16692 => x"00000000",
         16693 => x"00000000",
         16694 => x"00000000",
         16695 => x"00000000",
         16696 => x"00000000",
         16697 => x"00000000",
         16698 => x"00000000",
         16699 => x"00000000",
         16700 => x"00000000",
         16701 => x"00000000",
         16702 => x"00000000",
         16703 => x"00000000",
         16704 => x"00000000",
         16705 => x"00000000",
         16706 => x"00000000",
         16707 => x"00000000",
         16708 => x"00000000",
         16709 => x"00000000",
         16710 => x"00000000",
         16711 => x"00000000",
         16712 => x"00000000",
         16713 => x"00000000",
         16714 => x"00000000",
         16715 => x"00000000",
         16716 => x"00000000",
         16717 => x"00000000",
         16718 => x"00000000",
         16719 => x"00000000",
         16720 => x"00000000",
         16721 => x"00000000",
         16722 => x"00000000",
         16723 => x"00000000",
         16724 => x"00000000",
         16725 => x"00000000",
         16726 => x"00000000",
         16727 => x"00000000",
         16728 => x"00000000",
         16729 => x"00000000",
         16730 => x"00000000",
         16731 => x"00000000",
         16732 => x"00000000",
         16733 => x"00000000",
         16734 => x"00000000",
         16735 => x"00000000",
         16736 => x"00000000",
         16737 => x"00000000",
         16738 => x"00000000",
         16739 => x"00000000",
         16740 => x"00000000",
         16741 => x"00000000",
         16742 => x"00000000",
         16743 => x"00000000",
         16744 => x"00000000",
         16745 => x"00000000",
         16746 => x"00000000",
         16747 => x"00000000",
         16748 => x"00000000",
         16749 => x"00000000",
         16750 => x"00000000",
         16751 => x"00000000",
         16752 => x"00000000",
         16753 => x"00000000",
         16754 => x"00000000",
         16755 => x"00000000",
         16756 => x"00000000",
         16757 => x"00000000",
         16758 => x"00000000",
         16759 => x"00000000",
         16760 => x"00000000",
         16761 => x"00000000",
         16762 => x"00000000",
         16763 => x"00000000",
         16764 => x"00000000",
         16765 => x"00000000",
         16766 => x"00000000",
         16767 => x"00000000",
         16768 => x"00000000",
         16769 => x"00000000",
         16770 => x"00000000",
         16771 => x"00000000",
         16772 => x"00000000",
         16773 => x"00000000",
         16774 => x"00000000",
         16775 => x"00000000",
         16776 => x"00000000",
         16777 => x"00000000",
         16778 => x"00000000",
         16779 => x"00000000",
         16780 => x"00000000",
         16781 => x"00000000",
         16782 => x"00000000",
         16783 => x"00000000",
         16784 => x"00000000",
         16785 => x"00000000",
         16786 => x"00000000",
         16787 => x"00000000",
         16788 => x"00000000",
         16789 => x"00000000",
         16790 => x"00000000",
         16791 => x"00000000",
         16792 => x"00000000",
         16793 => x"00000000",
         16794 => x"00000000",
         16795 => x"00000000",
         16796 => x"00000000",
         16797 => x"00000000",
         16798 => x"00000000",
         16799 => x"00000000",
         16800 => x"00000000",
         16801 => x"00000000",
         16802 => x"00000000",
         16803 => x"00000000",
         16804 => x"00000000",
         16805 => x"00000000",
         16806 => x"00000000",
         16807 => x"00000000",
         16808 => x"00000000",
         16809 => x"00000000",
         16810 => x"00000000",
         16811 => x"00000000",
         16812 => x"00000000",
         16813 => x"00000000",
         16814 => x"00000000",
         16815 => x"00000000",
         16816 => x"00000000",
         16817 => x"00000000",
         16818 => x"00000000",
         16819 => x"00000000",
         16820 => x"00000000",
         16821 => x"00000000",
         16822 => x"00000000",
         16823 => x"00000000",
         16824 => x"00000000",
         16825 => x"00000000",
         16826 => x"00000000",
         16827 => x"00000000",
         16828 => x"00000000",
         16829 => x"00000000",
         16830 => x"00000000",
         16831 => x"00000000",
         16832 => x"00000000",
         16833 => x"00000000",
         16834 => x"00000000",
         16835 => x"00000000",
         16836 => x"00000000",
         16837 => x"00000000",
         16838 => x"00000000",
         16839 => x"00000000",
         16840 => x"00000000",
         16841 => x"00000000",
         16842 => x"00000000",
         16843 => x"00000000",
         16844 => x"00000000",
         16845 => x"00000000",
         16846 => x"00000000",
         16847 => x"00000000",
         16848 => x"00000000",
         16849 => x"00000000",
         16850 => x"00000000",
         16851 => x"00000000",
         16852 => x"00000000",
         16853 => x"00000000",
         16854 => x"00000000",
         16855 => x"00000000",
         16856 => x"00000000",
         16857 => x"00000000",
         16858 => x"00000000",
         16859 => x"00000000",
         16860 => x"00000000",
         16861 => x"00000000",
         16862 => x"00000000",
         16863 => x"00000000",
         16864 => x"00000000",
         16865 => x"00000000",
         16866 => x"00000000",
         16867 => x"00000000",
         16868 => x"00000000",
         16869 => x"00000000",
         16870 => x"00000000",
         16871 => x"00000000",
         16872 => x"00000000",
         16873 => x"00000000",
         16874 => x"00000000",
         16875 => x"00000000",
         16876 => x"00000000",
         16877 => x"00000000",
         16878 => x"00000000",
         16879 => x"00000000",
         16880 => x"00000000",
         16881 => x"00000000",
         16882 => x"00000000",
         16883 => x"00000000",
         16884 => x"00000000",
         16885 => x"00000000",
         16886 => x"00000000",
         16887 => x"00000000",
         16888 => x"00000000",
         16889 => x"00000000",
         16890 => x"00000000",
         16891 => x"00000000",
         16892 => x"00000000",
         16893 => x"00000000",
         16894 => x"00000000",
         16895 => x"00000000",
         16896 => x"00000000",
         16897 => x"00000000",
         16898 => x"00000000",
         16899 => x"00000000",
         16900 => x"00000000",
         16901 => x"00000000",
         16902 => x"00000000",
         16903 => x"00000000",
         16904 => x"00000000",
         16905 => x"00000000",
         16906 => x"00000000",
         16907 => x"00000000",
         16908 => x"00000000",
         16909 => x"00000000",
         16910 => x"00000000",
         16911 => x"00000000",
         16912 => x"00000000",
         16913 => x"00000000",
         16914 => x"00000000",
         16915 => x"00000000",
         16916 => x"00000000",
         16917 => x"00000000",
         16918 => x"00000000",
         16919 => x"00000000",
         16920 => x"00000000",
         16921 => x"00000000",
         16922 => x"00000000",
         16923 => x"00000000",
         16924 => x"00000000",
         16925 => x"00000000",
         16926 => x"00000000",
         16927 => x"00000000",
         16928 => x"00000000",
         16929 => x"00000000",
         16930 => x"00000000",
         16931 => x"00000000",
         16932 => x"00000000",
         16933 => x"00000000",
         16934 => x"00000000",
         16935 => x"00000000",
         16936 => x"00000000",
         16937 => x"00000000",
         16938 => x"00000000",
         16939 => x"00000000",
         16940 => x"00000000",
         16941 => x"00000000",
         16942 => x"00000000",
         16943 => x"00000000",
         16944 => x"00000000",
         16945 => x"00000000",
         16946 => x"00000000",
         16947 => x"00000000",
         16948 => x"00000000",
         16949 => x"00000000",
         16950 => x"00000000",
         16951 => x"00000000",
         16952 => x"00000000",
         16953 => x"00000000",
         16954 => x"00000000",
         16955 => x"00000000",
         16956 => x"00000000",
         16957 => x"00000000",
         16958 => x"00000000",
         16959 => x"00000000",
         16960 => x"00000000",
         16961 => x"00000000",
         16962 => x"00000000",
         16963 => x"00000000",
         16964 => x"00000000",
         16965 => x"00000000",
         16966 => x"00000000",
         16967 => x"00000000",
         16968 => x"00000000",
         16969 => x"00000000",
         16970 => x"00000000",
         16971 => x"00000000",
         16972 => x"00000000",
         16973 => x"00000000",
         16974 => x"00000000",
         16975 => x"00000000",
         16976 => x"00000000",
         16977 => x"00000000",
         16978 => x"00000000",
         16979 => x"00000000",
         16980 => x"00000000",
         16981 => x"00000000",
         16982 => x"00000000",
         16983 => x"00000000",
         16984 => x"00000000",
         16985 => x"00000000",
         16986 => x"00000000",
         16987 => x"00000000",
         16988 => x"00000000",
         16989 => x"00000000",
         16990 => x"00000000",
         16991 => x"00000000",
         16992 => x"00000000",
         16993 => x"00000000",
         16994 => x"00000000",
         16995 => x"00000000",
         16996 => x"00000000",
         16997 => x"00000000",
         16998 => x"00000000",
         16999 => x"00000000",
         17000 => x"00000000",
         17001 => x"00000000",
         17002 => x"00000000",
         17003 => x"00000000",
         17004 => x"00000000",
         17005 => x"00000000",
         17006 => x"00000000",
         17007 => x"00000000",
         17008 => x"00000000",
         17009 => x"00000000",
         17010 => x"00000000",
         17011 => x"00000000",
         17012 => x"00000000",
         17013 => x"00000000",
         17014 => x"00000000",
         17015 => x"00000000",
         17016 => x"00000000",
         17017 => x"00000000",
         17018 => x"00000000",
         17019 => x"00000000",
         17020 => x"00000000",
         17021 => x"00000000",
         17022 => x"00000000",
         17023 => x"00000000",
         17024 => x"00000000",
         17025 => x"00000000",
         17026 => x"00000000",
         17027 => x"00000000",
         17028 => x"00000000",
         17029 => x"00000000",
         17030 => x"00000000",
         17031 => x"00000000",
         17032 => x"00000000",
         17033 => x"00000000",
         17034 => x"00000000",
         17035 => x"00000000",
         17036 => x"00000000",
         17037 => x"00000000",
         17038 => x"00000000",
         17039 => x"00000000",
         17040 => x"00000000",
         17041 => x"00000000",
         17042 => x"00000000",
         17043 => x"00000000",
         17044 => x"00000000",
         17045 => x"00000000",
         17046 => x"00000000",
         17047 => x"00000000",
         17048 => x"00000000",
         17049 => x"00000000",
         17050 => x"00000000",
         17051 => x"00000000",
         17052 => x"00000000",
         17053 => x"00000000",
         17054 => x"00000000",
         17055 => x"00000000",
         17056 => x"00000000",
         17057 => x"00000000",
         17058 => x"00000000",
         17059 => x"00000000",
         17060 => x"00000000",
         17061 => x"00000000",
         17062 => x"00000000",
         17063 => x"00000000",
         17064 => x"00000000",
         17065 => x"00000000",
         17066 => x"00000000",
         17067 => x"00000000",
         17068 => x"00000000",
         17069 => x"00000000",
         17070 => x"00000000",
         17071 => x"00000000",
         17072 => x"00000000",
         17073 => x"00000000",
         17074 => x"00000000",
         17075 => x"00000000",
         17076 => x"00000000",
         17077 => x"00000000",
         17078 => x"00000000",
         17079 => x"00000000",
         17080 => x"00000000",
         17081 => x"00000000",
         17082 => x"00000000",
         17083 => x"00000000",
         17084 => x"00000000",
         17085 => x"00000000",
         17086 => x"00000000",
         17087 => x"00000000",
         17088 => x"00000000",
         17089 => x"00000000",
         17090 => x"00000000",
         17091 => x"00000000",
         17092 => x"00000000",
         17093 => x"00000000",
         17094 => x"00000000",
         17095 => x"00000000",
         17096 => x"00000000",
         17097 => x"00000000",
         17098 => x"00000000",
         17099 => x"00000000",
         17100 => x"00000000",
         17101 => x"00000000",
         17102 => x"00000000",
         17103 => x"00000000",
         17104 => x"00000000",
         17105 => x"00000000",
         17106 => x"00000000",
         17107 => x"00000000",
         17108 => x"00000000",
         17109 => x"00000000",
         17110 => x"00000000",
         17111 => x"00000000",
         17112 => x"00000000",
         17113 => x"00000000",
         17114 => x"00000000",
         17115 => x"00000000",
         17116 => x"00000000",
         17117 => x"00000000",
         17118 => x"00000000",
         17119 => x"00000000",
         17120 => x"00000000",
         17121 => x"00000000",
         17122 => x"00000000",
         17123 => x"00000000",
         17124 => x"00000000",
         17125 => x"00000000",
         17126 => x"00000000",
         17127 => x"00000000",
         17128 => x"00000000",
         17129 => x"00000000",
         17130 => x"00000000",
         17131 => x"00000000",
         17132 => x"00000000",
         17133 => x"00000000",
         17134 => x"00000000",
         17135 => x"00000000",
         17136 => x"00000000",
         17137 => x"00000000",
         17138 => x"00000000",
         17139 => x"00000000",
         17140 => x"00000000",
         17141 => x"00000000",
         17142 => x"00000000",
         17143 => x"00000000",
         17144 => x"00000000",
         17145 => x"00000000",
         17146 => x"00000000",
         17147 => x"00000000",
         17148 => x"00000000",
         17149 => x"00000000",
         17150 => x"00000000",
         17151 => x"00000000",
         17152 => x"00000000",
         17153 => x"00000000",
         17154 => x"00000000",
         17155 => x"00000000",
         17156 => x"00000000",
         17157 => x"00000000",
         17158 => x"00000000",
         17159 => x"00000000",
         17160 => x"00000000",
         17161 => x"00000000",
         17162 => x"00000000",
         17163 => x"00000000",
         17164 => x"00000000",
         17165 => x"00000000",
         17166 => x"00000000",
         17167 => x"00000000",
         17168 => x"00000000",
         17169 => x"00000000",
         17170 => x"00000000",
         17171 => x"00000000",
         17172 => x"00000000",
         17173 => x"00000000",
         17174 => x"00000000",
         17175 => x"00000000",
         17176 => x"00000000",
         17177 => x"00000000",
         17178 => x"00000000",
         17179 => x"00000000",
         17180 => x"00000000",
         17181 => x"00000000",
         17182 => x"00000000",
         17183 => x"00000000",
         17184 => x"00000000",
         17185 => x"00000000",
         17186 => x"00000000",
         17187 => x"00000000",
         17188 => x"00000000",
         17189 => x"00000000",
         17190 => x"00000000",
         17191 => x"00000000",
         17192 => x"00000000",
         17193 => x"00000000",
         17194 => x"00000000",
         17195 => x"00000000",
         17196 => x"00000000",
         17197 => x"00000000",
         17198 => x"00000000",
         17199 => x"00000000",
         17200 => x"00000000",
         17201 => x"00000000",
         17202 => x"00000000",
         17203 => x"00000000",
         17204 => x"00000000",
         17205 => x"00000000",
         17206 => x"00000000",
         17207 => x"00000000",
         17208 => x"00000000",
         17209 => x"00000000",
         17210 => x"00000000",
         17211 => x"00000000",
         17212 => x"00000000",
         17213 => x"00000000",
         17214 => x"00000000",
         17215 => x"00000000",
         17216 => x"00000000",
         17217 => x"00000000",
         17218 => x"00000000",
         17219 => x"00000000",
         17220 => x"00000000",
         17221 => x"00000000",
         17222 => x"00000000",
         17223 => x"00000000",
         17224 => x"00000000",
         17225 => x"00000000",
         17226 => x"00000000",
         17227 => x"00000000",
         17228 => x"00000000",
         17229 => x"00000000",
         17230 => x"00000000",
         17231 => x"00000000",
         17232 => x"00000000",
         17233 => x"00000000",
         17234 => x"00000000",
         17235 => x"00000000",
         17236 => x"00000000",
         17237 => x"00000000",
         17238 => x"00000000",
         17239 => x"00000000",
         17240 => x"00000000",
         17241 => x"00000000",
         17242 => x"00000000",
         17243 => x"00000000",
         17244 => x"00000000",
         17245 => x"00000000",
         17246 => x"00000000",
         17247 => x"00000000",
         17248 => x"00000000",
         17249 => x"00000000",
         17250 => x"00000000",
         17251 => x"00000000",
         17252 => x"00000000",
         17253 => x"00000000",
         17254 => x"00000000",
         17255 => x"00000000",
         17256 => x"00000000",
         17257 => x"00000000",
         17258 => x"00000000",
         17259 => x"00000000",
         17260 => x"00000000",
         17261 => x"00000000",
         17262 => x"00000000",
         17263 => x"00000000",
         17264 => x"00000000",
         17265 => x"00000000",
         17266 => x"00000000",
         17267 => x"00000000",
         17268 => x"00000000",
         17269 => x"00000000",
         17270 => x"00000000",
         17271 => x"00000000",
         17272 => x"00000000",
         17273 => x"00000000",
         17274 => x"00000000",
         17275 => x"00000000",
         17276 => x"00000000",
         17277 => x"00000000",
         17278 => x"00000000",
         17279 => x"00000000",
         17280 => x"00000000",
         17281 => x"00000000",
         17282 => x"00000000",
         17283 => x"00000000",
         17284 => x"00000000",
         17285 => x"00000000",
         17286 => x"00000000",
         17287 => x"00000000",
         17288 => x"00000000",
         17289 => x"00000000",
         17290 => x"00000000",
         17291 => x"00000000",
         17292 => x"00000000",
         17293 => x"00000000",
         17294 => x"00000000",
         17295 => x"00000000",
         17296 => x"00000000",
         17297 => x"00000000",
         17298 => x"00000000",
         17299 => x"00000000",
         17300 => x"00000000",
         17301 => x"00000000",
         17302 => x"00000000",
         17303 => x"00000000",
         17304 => x"00000000",
         17305 => x"00000000",
         17306 => x"00000000",
         17307 => x"00000000",
         17308 => x"00000000",
         17309 => x"00000000",
         17310 => x"00000000",
         17311 => x"00000000",
         17312 => x"00000000",
         17313 => x"00000000",
         17314 => x"00000000",
         17315 => x"00000000",
         17316 => x"00000000",
         17317 => x"00000000",
         17318 => x"00000000",
         17319 => x"00000000",
         17320 => x"00000000",
         17321 => x"00000000",
         17322 => x"00000000",
         17323 => x"00000000",
         17324 => x"00000000",
         17325 => x"00000000",
         17326 => x"00000000",
         17327 => x"00000000",
         17328 => x"00000000",
         17329 => x"00000000",
         17330 => x"00000000",
         17331 => x"00000000",
         17332 => x"00000000",
         17333 => x"00000000",
         17334 => x"00000000",
         17335 => x"00000000",
         17336 => x"00000000",
         17337 => x"00000000",
         17338 => x"00000000",
         17339 => x"00000000",
         17340 => x"00000000",
         17341 => x"00000000",
         17342 => x"00000000",
         17343 => x"00000000",
         17344 => x"00000000",
         17345 => x"00000000",
         17346 => x"00000000",
         17347 => x"00000000",
         17348 => x"00000000",
         17349 => x"00000000",
         17350 => x"00000000",
         17351 => x"00000000",
         17352 => x"00000000",
         17353 => x"00000000",
         17354 => x"00000000",
         17355 => x"00000000",
         17356 => x"00000000",
         17357 => x"00000000",
         17358 => x"00000000",
         17359 => x"00000000",
         17360 => x"00000000",
         17361 => x"00000000",
         17362 => x"00000000",
         17363 => x"00000000",
         17364 => x"00000000",
         17365 => x"00000000",
         17366 => x"00000000",
         17367 => x"00000000",
         17368 => x"00000000",
         17369 => x"00000000",
         17370 => x"00000000",
         17371 => x"00000000",
         17372 => x"00000000",
         17373 => x"00000000",
         17374 => x"00000000",
         17375 => x"00000000",
         17376 => x"00000000",
         17377 => x"00000000",
         17378 => x"00000000",
         17379 => x"00000000",
         17380 => x"00000000",
         17381 => x"00000000",
         17382 => x"00000000",
         17383 => x"00000000",
         17384 => x"00000000",
         17385 => x"00000000",
         17386 => x"00000000",
         17387 => x"00000000",
         17388 => x"00000000",
         17389 => x"00000000",
         17390 => x"00000000",
         17391 => x"00000000",
         17392 => x"00000000",
         17393 => x"00000000",
         17394 => x"00000000",
         17395 => x"00000000",
         17396 => x"00000000",
         17397 => x"00000000",
         17398 => x"00000000",
         17399 => x"00000000",
         17400 => x"00000000",
         17401 => x"00000000",
         17402 => x"00000000",
         17403 => x"00000000",
         17404 => x"00000000",
         17405 => x"00000000",
         17406 => x"00000000",
         17407 => x"00000000",
         17408 => x"00000000",
         17409 => x"00000000",
         17410 => x"00000000",
         17411 => x"00000000",
         17412 => x"00000000",
         17413 => x"00000000",
         17414 => x"00000000",
         17415 => x"00000000",
         17416 => x"00000000",
         17417 => x"00000000",
         17418 => x"00000000",
         17419 => x"00000000",
         17420 => x"00000000",
         17421 => x"00000000",
         17422 => x"00000000",
         17423 => x"00000000",
         17424 => x"00000000",
         17425 => x"00000000",
         17426 => x"00000000",
         17427 => x"00000000",
         17428 => x"00000000",
         17429 => x"00000000",
         17430 => x"00000000",
         17431 => x"00000000",
         17432 => x"00000000",
         17433 => x"00000000",
         17434 => x"00000000",
         17435 => x"00000000",
         17436 => x"00000000",
         17437 => x"00000000",
         17438 => x"00000000",
         17439 => x"00000000",
         17440 => x"00000000",
         17441 => x"00000000",
         17442 => x"00000000",
         17443 => x"00000000",
         17444 => x"00000000",
         17445 => x"00000000",
         17446 => x"00000000",
         17447 => x"00000000",
         17448 => x"00000000",
         17449 => x"00000000",
         17450 => x"00000000",
         17451 => x"00000000",
         17452 => x"00000000",
         17453 => x"00000000",
         17454 => x"00000000",
         17455 => x"00000000",
         17456 => x"00000000",
         17457 => x"00000000",
         17458 => x"00000000",
         17459 => x"00000000",
         17460 => x"00000000",
         17461 => x"00000000",
         17462 => x"00000000",
         17463 => x"00000000",
         17464 => x"00000000",
         17465 => x"00000000",
         17466 => x"00000000",
         17467 => x"00000000",
         17468 => x"00000000",
         17469 => x"00000000",
         17470 => x"00000000",
         17471 => x"00000000",
         17472 => x"00000000",
         17473 => x"00000000",
         17474 => x"00000000",
         17475 => x"00000000",
         17476 => x"00000000",
         17477 => x"00000000",
         17478 => x"00000000",
         17479 => x"00000000",
         17480 => x"00000000",
         17481 => x"00000000",
         17482 => x"00000000",
         17483 => x"00000000",
         17484 => x"00000000",
         17485 => x"00000000",
         17486 => x"00000000",
         17487 => x"00000000",
         17488 => x"00000000",
         17489 => x"00000000",
         17490 => x"00000000",
         17491 => x"00000000",
         17492 => x"00000000",
         17493 => x"00000000",
         17494 => x"00000000",
         17495 => x"00000000",
         17496 => x"00000000",
         17497 => x"00000000",
         17498 => x"00000000",
         17499 => x"00000000",
         17500 => x"00000000",
         17501 => x"00000000",
         17502 => x"00000000",
         17503 => x"00000000",
         17504 => x"00000000",
         17505 => x"00000000",
         17506 => x"00000000",
         17507 => x"00000000",
         17508 => x"00000000",
         17509 => x"00000000",
         17510 => x"00000000",
         17511 => x"00000000",
         17512 => x"00000000",
         17513 => x"00000000",
         17514 => x"00000000",
         17515 => x"00000000",
         17516 => x"00000000",
         17517 => x"00000000",
         17518 => x"00000000",
         17519 => x"00000000",
         17520 => x"00000000",
         17521 => x"00000000",
         17522 => x"00000000",
         17523 => x"00000000",
         17524 => x"00000000",
         17525 => x"00000000",
         17526 => x"00000000",
         17527 => x"00000000",
         17528 => x"00000000",
         17529 => x"00000000",
         17530 => x"00000000",
         17531 => x"00000000",
         17532 => x"00000000",
         17533 => x"00000000",
         17534 => x"00000000",
         17535 => x"00000000",
         17536 => x"00000000",
         17537 => x"00000000",
         17538 => x"00000000",
         17539 => x"00000000",
         17540 => x"00000000",
         17541 => x"00000000",
         17542 => x"00000000",
         17543 => x"00000000",
         17544 => x"00000000",
         17545 => x"00000000",
         17546 => x"00000000",
         17547 => x"00000000",
         17548 => x"00000000",
         17549 => x"00000000",
         17550 => x"00000000",
         17551 => x"00000000",
         17552 => x"00000000",
         17553 => x"00000000",
         17554 => x"00000000",
         17555 => x"00000000",
         17556 => x"00000000",
         17557 => x"00000000",
         17558 => x"00000000",
         17559 => x"00000000",
         17560 => x"00000000",
         17561 => x"00000000",
         17562 => x"00000000",
         17563 => x"00000000",
         17564 => x"00000000",
         17565 => x"00000000",
         17566 => x"00000000",
         17567 => x"00000000",
         17568 => x"00000000",
         17569 => x"00000000",
         17570 => x"00000000",
         17571 => x"00000000",
         17572 => x"00000000",
         17573 => x"00000000",
         17574 => x"00000000",
         17575 => x"00000000",
         17576 => x"00000000",
         17577 => x"00000000",
         17578 => x"00000000",
         17579 => x"00000000",
         17580 => x"00000000",
         17581 => x"00000000",
         17582 => x"00000000",
         17583 => x"00000000",
         17584 => x"00000000",
         17585 => x"00000000",
         17586 => x"00000000",
         17587 => x"00000000",
         17588 => x"00000000",
         17589 => x"00000000",
         17590 => x"00000000",
         17591 => x"00000000",
         17592 => x"00000000",
         17593 => x"00000000",
         17594 => x"00000000",
         17595 => x"00000000",
         17596 => x"00000000",
         17597 => x"00000000",
         17598 => x"00000000",
         17599 => x"00000000",
         17600 => x"00000000",
         17601 => x"00000000",
         17602 => x"00000000",
         17603 => x"00000000",
         17604 => x"00000000",
         17605 => x"00000000",
         17606 => x"00000000",
         17607 => x"00000000",
         17608 => x"00000000",
         17609 => x"00000000",
         17610 => x"00000000",
         17611 => x"00000000",
         17612 => x"00000000",
         17613 => x"00000000",
         17614 => x"00000000",
         17615 => x"00000000",
         17616 => x"00000000",
         17617 => x"00000000",
         17618 => x"00000000",
         17619 => x"00000000",
         17620 => x"00000000",
         17621 => x"00000000",
         17622 => x"00000000",
         17623 => x"00000000",
         17624 => x"00000000",
         17625 => x"00000000",
         17626 => x"00000000",
         17627 => x"00000000",
         17628 => x"00000000",
         17629 => x"00000000",
         17630 => x"00000000",
         17631 => x"00000000",
         17632 => x"00000000",
         17633 => x"00000000",
         17634 => x"00000000",
         17635 => x"00000000",
         17636 => x"00000000",
         17637 => x"00000000",
         17638 => x"00000000",
         17639 => x"00000000",
         17640 => x"00000000",
         17641 => x"00000000",
         17642 => x"00000000",
         17643 => x"00000000",
         17644 => x"00000000",
         17645 => x"00000000",
         17646 => x"00000000",
         17647 => x"00000000",
         17648 => x"00000000",
         17649 => x"00000000",
         17650 => x"00000000",
         17651 => x"00000000",
         17652 => x"00000000",
         17653 => x"00000000",
         17654 => x"00000000",
         17655 => x"00000000",
         17656 => x"00000000",
         17657 => x"00000000",
         17658 => x"00000000",
         17659 => x"00000000",
         17660 => x"00000000",
         17661 => x"00000000",
         17662 => x"00000000",
         17663 => x"00000000",
         17664 => x"00000000",
         17665 => x"00000000",
         17666 => x"00000000",
         17667 => x"00000000",
         17668 => x"00000000",
         17669 => x"00000000",
         17670 => x"00000000",
         17671 => x"00000000",
         17672 => x"00000000",
         17673 => x"00000000",
         17674 => x"00000000",
         17675 => x"00000000",
         17676 => x"00000000",
         17677 => x"00000000",
         17678 => x"00000000",
         17679 => x"00000000",
         17680 => x"00000000",
         17681 => x"00000000",
         17682 => x"00000000",
         17683 => x"00000000",
         17684 => x"00000000",
         17685 => x"00000000",
         17686 => x"00000000",
         17687 => x"00000000",
         17688 => x"00000000",
         17689 => x"00000000",
         17690 => x"00000000",
         17691 => x"00000000",
         17692 => x"00000000",
         17693 => x"00000000",
         17694 => x"00000000",
         17695 => x"00000000",
         17696 => x"00000000",
         17697 => x"00000000",
         17698 => x"00000000",
         17699 => x"00000000",
         17700 => x"00000000",
         17701 => x"00000000",
         17702 => x"00000000",
         17703 => x"00000000",
         17704 => x"00000000",
         17705 => x"00000000",
         17706 => x"00000000",
         17707 => x"00000000",
         17708 => x"00000000",
         17709 => x"00000000",
         17710 => x"00000000",
         17711 => x"00000000",
         17712 => x"00000000",
         17713 => x"00000000",
         17714 => x"00000000",
         17715 => x"00000000",
         17716 => x"00000000",
         17717 => x"00000000",
         17718 => x"00000000",
         17719 => x"00000000",
         17720 => x"00000000",
         17721 => x"00000000",
         17722 => x"00000000",
         17723 => x"00000000",
         17724 => x"00000000",
         17725 => x"00000000",
         17726 => x"00000000",
         17727 => x"00000000",
         17728 => x"00000000",
         17729 => x"00000000",
         17730 => x"00000000",
         17731 => x"00000000",
         17732 => x"00000000",
         17733 => x"00000000",
         17734 => x"00000000",
         17735 => x"00000000",
         17736 => x"00000000",
         17737 => x"00000000",
         17738 => x"00000000",
         17739 => x"00000000",
         17740 => x"00000000",
         17741 => x"00000000",
         17742 => x"00000000",
         17743 => x"00000000",
         17744 => x"00000000",
         17745 => x"00000000",
         17746 => x"00000000",
         17747 => x"00000000",
         17748 => x"00000000",
         17749 => x"00000000",
         17750 => x"00000000",
         17751 => x"00000000",
         17752 => x"00000000",
         17753 => x"00000000",
         17754 => x"00000000",
         17755 => x"00000000",
         17756 => x"00000000",
         17757 => x"00000000",
         17758 => x"00000000",
         17759 => x"00000000",
         17760 => x"00000000",
         17761 => x"00000000",
         17762 => x"00000000",
         17763 => x"00000000",
         17764 => x"00000000",
         17765 => x"00000000",
         17766 => x"00000000",
         17767 => x"00000000",
         17768 => x"00000000",
         17769 => x"00000000",
         17770 => x"00000000",
         17771 => x"00000000",
         17772 => x"00000000",
         17773 => x"00000000",
         17774 => x"00000000",
         17775 => x"00000000",
         17776 => x"00000000",
         17777 => x"00000000",
         17778 => x"00000000",
         17779 => x"00000000",
         17780 => x"00000000",
         17781 => x"00000000",
         17782 => x"00000000",
         17783 => x"00000000",
         17784 => x"00000000",
         17785 => x"00000000",
         17786 => x"00000000",
         17787 => x"00000000",
         17788 => x"00000000",
         17789 => x"00000000",
         17790 => x"00000000",
         17791 => x"00000000",
         17792 => x"00000000",
         17793 => x"00000000",
         17794 => x"00000000",
         17795 => x"00000000",
         17796 => x"00000000",
         17797 => x"00000000",
         17798 => x"00000000",
         17799 => x"00000000",
         17800 => x"00000000",
         17801 => x"00000000",
         17802 => x"00000000",
         17803 => x"00000000",
         17804 => x"00000000",
         17805 => x"00000000",
         17806 => x"00000000",
         17807 => x"00000000",
         17808 => x"00000000",
         17809 => x"00000000",
         17810 => x"00000000",
         17811 => x"00000000",
         17812 => x"00000000",
         17813 => x"00000000",
         17814 => x"00000000",
         17815 => x"00000000",
         17816 => x"00000000",
         17817 => x"00000000",
         17818 => x"00000000",
         17819 => x"00000000",
         17820 => x"00000000",
         17821 => x"00000000",
         17822 => x"00000000",
         17823 => x"00000000",
         17824 => x"00000000",
         17825 => x"00000000",
         17826 => x"00000000",
         17827 => x"00000000",
         17828 => x"00000000",
         17829 => x"00000000",
         17830 => x"00000000",
         17831 => x"00000000",
         17832 => x"00000000",
         17833 => x"00000000",
         17834 => x"00000000",
         17835 => x"00000000",
         17836 => x"00000000",
         17837 => x"00000000",
         17838 => x"00000000",
         17839 => x"00000000",
         17840 => x"00000000",
         17841 => x"00000000",
         17842 => x"00000000",
         17843 => x"00000000",
         17844 => x"00000000",
         17845 => x"00000000",
         17846 => x"00000000",
         17847 => x"00000000",
         17848 => x"00000000",
         17849 => x"00000000",
         17850 => x"00000000",
         17851 => x"00000000",
         17852 => x"00000000",
         17853 => x"00000000",
         17854 => x"00000000",
         17855 => x"00000000",
         17856 => x"00000000",
         17857 => x"00000000",
         17858 => x"00000000",
         17859 => x"00000000",
         17860 => x"00000000",
         17861 => x"00000000",
         17862 => x"00000000",
         17863 => x"00000000",
         17864 => x"00000000",
         17865 => x"00000000",
         17866 => x"00000000",
         17867 => x"00000000",
         17868 => x"00000000",
         17869 => x"00000000",
         17870 => x"00000000",
         17871 => x"00000000",
         17872 => x"00000000",
         17873 => x"00000000",
         17874 => x"00000000",
         17875 => x"00000000",
         17876 => x"00000000",
         17877 => x"00000000",
         17878 => x"00000000",
         17879 => x"00000000",
         17880 => x"00000000",
         17881 => x"00000000",
         17882 => x"00000000",
         17883 => x"00000000",
         17884 => x"00000000",
         17885 => x"00000000",
         17886 => x"00000000",
         17887 => x"00000000",
         17888 => x"00000000",
         17889 => x"00000000",
         17890 => x"00000000",
         17891 => x"00000000",
         17892 => x"00000000",
         17893 => x"00000000",
         17894 => x"00000000",
         17895 => x"00000000",
         17896 => x"00000000",
         17897 => x"00000000",
         17898 => x"00000000",
         17899 => x"00000000",
         17900 => x"00000000",
         17901 => x"00000000",
         17902 => x"00000000",
         17903 => x"00000000",
         17904 => x"00000000",
         17905 => x"00000000",
         17906 => x"00000000",
         17907 => x"00000000",
         17908 => x"00000000",
         17909 => x"00000000",
         17910 => x"00000000",
         17911 => x"00000000",
         17912 => x"00000000",
         17913 => x"00000000",
         17914 => x"00000000",
         17915 => x"00000000",
         17916 => x"00000000",
         17917 => x"00000000",
         17918 => x"00000000",
         17919 => x"00000000",
         17920 => x"00000000",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"00000000",
         17924 => x"00000000",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"00000000",
         17928 => x"00000000",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"00000000",
         17932 => x"00000000",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"00000000",
         17936 => x"00000000",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"00000000",
         17940 => x"00000000",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"00000000",
         17944 => x"00000000",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"00000000",
         17948 => x"00000000",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"00000000",
         17952 => x"00000000",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"00000000",
         17956 => x"00000000",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"00000000",
         17962 => x"00000000",
         17963 => x"00000000",
         17964 => x"00000000",
         17965 => x"00000000",
         17966 => x"00000000",
         17967 => x"00000000",
         17968 => x"00000000",
         17969 => x"00000000",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"00000000",
         17973 => x"00000000",
         17974 => x"00000000",
         17975 => x"00000000",
         17976 => x"00000000",
         17977 => x"00000000",
         17978 => x"00000000",
         17979 => x"00000000",
         17980 => x"00000000",
         17981 => x"00000000",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00000000",
         18004 => x"00000000",
         18005 => x"00000000",
         18006 => x"00000000",
         18007 => x"00000000",
         18008 => x"00000000",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"00000000",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"00000000",
         18016 => x"00000000",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"00000000",
         18020 => x"00000000",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"00000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00000000",
         18034 => x"00000000",
         18035 => x"00000000",
         18036 => x"00000000",
         18037 => x"00000000",
         18038 => x"00000000",
         18039 => x"00000000",
         18040 => x"00000000",
         18041 => x"00000000",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00000000",
         18045 => x"00000000",
         18046 => x"00000000",
         18047 => x"00000000",
         18048 => x"00000000",
         18049 => x"00000000",
         18050 => x"00000000",
         18051 => x"00000000",
         18052 => x"00000000",
         18053 => x"00000000",
         18054 => x"00000000",
         18055 => x"00000000",
         18056 => x"00000000",
         18057 => x"00000000",
         18058 => x"00000000",
         18059 => x"00000000",
         18060 => x"00000000",
         18061 => x"00000000",
         18062 => x"00000000",
         18063 => x"00000000",
         18064 => x"00000000",
         18065 => x"00000000",
         18066 => x"00000000",
         18067 => x"00000000",
         18068 => x"00000000",
         18069 => x"00000000",
         18070 => x"00000000",
         18071 => x"00000000",
         18072 => x"00000000",
         18073 => x"00000000",
         18074 => x"00000000",
         18075 => x"00000000",
         18076 => x"00000000",
         18077 => x"00000000",
         18078 => x"00000000",
         18079 => x"00000000",
         18080 => x"00000000",
         18081 => x"00000000",
         18082 => x"00000000",
         18083 => x"00000000",
         18084 => x"00000000",
         18085 => x"00000000",
         18086 => x"00000000",
         18087 => x"00000000",
         18088 => x"00000000",
         18089 => x"00000000",
         18090 => x"00000000",
         18091 => x"00000000",
         18092 => x"00000000",
         18093 => x"00000000",
         18094 => x"00000000",
         18095 => x"00000000",
         18096 => x"00000000",
         18097 => x"00000000",
         18098 => x"00000000",
         18099 => x"00000000",
         18100 => x"00000000",
         18101 => x"00000000",
         18102 => x"00000000",
         18103 => x"00000000",
         18104 => x"00000000",
         18105 => x"00000000",
         18106 => x"00000000",
         18107 => x"00000000",
         18108 => x"00000000",
         18109 => x"00000000",
         18110 => x"00000000",
         18111 => x"00000000",
         18112 => x"00000000",
         18113 => x"00000000",
         18114 => x"00000000",
         18115 => x"00000000",
         18116 => x"00000000",
         18117 => x"00000000",
         18118 => x"00000000",
         18119 => x"00000000",
         18120 => x"00000000",
         18121 => x"00000000",
         18122 => x"00000000",
         18123 => x"00000000",
         18124 => x"00000000",
         18125 => x"00000000",
         18126 => x"00000000",
         18127 => x"00000000",
         18128 => x"00000000",
         18129 => x"00000000",
         18130 => x"00000000",
         18131 => x"00000000",
         18132 => x"00000000",
         18133 => x"00003219",
         18134 => x"50000100",
         18135 => x"00000000",
         18136 => x"cce0f2f3",
         18137 => x"cecff6f7",
         18138 => x"f8f9fafb",
         18139 => x"fcfdfeff",
         18140 => x"e1c1c2c3",
         18141 => x"c4c5c6e2",
         18142 => x"e3e4e5e6",
         18143 => x"ebeeeff4",
         18144 => x"00616263",
         18145 => x"64656667",
         18146 => x"68696b6a",
         18147 => x"2f2a2e2d",
         18148 => x"20212223",
         18149 => x"24252627",
         18150 => x"28294f2c",
         18151 => x"512b5749",
         18152 => x"55010203",
         18153 => x"04050607",
         18154 => x"08090a0b",
         18155 => x"0c0d0e0f",
         18156 => x"10111213",
         18157 => x"14151617",
         18158 => x"18191a52",
         18159 => x"5954be3c",
         18160 => x"c7818283",
         18161 => x"84858687",
         18162 => x"88898a8b",
         18163 => x"8c8d8e8f",
         18164 => x"90919293",
         18165 => x"94959697",
         18166 => x"98999abc",
         18167 => x"8040a5c0",
         18168 => x"00000000",
         18169 => x"00000000",
         18170 => x"00000000",
         18171 => x"00000000",
         18172 => x"00000000",
         18173 => x"00000000",
         18174 => x"00000000",
         18175 => x"00000000",
         18176 => x"00000000",
         18177 => x"00000000",
         18178 => x"00000000",
         18179 => x"00000000",
         18180 => x"00000000",
         18181 => x"00000000",
         18182 => x"00000000",
         18183 => x"00000000",
         18184 => x"00000000",
         18185 => x"00000000",
         18186 => x"00000000",
         18187 => x"00000000",
         18188 => x"00000000",
         18189 => x"00000000",
         18190 => x"00000000",
         18191 => x"00000000",
         18192 => x"00000000",
         18193 => x"00000000",
         18194 => x"00000000",
         18195 => x"00000000",
         18196 => x"00000000",
         18197 => x"00000000",
         18198 => x"00020003",
         18199 => x"00040101",
         18200 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

