-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"fe",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"94",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"cf",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"d1",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"b4",
           386 => x"c6",
           387 => x"b4",
           388 => x"90",
           389 => x"b4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"82",
           396 => x"82",
           397 => x"b4",
           398 => x"b5",
           399 => x"d0",
           400 => x"b5",
           401 => x"ab",
           402 => x"b4",
           403 => x"90",
           404 => x"b4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"82",
           410 => x"82",
           411 => x"82",
           412 => x"af",
           413 => x"b5",
           414 => x"d0",
           415 => x"b5",
           416 => x"d6",
           417 => x"b4",
           418 => x"90",
           419 => x"b4",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"82",
           425 => x"82",
           426 => x"82",
           427 => x"80",
           428 => x"82",
           429 => x"82",
           430 => x"82",
           431 => x"80",
           432 => x"82",
           433 => x"82",
           434 => x"82",
           435 => x"80",
           436 => x"82",
           437 => x"82",
           438 => x"82",
           439 => x"80",
           440 => x"82",
           441 => x"82",
           442 => x"82",
           443 => x"80",
           444 => x"82",
           445 => x"82",
           446 => x"82",
           447 => x"81",
           448 => x"82",
           449 => x"82",
           450 => x"82",
           451 => x"81",
           452 => x"82",
           453 => x"82",
           454 => x"82",
           455 => x"81",
           456 => x"82",
           457 => x"82",
           458 => x"82",
           459 => x"81",
           460 => x"82",
           461 => x"82",
           462 => x"82",
           463 => x"81",
           464 => x"82",
           465 => x"82",
           466 => x"82",
           467 => x"81",
           468 => x"82",
           469 => x"82",
           470 => x"82",
           471 => x"81",
           472 => x"82",
           473 => x"82",
           474 => x"82",
           475 => x"81",
           476 => x"82",
           477 => x"82",
           478 => x"82",
           479 => x"81",
           480 => x"82",
           481 => x"82",
           482 => x"82",
           483 => x"81",
           484 => x"82",
           485 => x"82",
           486 => x"82",
           487 => x"81",
           488 => x"82",
           489 => x"82",
           490 => x"82",
           491 => x"81",
           492 => x"82",
           493 => x"82",
           494 => x"82",
           495 => x"81",
           496 => x"82",
           497 => x"82",
           498 => x"82",
           499 => x"81",
           500 => x"82",
           501 => x"82",
           502 => x"82",
           503 => x"81",
           504 => x"82",
           505 => x"82",
           506 => x"82",
           507 => x"81",
           508 => x"82",
           509 => x"82",
           510 => x"82",
           511 => x"81",
           512 => x"82",
           513 => x"82",
           514 => x"82",
           515 => x"81",
           516 => x"82",
           517 => x"82",
           518 => x"82",
           519 => x"81",
           520 => x"82",
           521 => x"82",
           522 => x"82",
           523 => x"81",
           524 => x"82",
           525 => x"82",
           526 => x"82",
           527 => x"81",
           528 => x"82",
           529 => x"82",
           530 => x"82",
           531 => x"81",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"81",
           540 => x"82",
           541 => x"82",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"82",
           555 => x"81",
           556 => x"82",
           557 => x"82",
           558 => x"82",
           559 => x"81",
           560 => x"82",
           561 => x"82",
           562 => x"82",
           563 => x"81",
           564 => x"82",
           565 => x"82",
           566 => x"82",
           567 => x"80",
           568 => x"82",
           569 => x"82",
           570 => x"82",
           571 => x"80",
           572 => x"82",
           573 => x"82",
           574 => x"82",
           575 => x"80",
           576 => x"82",
           577 => x"82",
           578 => x"82",
           579 => x"80",
           580 => x"82",
           581 => x"82",
           582 => x"82",
           583 => x"81",
           584 => x"82",
           585 => x"82",
           586 => x"82",
           587 => x"81",
           588 => x"82",
           589 => x"82",
           590 => x"82",
           591 => x"81",
           592 => x"82",
           593 => x"82",
           594 => x"82",
           595 => x"81",
           596 => x"82",
           597 => x"82",
           598 => x"3c",
           599 => x"10",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"51",
           608 => x"73",
           609 => x"73",
           610 => x"81",
           611 => x"10",
           612 => x"07",
           613 => x"0c",
           614 => x"72",
           615 => x"81",
           616 => x"09",
           617 => x"71",
           618 => x"0a",
           619 => x"72",
           620 => x"51",
           621 => x"82",
           622 => x"82",
           623 => x"8e",
           624 => x"70",
           625 => x"0c",
           626 => x"93",
           627 => x"81",
           628 => x"cb",
           629 => x"b5",
           630 => x"82",
           631 => x"fb",
           632 => x"b5",
           633 => x"05",
           634 => x"b4",
           635 => x"0c",
           636 => x"08",
           637 => x"54",
           638 => x"08",
           639 => x"53",
           640 => x"08",
           641 => x"9a",
           642 => x"a8",
           643 => x"b5",
           644 => x"05",
           645 => x"b4",
           646 => x"08",
           647 => x"a8",
           648 => x"87",
           649 => x"b5",
           650 => x"82",
           651 => x"02",
           652 => x"0c",
           653 => x"82",
           654 => x"90",
           655 => x"11",
           656 => x"32",
           657 => x"51",
           658 => x"71",
           659 => x"0b",
           660 => x"08",
           661 => x"25",
           662 => x"39",
           663 => x"b5",
           664 => x"05",
           665 => x"39",
           666 => x"08",
           667 => x"ff",
           668 => x"b4",
           669 => x"0c",
           670 => x"b5",
           671 => x"05",
           672 => x"b4",
           673 => x"08",
           674 => x"08",
           675 => x"82",
           676 => x"f8",
           677 => x"2e",
           678 => x"80",
           679 => x"b4",
           680 => x"08",
           681 => x"38",
           682 => x"08",
           683 => x"51",
           684 => x"82",
           685 => x"70",
           686 => x"08",
           687 => x"52",
           688 => x"08",
           689 => x"ff",
           690 => x"06",
           691 => x"0b",
           692 => x"08",
           693 => x"80",
           694 => x"b5",
           695 => x"05",
           696 => x"b4",
           697 => x"08",
           698 => x"73",
           699 => x"b4",
           700 => x"08",
           701 => x"b5",
           702 => x"05",
           703 => x"b4",
           704 => x"08",
           705 => x"b5",
           706 => x"05",
           707 => x"39",
           708 => x"08",
           709 => x"52",
           710 => x"82",
           711 => x"88",
           712 => x"82",
           713 => x"f4",
           714 => x"82",
           715 => x"f4",
           716 => x"b5",
           717 => x"3d",
           718 => x"b4",
           719 => x"b5",
           720 => x"82",
           721 => x"f4",
           722 => x"0b",
           723 => x"08",
           724 => x"82",
           725 => x"88",
           726 => x"b5",
           727 => x"05",
           728 => x"0b",
           729 => x"08",
           730 => x"82",
           731 => x"90",
           732 => x"b5",
           733 => x"05",
           734 => x"b4",
           735 => x"08",
           736 => x"b4",
           737 => x"08",
           738 => x"b4",
           739 => x"70",
           740 => x"81",
           741 => x"b5",
           742 => x"82",
           743 => x"dc",
           744 => x"b5",
           745 => x"05",
           746 => x"b4",
           747 => x"08",
           748 => x"80",
           749 => x"b5",
           750 => x"05",
           751 => x"b5",
           752 => x"8e",
           753 => x"b5",
           754 => x"82",
           755 => x"02",
           756 => x"0c",
           757 => x"82",
           758 => x"90",
           759 => x"b5",
           760 => x"05",
           761 => x"b4",
           762 => x"08",
           763 => x"b4",
           764 => x"08",
           765 => x"b4",
           766 => x"08",
           767 => x"3f",
           768 => x"08",
           769 => x"b4",
           770 => x"0c",
           771 => x"08",
           772 => x"70",
           773 => x"0c",
           774 => x"3d",
           775 => x"b4",
           776 => x"b5",
           777 => x"82",
           778 => x"ed",
           779 => x"0b",
           780 => x"08",
           781 => x"82",
           782 => x"88",
           783 => x"80",
           784 => x"0c",
           785 => x"08",
           786 => x"85",
           787 => x"81",
           788 => x"32",
           789 => x"51",
           790 => x"53",
           791 => x"8d",
           792 => x"82",
           793 => x"e0",
           794 => x"ac",
           795 => x"b4",
           796 => x"08",
           797 => x"53",
           798 => x"b4",
           799 => x"34",
           800 => x"06",
           801 => x"2e",
           802 => x"82",
           803 => x"8c",
           804 => x"05",
           805 => x"08",
           806 => x"82",
           807 => x"e4",
           808 => x"81",
           809 => x"72",
           810 => x"8b",
           811 => x"b4",
           812 => x"33",
           813 => x"27",
           814 => x"82",
           815 => x"f8",
           816 => x"72",
           817 => x"ee",
           818 => x"b4",
           819 => x"33",
           820 => x"2e",
           821 => x"80",
           822 => x"b5",
           823 => x"05",
           824 => x"2b",
           825 => x"51",
           826 => x"b2",
           827 => x"b4",
           828 => x"22",
           829 => x"70",
           830 => x"81",
           831 => x"51",
           832 => x"2e",
           833 => x"b5",
           834 => x"05",
           835 => x"80",
           836 => x"72",
           837 => x"08",
           838 => x"fe",
           839 => x"b5",
           840 => x"05",
           841 => x"2b",
           842 => x"70",
           843 => x"72",
           844 => x"51",
           845 => x"51",
           846 => x"82",
           847 => x"e8",
           848 => x"b5",
           849 => x"05",
           850 => x"b5",
           851 => x"05",
           852 => x"d0",
           853 => x"53",
           854 => x"b4",
           855 => x"34",
           856 => x"08",
           857 => x"70",
           858 => x"98",
           859 => x"53",
           860 => x"8b",
           861 => x"0b",
           862 => x"08",
           863 => x"82",
           864 => x"e4",
           865 => x"83",
           866 => x"06",
           867 => x"72",
           868 => x"82",
           869 => x"e8",
           870 => x"88",
           871 => x"2b",
           872 => x"70",
           873 => x"51",
           874 => x"72",
           875 => x"08",
           876 => x"fd",
           877 => x"b5",
           878 => x"05",
           879 => x"2a",
           880 => x"51",
           881 => x"80",
           882 => x"82",
           883 => x"e8",
           884 => x"98",
           885 => x"2c",
           886 => x"72",
           887 => x"0b",
           888 => x"08",
           889 => x"82",
           890 => x"f8",
           891 => x"11",
           892 => x"08",
           893 => x"53",
           894 => x"08",
           895 => x"80",
           896 => x"94",
           897 => x"b4",
           898 => x"08",
           899 => x"82",
           900 => x"70",
           901 => x"51",
           902 => x"82",
           903 => x"e4",
           904 => x"90",
           905 => x"72",
           906 => x"08",
           907 => x"82",
           908 => x"e4",
           909 => x"a0",
           910 => x"72",
           911 => x"08",
           912 => x"fc",
           913 => x"b5",
           914 => x"05",
           915 => x"80",
           916 => x"72",
           917 => x"08",
           918 => x"fc",
           919 => x"b5",
           920 => x"05",
           921 => x"c0",
           922 => x"72",
           923 => x"08",
           924 => x"fb",
           925 => x"b5",
           926 => x"05",
           927 => x"07",
           928 => x"82",
           929 => x"e4",
           930 => x"0b",
           931 => x"08",
           932 => x"fb",
           933 => x"b5",
           934 => x"05",
           935 => x"07",
           936 => x"82",
           937 => x"e4",
           938 => x"c1",
           939 => x"82",
           940 => x"fc",
           941 => x"b5",
           942 => x"05",
           943 => x"51",
           944 => x"b5",
           945 => x"05",
           946 => x"0b",
           947 => x"08",
           948 => x"8d",
           949 => x"b5",
           950 => x"05",
           951 => x"b4",
           952 => x"08",
           953 => x"b5",
           954 => x"05",
           955 => x"51",
           956 => x"b5",
           957 => x"05",
           958 => x"b4",
           959 => x"22",
           960 => x"53",
           961 => x"b4",
           962 => x"23",
           963 => x"82",
           964 => x"90",
           965 => x"b5",
           966 => x"05",
           967 => x"82",
           968 => x"90",
           969 => x"08",
           970 => x"08",
           971 => x"82",
           972 => x"e4",
           973 => x"83",
           974 => x"06",
           975 => x"53",
           976 => x"ab",
           977 => x"b4",
           978 => x"33",
           979 => x"53",
           980 => x"53",
           981 => x"08",
           982 => x"52",
           983 => x"3f",
           984 => x"08",
           985 => x"b5",
           986 => x"05",
           987 => x"82",
           988 => x"fc",
           989 => x"a8",
           990 => x"b5",
           991 => x"72",
           992 => x"08",
           993 => x"82",
           994 => x"ec",
           995 => x"82",
           996 => x"f4",
           997 => x"71",
           998 => x"72",
           999 => x"08",
          1000 => x"8b",
          1001 => x"b5",
          1002 => x"05",
          1003 => x"b4",
          1004 => x"08",
          1005 => x"b5",
          1006 => x"05",
          1007 => x"82",
          1008 => x"fc",
          1009 => x"b5",
          1010 => x"05",
          1011 => x"2a",
          1012 => x"51",
          1013 => x"72",
          1014 => x"38",
          1015 => x"08",
          1016 => x"70",
          1017 => x"72",
          1018 => x"82",
          1019 => x"fc",
          1020 => x"53",
          1021 => x"82",
          1022 => x"53",
          1023 => x"b4",
          1024 => x"23",
          1025 => x"b5",
          1026 => x"05",
          1027 => x"95",
          1028 => x"a8",
          1029 => x"82",
          1030 => x"f4",
          1031 => x"b5",
          1032 => x"05",
          1033 => x"b5",
          1034 => x"05",
          1035 => x"31",
          1036 => x"82",
          1037 => x"ec",
          1038 => x"c1",
          1039 => x"b4",
          1040 => x"22",
          1041 => x"70",
          1042 => x"51",
          1043 => x"2e",
          1044 => x"b5",
          1045 => x"05",
          1046 => x"b4",
          1047 => x"08",
          1048 => x"b5",
          1049 => x"05",
          1050 => x"82",
          1051 => x"dc",
          1052 => x"a2",
          1053 => x"b4",
          1054 => x"08",
          1055 => x"08",
          1056 => x"84",
          1057 => x"b4",
          1058 => x"0c",
          1059 => x"b5",
          1060 => x"05",
          1061 => x"b5",
          1062 => x"05",
          1063 => x"b4",
          1064 => x"0c",
          1065 => x"08",
          1066 => x"80",
          1067 => x"82",
          1068 => x"e4",
          1069 => x"82",
          1070 => x"72",
          1071 => x"08",
          1072 => x"82",
          1073 => x"fc",
          1074 => x"82",
          1075 => x"fc",
          1076 => x"b5",
          1077 => x"05",
          1078 => x"bf",
          1079 => x"72",
          1080 => x"08",
          1081 => x"81",
          1082 => x"0b",
          1083 => x"08",
          1084 => x"a9",
          1085 => x"b4",
          1086 => x"22",
          1087 => x"07",
          1088 => x"82",
          1089 => x"e4",
          1090 => x"f8",
          1091 => x"b4",
          1092 => x"34",
          1093 => x"b5",
          1094 => x"05",
          1095 => x"b4",
          1096 => x"22",
          1097 => x"70",
          1098 => x"51",
          1099 => x"2e",
          1100 => x"b5",
          1101 => x"05",
          1102 => x"b4",
          1103 => x"08",
          1104 => x"b5",
          1105 => x"05",
          1106 => x"82",
          1107 => x"d8",
          1108 => x"a2",
          1109 => x"b4",
          1110 => x"08",
          1111 => x"08",
          1112 => x"84",
          1113 => x"b4",
          1114 => x"0c",
          1115 => x"b5",
          1116 => x"05",
          1117 => x"b5",
          1118 => x"05",
          1119 => x"b4",
          1120 => x"0c",
          1121 => x"08",
          1122 => x"70",
          1123 => x"53",
          1124 => x"b4",
          1125 => x"23",
          1126 => x"0b",
          1127 => x"08",
          1128 => x"82",
          1129 => x"f0",
          1130 => x"b5",
          1131 => x"05",
          1132 => x"b4",
          1133 => x"08",
          1134 => x"54",
          1135 => x"af",
          1136 => x"b5",
          1137 => x"72",
          1138 => x"b5",
          1139 => x"05",
          1140 => x"b4",
          1141 => x"0c",
          1142 => x"08",
          1143 => x"70",
          1144 => x"89",
          1145 => x"38",
          1146 => x"08",
          1147 => x"53",
          1148 => x"82",
          1149 => x"f8",
          1150 => x"15",
          1151 => x"51",
          1152 => x"b5",
          1153 => x"05",
          1154 => x"82",
          1155 => x"f0",
          1156 => x"72",
          1157 => x"51",
          1158 => x"b5",
          1159 => x"05",
          1160 => x"b4",
          1161 => x"08",
          1162 => x"b4",
          1163 => x"33",
          1164 => x"b5",
          1165 => x"05",
          1166 => x"82",
          1167 => x"f0",
          1168 => x"b5",
          1169 => x"05",
          1170 => x"82",
          1171 => x"fc",
          1172 => x"53",
          1173 => x"82",
          1174 => x"70",
          1175 => x"08",
          1176 => x"53",
          1177 => x"08",
          1178 => x"80",
          1179 => x"fe",
          1180 => x"b5",
          1181 => x"05",
          1182 => x"b8",
          1183 => x"54",
          1184 => x"31",
          1185 => x"82",
          1186 => x"fc",
          1187 => x"b5",
          1188 => x"05",
          1189 => x"06",
          1190 => x"80",
          1191 => x"82",
          1192 => x"ec",
          1193 => x"11",
          1194 => x"82",
          1195 => x"ec",
          1196 => x"b5",
          1197 => x"05",
          1198 => x"2a",
          1199 => x"51",
          1200 => x"80",
          1201 => x"38",
          1202 => x"08",
          1203 => x"70",
          1204 => x"b5",
          1205 => x"05",
          1206 => x"b4",
          1207 => x"08",
          1208 => x"b5",
          1209 => x"05",
          1210 => x"b4",
          1211 => x"22",
          1212 => x"90",
          1213 => x"06",
          1214 => x"b5",
          1215 => x"05",
          1216 => x"53",
          1217 => x"b4",
          1218 => x"23",
          1219 => x"b5",
          1220 => x"05",
          1221 => x"53",
          1222 => x"b4",
          1223 => x"23",
          1224 => x"08",
          1225 => x"82",
          1226 => x"ec",
          1227 => x"b5",
          1228 => x"05",
          1229 => x"2a",
          1230 => x"51",
          1231 => x"80",
          1232 => x"38",
          1233 => x"08",
          1234 => x"70",
          1235 => x"98",
          1236 => x"b4",
          1237 => x"33",
          1238 => x"53",
          1239 => x"97",
          1240 => x"b4",
          1241 => x"22",
          1242 => x"51",
          1243 => x"b5",
          1244 => x"05",
          1245 => x"82",
          1246 => x"e8",
          1247 => x"82",
          1248 => x"fc",
          1249 => x"71",
          1250 => x"72",
          1251 => x"08",
          1252 => x"82",
          1253 => x"e4",
          1254 => x"83",
          1255 => x"06",
          1256 => x"72",
          1257 => x"38",
          1258 => x"08",
          1259 => x"70",
          1260 => x"90",
          1261 => x"2c",
          1262 => x"51",
          1263 => x"53",
          1264 => x"b5",
          1265 => x"05",
          1266 => x"31",
          1267 => x"82",
          1268 => x"ec",
          1269 => x"39",
          1270 => x"08",
          1271 => x"70",
          1272 => x"90",
          1273 => x"2c",
          1274 => x"51",
          1275 => x"53",
          1276 => x"b5",
          1277 => x"05",
          1278 => x"31",
          1279 => x"82",
          1280 => x"ec",
          1281 => x"b5",
          1282 => x"05",
          1283 => x"80",
          1284 => x"72",
          1285 => x"b5",
          1286 => x"05",
          1287 => x"54",
          1288 => x"b5",
          1289 => x"05",
          1290 => x"2b",
          1291 => x"51",
          1292 => x"25",
          1293 => x"b5",
          1294 => x"05",
          1295 => x"51",
          1296 => x"d2",
          1297 => x"b4",
          1298 => x"22",
          1299 => x"70",
          1300 => x"51",
          1301 => x"2e",
          1302 => x"b5",
          1303 => x"05",
          1304 => x"51",
          1305 => x"80",
          1306 => x"b5",
          1307 => x"05",
          1308 => x"2a",
          1309 => x"51",
          1310 => x"80",
          1311 => x"82",
          1312 => x"88",
          1313 => x"ab",
          1314 => x"3f",
          1315 => x"b5",
          1316 => x"05",
          1317 => x"2a",
          1318 => x"51",
          1319 => x"80",
          1320 => x"82",
          1321 => x"88",
          1322 => x"a0",
          1323 => x"3f",
          1324 => x"08",
          1325 => x"70",
          1326 => x"81",
          1327 => x"53",
          1328 => x"b1",
          1329 => x"b4",
          1330 => x"08",
          1331 => x"95",
          1332 => x"b5",
          1333 => x"05",
          1334 => x"90",
          1335 => x"06",
          1336 => x"b5",
          1337 => x"05",
          1338 => x"b5",
          1339 => x"05",
          1340 => x"de",
          1341 => x"b4",
          1342 => x"22",
          1343 => x"70",
          1344 => x"51",
          1345 => x"2e",
          1346 => x"b5",
          1347 => x"05",
          1348 => x"54",
          1349 => x"b5",
          1350 => x"05",
          1351 => x"2b",
          1352 => x"51",
          1353 => x"25",
          1354 => x"b5",
          1355 => x"05",
          1356 => x"51",
          1357 => x"d2",
          1358 => x"b4",
          1359 => x"22",
          1360 => x"70",
          1361 => x"51",
          1362 => x"2e",
          1363 => x"b5",
          1364 => x"05",
          1365 => x"54",
          1366 => x"b5",
          1367 => x"05",
          1368 => x"2b",
          1369 => x"51",
          1370 => x"25",
          1371 => x"b5",
          1372 => x"05",
          1373 => x"51",
          1374 => x"d2",
          1375 => x"b4",
          1376 => x"22",
          1377 => x"70",
          1378 => x"51",
          1379 => x"38",
          1380 => x"08",
          1381 => x"ff",
          1382 => x"72",
          1383 => x"08",
          1384 => x"73",
          1385 => x"90",
          1386 => x"80",
          1387 => x"38",
          1388 => x"08",
          1389 => x"52",
          1390 => x"96",
          1391 => x"82",
          1392 => x"f8",
          1393 => x"72",
          1394 => x"09",
          1395 => x"38",
          1396 => x"08",
          1397 => x"52",
          1398 => x"08",
          1399 => x"51",
          1400 => x"81",
          1401 => x"b5",
          1402 => x"05",
          1403 => x"80",
          1404 => x"81",
          1405 => x"38",
          1406 => x"08",
          1407 => x"ff",
          1408 => x"72",
          1409 => x"08",
          1410 => x"72",
          1411 => x"06",
          1412 => x"ff",
          1413 => x"bb",
          1414 => x"b4",
          1415 => x"08",
          1416 => x"b4",
          1417 => x"08",
          1418 => x"82",
          1419 => x"fc",
          1420 => x"05",
          1421 => x"08",
          1422 => x"53",
          1423 => x"ff",
          1424 => x"b5",
          1425 => x"05",
          1426 => x"80",
          1427 => x"81",
          1428 => x"38",
          1429 => x"08",
          1430 => x"ff",
          1431 => x"72",
          1432 => x"08",
          1433 => x"72",
          1434 => x"06",
          1435 => x"ff",
          1436 => x"df",
          1437 => x"b4",
          1438 => x"08",
          1439 => x"b4",
          1440 => x"08",
          1441 => x"53",
          1442 => x"82",
          1443 => x"fc",
          1444 => x"05",
          1445 => x"08",
          1446 => x"ff",
          1447 => x"b5",
          1448 => x"05",
          1449 => x"b8",
          1450 => x"82",
          1451 => x"88",
          1452 => x"82",
          1453 => x"f0",
          1454 => x"05",
          1455 => x"08",
          1456 => x"82",
          1457 => x"f0",
          1458 => x"33",
          1459 => x"82",
          1460 => x"82",
          1461 => x"e4",
          1462 => x"87",
          1463 => x"06",
          1464 => x"72",
          1465 => x"c3",
          1466 => x"b4",
          1467 => x"22",
          1468 => x"54",
          1469 => x"b4",
          1470 => x"23",
          1471 => x"70",
          1472 => x"53",
          1473 => x"a3",
          1474 => x"b4",
          1475 => x"08",
          1476 => x"90",
          1477 => x"39",
          1478 => x"08",
          1479 => x"52",
          1480 => x"08",
          1481 => x"51",
          1482 => x"80",
          1483 => x"b4",
          1484 => x"23",
          1485 => x"82",
          1486 => x"f8",
          1487 => x"72",
          1488 => x"81",
          1489 => x"81",
          1490 => x"b4",
          1491 => x"23",
          1492 => x"b5",
          1493 => x"05",
          1494 => x"82",
          1495 => x"e8",
          1496 => x"0b",
          1497 => x"08",
          1498 => x"ea",
          1499 => x"b5",
          1500 => x"05",
          1501 => x"b5",
          1502 => x"05",
          1503 => x"d2",
          1504 => x"39",
          1505 => x"08",
          1506 => x"8c",
          1507 => x"82",
          1508 => x"e0",
          1509 => x"53",
          1510 => x"08",
          1511 => x"82",
          1512 => x"95",
          1513 => x"b5",
          1514 => x"82",
          1515 => x"02",
          1516 => x"0c",
          1517 => x"80",
          1518 => x"b4",
          1519 => x"34",
          1520 => x"08",
          1521 => x"53",
          1522 => x"82",
          1523 => x"88",
          1524 => x"08",
          1525 => x"33",
          1526 => x"b5",
          1527 => x"05",
          1528 => x"ff",
          1529 => x"a0",
          1530 => x"06",
          1531 => x"b5",
          1532 => x"05",
          1533 => x"81",
          1534 => x"53",
          1535 => x"b5",
          1536 => x"05",
          1537 => x"ad",
          1538 => x"06",
          1539 => x"0b",
          1540 => x"08",
          1541 => x"82",
          1542 => x"88",
          1543 => x"08",
          1544 => x"0c",
          1545 => x"53",
          1546 => x"b5",
          1547 => x"05",
          1548 => x"b4",
          1549 => x"33",
          1550 => x"2e",
          1551 => x"81",
          1552 => x"b5",
          1553 => x"05",
          1554 => x"81",
          1555 => x"70",
          1556 => x"72",
          1557 => x"b4",
          1558 => x"34",
          1559 => x"08",
          1560 => x"82",
          1561 => x"e8",
          1562 => x"b5",
          1563 => x"05",
          1564 => x"2e",
          1565 => x"b5",
          1566 => x"05",
          1567 => x"2e",
          1568 => x"cd",
          1569 => x"82",
          1570 => x"f4",
          1571 => x"b5",
          1572 => x"05",
          1573 => x"81",
          1574 => x"70",
          1575 => x"72",
          1576 => x"b4",
          1577 => x"34",
          1578 => x"82",
          1579 => x"b4",
          1580 => x"34",
          1581 => x"08",
          1582 => x"70",
          1583 => x"71",
          1584 => x"51",
          1585 => x"82",
          1586 => x"f8",
          1587 => x"fe",
          1588 => x"b4",
          1589 => x"33",
          1590 => x"26",
          1591 => x"0b",
          1592 => x"08",
          1593 => x"83",
          1594 => x"b5",
          1595 => x"05",
          1596 => x"73",
          1597 => x"82",
          1598 => x"f8",
          1599 => x"72",
          1600 => x"38",
          1601 => x"0b",
          1602 => x"08",
          1603 => x"82",
          1604 => x"0b",
          1605 => x"08",
          1606 => x"b2",
          1607 => x"b4",
          1608 => x"33",
          1609 => x"27",
          1610 => x"b5",
          1611 => x"05",
          1612 => x"b9",
          1613 => x"8d",
          1614 => x"82",
          1615 => x"ec",
          1616 => x"a5",
          1617 => x"82",
          1618 => x"f4",
          1619 => x"0b",
          1620 => x"08",
          1621 => x"82",
          1622 => x"f8",
          1623 => x"a0",
          1624 => x"cf",
          1625 => x"b4",
          1626 => x"33",
          1627 => x"73",
          1628 => x"82",
          1629 => x"f8",
          1630 => x"11",
          1631 => x"82",
          1632 => x"f8",
          1633 => x"b5",
          1634 => x"05",
          1635 => x"51",
          1636 => x"b5",
          1637 => x"05",
          1638 => x"b4",
          1639 => x"33",
          1640 => x"27",
          1641 => x"b5",
          1642 => x"05",
          1643 => x"51",
          1644 => x"b5",
          1645 => x"05",
          1646 => x"b4",
          1647 => x"33",
          1648 => x"26",
          1649 => x"0b",
          1650 => x"08",
          1651 => x"81",
          1652 => x"b5",
          1653 => x"05",
          1654 => x"b4",
          1655 => x"33",
          1656 => x"74",
          1657 => x"80",
          1658 => x"b4",
          1659 => x"0c",
          1660 => x"82",
          1661 => x"f4",
          1662 => x"82",
          1663 => x"fc",
          1664 => x"82",
          1665 => x"f8",
          1666 => x"12",
          1667 => x"08",
          1668 => x"82",
          1669 => x"88",
          1670 => x"08",
          1671 => x"0c",
          1672 => x"51",
          1673 => x"72",
          1674 => x"b4",
          1675 => x"34",
          1676 => x"82",
          1677 => x"f0",
          1678 => x"72",
          1679 => x"38",
          1680 => x"08",
          1681 => x"30",
          1682 => x"08",
          1683 => x"82",
          1684 => x"8c",
          1685 => x"b5",
          1686 => x"05",
          1687 => x"53",
          1688 => x"b5",
          1689 => x"05",
          1690 => x"b4",
          1691 => x"08",
          1692 => x"0c",
          1693 => x"82",
          1694 => x"04",
          1695 => x"08",
          1696 => x"b4",
          1697 => x"0d",
          1698 => x"08",
          1699 => x"b4",
          1700 => x"08",
          1701 => x"b4",
          1702 => x"08",
          1703 => x"3f",
          1704 => x"08",
          1705 => x"a8",
          1706 => x"3d",
          1707 => x"b4",
          1708 => x"b5",
          1709 => x"82",
          1710 => x"f7",
          1711 => x"0b",
          1712 => x"08",
          1713 => x"82",
          1714 => x"8c",
          1715 => x"80",
          1716 => x"b5",
          1717 => x"05",
          1718 => x"51",
          1719 => x"53",
          1720 => x"b4",
          1721 => x"34",
          1722 => x"06",
          1723 => x"2e",
          1724 => x"91",
          1725 => x"b4",
          1726 => x"08",
          1727 => x"05",
          1728 => x"ce",
          1729 => x"b4",
          1730 => x"33",
          1731 => x"2e",
          1732 => x"a4",
          1733 => x"82",
          1734 => x"f0",
          1735 => x"b5",
          1736 => x"05",
          1737 => x"81",
          1738 => x"70",
          1739 => x"72",
          1740 => x"b4",
          1741 => x"34",
          1742 => x"08",
          1743 => x"53",
          1744 => x"09",
          1745 => x"dc",
          1746 => x"b4",
          1747 => x"08",
          1748 => x"05",
          1749 => x"08",
          1750 => x"33",
          1751 => x"08",
          1752 => x"82",
          1753 => x"f8",
          1754 => x"b5",
          1755 => x"05",
          1756 => x"b4",
          1757 => x"08",
          1758 => x"b6",
          1759 => x"b4",
          1760 => x"08",
          1761 => x"84",
          1762 => x"39",
          1763 => x"b5",
          1764 => x"05",
          1765 => x"b4",
          1766 => x"08",
          1767 => x"05",
          1768 => x"08",
          1769 => x"33",
          1770 => x"08",
          1771 => x"81",
          1772 => x"0b",
          1773 => x"08",
          1774 => x"82",
          1775 => x"88",
          1776 => x"08",
          1777 => x"0c",
          1778 => x"53",
          1779 => x"b5",
          1780 => x"05",
          1781 => x"39",
          1782 => x"08",
          1783 => x"53",
          1784 => x"8d",
          1785 => x"82",
          1786 => x"ec",
          1787 => x"80",
          1788 => x"b4",
          1789 => x"33",
          1790 => x"27",
          1791 => x"b5",
          1792 => x"05",
          1793 => x"b9",
          1794 => x"8d",
          1795 => x"82",
          1796 => x"ec",
          1797 => x"d8",
          1798 => x"82",
          1799 => x"f4",
          1800 => x"39",
          1801 => x"08",
          1802 => x"53",
          1803 => x"90",
          1804 => x"b4",
          1805 => x"33",
          1806 => x"26",
          1807 => x"39",
          1808 => x"b5",
          1809 => x"05",
          1810 => x"39",
          1811 => x"b5",
          1812 => x"05",
          1813 => x"82",
          1814 => x"fc",
          1815 => x"b5",
          1816 => x"05",
          1817 => x"73",
          1818 => x"38",
          1819 => x"08",
          1820 => x"53",
          1821 => x"27",
          1822 => x"b5",
          1823 => x"05",
          1824 => x"51",
          1825 => x"b5",
          1826 => x"05",
          1827 => x"b4",
          1828 => x"33",
          1829 => x"53",
          1830 => x"b4",
          1831 => x"34",
          1832 => x"08",
          1833 => x"53",
          1834 => x"ad",
          1835 => x"b4",
          1836 => x"33",
          1837 => x"53",
          1838 => x"b4",
          1839 => x"34",
          1840 => x"08",
          1841 => x"53",
          1842 => x"8d",
          1843 => x"82",
          1844 => x"ec",
          1845 => x"98",
          1846 => x"b4",
          1847 => x"33",
          1848 => x"08",
          1849 => x"54",
          1850 => x"26",
          1851 => x"0b",
          1852 => x"08",
          1853 => x"80",
          1854 => x"b5",
          1855 => x"05",
          1856 => x"b5",
          1857 => x"05",
          1858 => x"b5",
          1859 => x"05",
          1860 => x"82",
          1861 => x"fc",
          1862 => x"b5",
          1863 => x"05",
          1864 => x"81",
          1865 => x"70",
          1866 => x"52",
          1867 => x"33",
          1868 => x"08",
          1869 => x"fe",
          1870 => x"b5",
          1871 => x"05",
          1872 => x"80",
          1873 => x"82",
          1874 => x"fc",
          1875 => x"82",
          1876 => x"fc",
          1877 => x"b5",
          1878 => x"05",
          1879 => x"b4",
          1880 => x"08",
          1881 => x"81",
          1882 => x"b4",
          1883 => x"0c",
          1884 => x"08",
          1885 => x"82",
          1886 => x"8b",
          1887 => x"b5",
          1888 => x"82",
          1889 => x"02",
          1890 => x"0c",
          1891 => x"80",
          1892 => x"b4",
          1893 => x"0c",
          1894 => x"08",
          1895 => x"70",
          1896 => x"81",
          1897 => x"06",
          1898 => x"51",
          1899 => x"2e",
          1900 => x"0b",
          1901 => x"08",
          1902 => x"81",
          1903 => x"b5",
          1904 => x"05",
          1905 => x"33",
          1906 => x"08",
          1907 => x"81",
          1908 => x"b4",
          1909 => x"0c",
          1910 => x"b5",
          1911 => x"05",
          1912 => x"ff",
          1913 => x"80",
          1914 => x"82",
          1915 => x"82",
          1916 => x"53",
          1917 => x"08",
          1918 => x"52",
          1919 => x"51",
          1920 => x"82",
          1921 => x"53",
          1922 => x"ff",
          1923 => x"0b",
          1924 => x"08",
          1925 => x"ff",
          1926 => x"cc",
          1927 => x"cc",
          1928 => x"53",
          1929 => x"13",
          1930 => x"2d",
          1931 => x"08",
          1932 => x"2e",
          1933 => x"0b",
          1934 => x"08",
          1935 => x"82",
          1936 => x"f8",
          1937 => x"82",
          1938 => x"f4",
          1939 => x"82",
          1940 => x"f4",
          1941 => x"b5",
          1942 => x"3d",
          1943 => x"b4",
          1944 => x"b5",
          1945 => x"82",
          1946 => x"fb",
          1947 => x"0b",
          1948 => x"08",
          1949 => x"82",
          1950 => x"8c",
          1951 => x"11",
          1952 => x"2a",
          1953 => x"70",
          1954 => x"51",
          1955 => x"72",
          1956 => x"38",
          1957 => x"b5",
          1958 => x"05",
          1959 => x"39",
          1960 => x"08",
          1961 => x"53",
          1962 => x"b5",
          1963 => x"05",
          1964 => x"82",
          1965 => x"88",
          1966 => x"72",
          1967 => x"08",
          1968 => x"72",
          1969 => x"53",
          1970 => x"b6",
          1971 => x"b4",
          1972 => x"08",
          1973 => x"08",
          1974 => x"53",
          1975 => x"08",
          1976 => x"52",
          1977 => x"51",
          1978 => x"82",
          1979 => x"53",
          1980 => x"ff",
          1981 => x"0b",
          1982 => x"08",
          1983 => x"ff",
          1984 => x"b5",
          1985 => x"05",
          1986 => x"b5",
          1987 => x"05",
          1988 => x"b5",
          1989 => x"05",
          1990 => x"a8",
          1991 => x"0d",
          1992 => x"0c",
          1993 => x"b4",
          1994 => x"b5",
          1995 => x"3d",
          1996 => x"fc",
          1997 => x"b5",
          1998 => x"05",
          1999 => x"3f",
          2000 => x"08",
          2001 => x"a8",
          2002 => x"3d",
          2003 => x"b4",
          2004 => x"b5",
          2005 => x"82",
          2006 => x"fb",
          2007 => x"b5",
          2008 => x"05",
          2009 => x"33",
          2010 => x"70",
          2011 => x"81",
          2012 => x"51",
          2013 => x"80",
          2014 => x"ff",
          2015 => x"b4",
          2016 => x"0c",
          2017 => x"82",
          2018 => x"8c",
          2019 => x"11",
          2020 => x"2a",
          2021 => x"51",
          2022 => x"72",
          2023 => x"db",
          2024 => x"b4",
          2025 => x"08",
          2026 => x"08",
          2027 => x"54",
          2028 => x"08",
          2029 => x"25",
          2030 => x"b5",
          2031 => x"05",
          2032 => x"70",
          2033 => x"08",
          2034 => x"52",
          2035 => x"72",
          2036 => x"08",
          2037 => x"0c",
          2038 => x"08",
          2039 => x"8c",
          2040 => x"05",
          2041 => x"82",
          2042 => x"88",
          2043 => x"82",
          2044 => x"fc",
          2045 => x"53",
          2046 => x"82",
          2047 => x"8c",
          2048 => x"b5",
          2049 => x"05",
          2050 => x"b5",
          2051 => x"05",
          2052 => x"ff",
          2053 => x"12",
          2054 => x"54",
          2055 => x"b5",
          2056 => x"72",
          2057 => x"b5",
          2058 => x"05",
          2059 => x"08",
          2060 => x"12",
          2061 => x"b4",
          2062 => x"08",
          2063 => x"b4",
          2064 => x"0c",
          2065 => x"39",
          2066 => x"b5",
          2067 => x"05",
          2068 => x"b4",
          2069 => x"08",
          2070 => x"0c",
          2071 => x"82",
          2072 => x"04",
          2073 => x"08",
          2074 => x"b4",
          2075 => x"0d",
          2076 => x"08",
          2077 => x"85",
          2078 => x"81",
          2079 => x"06",
          2080 => x"52",
          2081 => x"8d",
          2082 => x"82",
          2083 => x"f8",
          2084 => x"94",
          2085 => x"b4",
          2086 => x"08",
          2087 => x"70",
          2088 => x"81",
          2089 => x"51",
          2090 => x"2e",
          2091 => x"82",
          2092 => x"88",
          2093 => x"b5",
          2094 => x"05",
          2095 => x"85",
          2096 => x"ff",
          2097 => x"52",
          2098 => x"34",
          2099 => x"08",
          2100 => x"8c",
          2101 => x"05",
          2102 => x"82",
          2103 => x"88",
          2104 => x"11",
          2105 => x"b5",
          2106 => x"05",
          2107 => x"52",
          2108 => x"82",
          2109 => x"88",
          2110 => x"11",
          2111 => x"2a",
          2112 => x"51",
          2113 => x"71",
          2114 => x"d7",
          2115 => x"b4",
          2116 => x"08",
          2117 => x"33",
          2118 => x"08",
          2119 => x"51",
          2120 => x"b4",
          2121 => x"08",
          2122 => x"b5",
          2123 => x"05",
          2124 => x"b4",
          2125 => x"08",
          2126 => x"12",
          2127 => x"07",
          2128 => x"85",
          2129 => x"0b",
          2130 => x"08",
          2131 => x"81",
          2132 => x"b5",
          2133 => x"05",
          2134 => x"81",
          2135 => x"52",
          2136 => x"82",
          2137 => x"88",
          2138 => x"b5",
          2139 => x"05",
          2140 => x"11",
          2141 => x"71",
          2142 => x"a8",
          2143 => x"b5",
          2144 => x"05",
          2145 => x"b5",
          2146 => x"05",
          2147 => x"80",
          2148 => x"b5",
          2149 => x"05",
          2150 => x"b4",
          2151 => x"0c",
          2152 => x"08",
          2153 => x"85",
          2154 => x"b5",
          2155 => x"05",
          2156 => x"b5",
          2157 => x"05",
          2158 => x"09",
          2159 => x"38",
          2160 => x"08",
          2161 => x"90",
          2162 => x"82",
          2163 => x"ec",
          2164 => x"39",
          2165 => x"08",
          2166 => x"a0",
          2167 => x"82",
          2168 => x"ec",
          2169 => x"b5",
          2170 => x"05",
          2171 => x"b5",
          2172 => x"05",
          2173 => x"34",
          2174 => x"b5",
          2175 => x"05",
          2176 => x"82",
          2177 => x"88",
          2178 => x"11",
          2179 => x"8c",
          2180 => x"b5",
          2181 => x"05",
          2182 => x"ff",
          2183 => x"b5",
          2184 => x"05",
          2185 => x"52",
          2186 => x"08",
          2187 => x"82",
          2188 => x"89",
          2189 => x"b5",
          2190 => x"82",
          2191 => x"02",
          2192 => x"0c",
          2193 => x"82",
          2194 => x"88",
          2195 => x"b5",
          2196 => x"05",
          2197 => x"b4",
          2198 => x"08",
          2199 => x"08",
          2200 => x"82",
          2201 => x"90",
          2202 => x"2e",
          2203 => x"82",
          2204 => x"f8",
          2205 => x"b5",
          2206 => x"05",
          2207 => x"ac",
          2208 => x"b4",
          2209 => x"08",
          2210 => x"08",
          2211 => x"05",
          2212 => x"b4",
          2213 => x"08",
          2214 => x"90",
          2215 => x"b4",
          2216 => x"08",
          2217 => x"08",
          2218 => x"05",
          2219 => x"08",
          2220 => x"82",
          2221 => x"f8",
          2222 => x"b5",
          2223 => x"05",
          2224 => x"b5",
          2225 => x"05",
          2226 => x"b4",
          2227 => x"08",
          2228 => x"b5",
          2229 => x"05",
          2230 => x"b4",
          2231 => x"08",
          2232 => x"b5",
          2233 => x"05",
          2234 => x"b4",
          2235 => x"08",
          2236 => x"9c",
          2237 => x"b4",
          2238 => x"08",
          2239 => x"b5",
          2240 => x"05",
          2241 => x"b4",
          2242 => x"08",
          2243 => x"b5",
          2244 => x"05",
          2245 => x"b4",
          2246 => x"08",
          2247 => x"08",
          2248 => x"53",
          2249 => x"71",
          2250 => x"39",
          2251 => x"08",
          2252 => x"81",
          2253 => x"b4",
          2254 => x"0c",
          2255 => x"08",
          2256 => x"ff",
          2257 => x"b4",
          2258 => x"0c",
          2259 => x"08",
          2260 => x"80",
          2261 => x"82",
          2262 => x"f8",
          2263 => x"70",
          2264 => x"b4",
          2265 => x"08",
          2266 => x"b5",
          2267 => x"05",
          2268 => x"b4",
          2269 => x"08",
          2270 => x"71",
          2271 => x"b4",
          2272 => x"08",
          2273 => x"b5",
          2274 => x"05",
          2275 => x"39",
          2276 => x"08",
          2277 => x"70",
          2278 => x"0c",
          2279 => x"0d",
          2280 => x"0c",
          2281 => x"b4",
          2282 => x"b5",
          2283 => x"3d",
          2284 => x"b4",
          2285 => x"08",
          2286 => x"08",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"71",
          2290 => x"b4",
          2291 => x"08",
          2292 => x"b5",
          2293 => x"05",
          2294 => x"ff",
          2295 => x"70",
          2296 => x"38",
          2297 => x"b5",
          2298 => x"05",
          2299 => x"82",
          2300 => x"fc",
          2301 => x"b5",
          2302 => x"05",
          2303 => x"b4",
          2304 => x"08",
          2305 => x"b5",
          2306 => x"84",
          2307 => x"b5",
          2308 => x"82",
          2309 => x"02",
          2310 => x"0c",
          2311 => x"82",
          2312 => x"88",
          2313 => x"b5",
          2314 => x"05",
          2315 => x"b4",
          2316 => x"08",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"05",
          2320 => x"08",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"51",
          2324 => x"82",
          2325 => x"fc",
          2326 => x"05",
          2327 => x"08",
          2328 => x"70",
          2329 => x"51",
          2330 => x"84",
          2331 => x"39",
          2332 => x"08",
          2333 => x"70",
          2334 => x"0c",
          2335 => x"0d",
          2336 => x"0c",
          2337 => x"b4",
          2338 => x"b5",
          2339 => x"3d",
          2340 => x"b4",
          2341 => x"08",
          2342 => x"08",
          2343 => x"82",
          2344 => x"8c",
          2345 => x"b5",
          2346 => x"05",
          2347 => x"b4",
          2348 => x"08",
          2349 => x"e5",
          2350 => x"b4",
          2351 => x"08",
          2352 => x"b5",
          2353 => x"05",
          2354 => x"b4",
          2355 => x"08",
          2356 => x"b5",
          2357 => x"05",
          2358 => x"b4",
          2359 => x"08",
          2360 => x"38",
          2361 => x"08",
          2362 => x"51",
          2363 => x"b5",
          2364 => x"05",
          2365 => x"82",
          2366 => x"f8",
          2367 => x"b5",
          2368 => x"05",
          2369 => x"71",
          2370 => x"b5",
          2371 => x"05",
          2372 => x"82",
          2373 => x"fc",
          2374 => x"ad",
          2375 => x"b4",
          2376 => x"08",
          2377 => x"a8",
          2378 => x"3d",
          2379 => x"b4",
          2380 => x"b5",
          2381 => x"82",
          2382 => x"fd",
          2383 => x"b5",
          2384 => x"05",
          2385 => x"81",
          2386 => x"b5",
          2387 => x"05",
          2388 => x"33",
          2389 => x"08",
          2390 => x"81",
          2391 => x"b4",
          2392 => x"0c",
          2393 => x"08",
          2394 => x"70",
          2395 => x"ff",
          2396 => x"54",
          2397 => x"2e",
          2398 => x"ce",
          2399 => x"b4",
          2400 => x"08",
          2401 => x"82",
          2402 => x"88",
          2403 => x"05",
          2404 => x"08",
          2405 => x"70",
          2406 => x"51",
          2407 => x"38",
          2408 => x"b5",
          2409 => x"05",
          2410 => x"39",
          2411 => x"08",
          2412 => x"ff",
          2413 => x"b4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"ff",
          2418 => x"b5",
          2419 => x"05",
          2420 => x"80",
          2421 => x"b5",
          2422 => x"05",
          2423 => x"52",
          2424 => x"38",
          2425 => x"b5",
          2426 => x"05",
          2427 => x"39",
          2428 => x"08",
          2429 => x"ff",
          2430 => x"b4",
          2431 => x"0c",
          2432 => x"08",
          2433 => x"70",
          2434 => x"70",
          2435 => x"0b",
          2436 => x"08",
          2437 => x"ae",
          2438 => x"b4",
          2439 => x"08",
          2440 => x"b5",
          2441 => x"05",
          2442 => x"72",
          2443 => x"82",
          2444 => x"fc",
          2445 => x"55",
          2446 => x"8a",
          2447 => x"82",
          2448 => x"fc",
          2449 => x"b5",
          2450 => x"05",
          2451 => x"a8",
          2452 => x"0d",
          2453 => x"0c",
          2454 => x"b4",
          2455 => x"b5",
          2456 => x"3d",
          2457 => x"b4",
          2458 => x"08",
          2459 => x"08",
          2460 => x"82",
          2461 => x"8c",
          2462 => x"38",
          2463 => x"b5",
          2464 => x"05",
          2465 => x"39",
          2466 => x"08",
          2467 => x"52",
          2468 => x"b5",
          2469 => x"05",
          2470 => x"82",
          2471 => x"f8",
          2472 => x"81",
          2473 => x"51",
          2474 => x"9f",
          2475 => x"b4",
          2476 => x"08",
          2477 => x"b5",
          2478 => x"05",
          2479 => x"b4",
          2480 => x"08",
          2481 => x"38",
          2482 => x"82",
          2483 => x"f8",
          2484 => x"05",
          2485 => x"08",
          2486 => x"82",
          2487 => x"f8",
          2488 => x"b5",
          2489 => x"05",
          2490 => x"82",
          2491 => x"fc",
          2492 => x"82",
          2493 => x"fc",
          2494 => x"b5",
          2495 => x"3d",
          2496 => x"b4",
          2497 => x"b5",
          2498 => x"82",
          2499 => x"fe",
          2500 => x"b5",
          2501 => x"05",
          2502 => x"b4",
          2503 => x"0c",
          2504 => x"08",
          2505 => x"80",
          2506 => x"38",
          2507 => x"08",
          2508 => x"81",
          2509 => x"b4",
          2510 => x"0c",
          2511 => x"08",
          2512 => x"ff",
          2513 => x"b4",
          2514 => x"0c",
          2515 => x"08",
          2516 => x"80",
          2517 => x"82",
          2518 => x"8c",
          2519 => x"70",
          2520 => x"08",
          2521 => x"52",
          2522 => x"34",
          2523 => x"08",
          2524 => x"81",
          2525 => x"b4",
          2526 => x"0c",
          2527 => x"82",
          2528 => x"88",
          2529 => x"82",
          2530 => x"51",
          2531 => x"82",
          2532 => x"04",
          2533 => x"08",
          2534 => x"b4",
          2535 => x"0d",
          2536 => x"b5",
          2537 => x"05",
          2538 => x"b4",
          2539 => x"08",
          2540 => x"38",
          2541 => x"08",
          2542 => x"30",
          2543 => x"08",
          2544 => x"80",
          2545 => x"b4",
          2546 => x"0c",
          2547 => x"08",
          2548 => x"8a",
          2549 => x"82",
          2550 => x"f4",
          2551 => x"b5",
          2552 => x"05",
          2553 => x"b4",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"80",
          2557 => x"82",
          2558 => x"8c",
          2559 => x"82",
          2560 => x"8c",
          2561 => x"0b",
          2562 => x"08",
          2563 => x"82",
          2564 => x"fc",
          2565 => x"38",
          2566 => x"b5",
          2567 => x"05",
          2568 => x"b4",
          2569 => x"08",
          2570 => x"08",
          2571 => x"80",
          2572 => x"b4",
          2573 => x"08",
          2574 => x"b4",
          2575 => x"08",
          2576 => x"3f",
          2577 => x"08",
          2578 => x"b4",
          2579 => x"0c",
          2580 => x"b4",
          2581 => x"08",
          2582 => x"38",
          2583 => x"08",
          2584 => x"30",
          2585 => x"08",
          2586 => x"82",
          2587 => x"f8",
          2588 => x"82",
          2589 => x"54",
          2590 => x"82",
          2591 => x"04",
          2592 => x"08",
          2593 => x"b4",
          2594 => x"0d",
          2595 => x"b5",
          2596 => x"05",
          2597 => x"b4",
          2598 => x"08",
          2599 => x"38",
          2600 => x"08",
          2601 => x"30",
          2602 => x"08",
          2603 => x"81",
          2604 => x"b4",
          2605 => x"0c",
          2606 => x"08",
          2607 => x"80",
          2608 => x"82",
          2609 => x"8c",
          2610 => x"82",
          2611 => x"8c",
          2612 => x"53",
          2613 => x"08",
          2614 => x"52",
          2615 => x"08",
          2616 => x"51",
          2617 => x"82",
          2618 => x"70",
          2619 => x"08",
          2620 => x"54",
          2621 => x"08",
          2622 => x"80",
          2623 => x"82",
          2624 => x"f8",
          2625 => x"82",
          2626 => x"f8",
          2627 => x"b5",
          2628 => x"05",
          2629 => x"b5",
          2630 => x"87",
          2631 => x"b5",
          2632 => x"82",
          2633 => x"02",
          2634 => x"0c",
          2635 => x"80",
          2636 => x"b4",
          2637 => x"08",
          2638 => x"b4",
          2639 => x"08",
          2640 => x"3f",
          2641 => x"08",
          2642 => x"a8",
          2643 => x"3d",
          2644 => x"b4",
          2645 => x"b5",
          2646 => x"82",
          2647 => x"fd",
          2648 => x"53",
          2649 => x"08",
          2650 => x"52",
          2651 => x"08",
          2652 => x"51",
          2653 => x"b5",
          2654 => x"82",
          2655 => x"54",
          2656 => x"82",
          2657 => x"04",
          2658 => x"08",
          2659 => x"b4",
          2660 => x"0d",
          2661 => x"b5",
          2662 => x"05",
          2663 => x"82",
          2664 => x"f8",
          2665 => x"b5",
          2666 => x"05",
          2667 => x"b4",
          2668 => x"08",
          2669 => x"82",
          2670 => x"fc",
          2671 => x"2e",
          2672 => x"0b",
          2673 => x"08",
          2674 => x"24",
          2675 => x"b5",
          2676 => x"05",
          2677 => x"b5",
          2678 => x"05",
          2679 => x"b4",
          2680 => x"08",
          2681 => x"b4",
          2682 => x"0c",
          2683 => x"82",
          2684 => x"fc",
          2685 => x"2e",
          2686 => x"82",
          2687 => x"8c",
          2688 => x"b5",
          2689 => x"05",
          2690 => x"38",
          2691 => x"08",
          2692 => x"82",
          2693 => x"8c",
          2694 => x"82",
          2695 => x"88",
          2696 => x"b5",
          2697 => x"05",
          2698 => x"b4",
          2699 => x"08",
          2700 => x"b4",
          2701 => x"0c",
          2702 => x"08",
          2703 => x"81",
          2704 => x"b4",
          2705 => x"0c",
          2706 => x"08",
          2707 => x"81",
          2708 => x"b4",
          2709 => x"0c",
          2710 => x"82",
          2711 => x"90",
          2712 => x"2e",
          2713 => x"b5",
          2714 => x"05",
          2715 => x"b5",
          2716 => x"05",
          2717 => x"39",
          2718 => x"08",
          2719 => x"70",
          2720 => x"08",
          2721 => x"51",
          2722 => x"08",
          2723 => x"82",
          2724 => x"85",
          2725 => x"b5",
          2726 => x"f9",
          2727 => x"70",
          2728 => x"56",
          2729 => x"2e",
          2730 => x"95",
          2731 => x"51",
          2732 => x"82",
          2733 => x"15",
          2734 => x"16",
          2735 => x"cd",
          2736 => x"54",
          2737 => x"09",
          2738 => x"38",
          2739 => x"f1",
          2740 => x"76",
          2741 => x"b0",
          2742 => x"08",
          2743 => x"c5",
          2744 => x"a8",
          2745 => x"52",
          2746 => x"f4",
          2747 => x"b5",
          2748 => x"38",
          2749 => x"54",
          2750 => x"ff",
          2751 => x"17",
          2752 => x"06",
          2753 => x"77",
          2754 => x"ff",
          2755 => x"b5",
          2756 => x"3d",
          2757 => x"3d",
          2758 => x"71",
          2759 => x"8e",
          2760 => x"29",
          2761 => x"05",
          2762 => x"04",
          2763 => x"51",
          2764 => x"82",
          2765 => x"80",
          2766 => x"9a",
          2767 => x"f2",
          2768 => x"c0",
          2769 => x"39",
          2770 => x"51",
          2771 => x"82",
          2772 => x"80",
          2773 => x"9a",
          2774 => x"d6",
          2775 => x"84",
          2776 => x"39",
          2777 => x"51",
          2778 => x"82",
          2779 => x"80",
          2780 => x"9b",
          2781 => x"39",
          2782 => x"51",
          2783 => x"9b",
          2784 => x"39",
          2785 => x"51",
          2786 => x"9c",
          2787 => x"39",
          2788 => x"51",
          2789 => x"9c",
          2790 => x"39",
          2791 => x"51",
          2792 => x"9d",
          2793 => x"39",
          2794 => x"51",
          2795 => x"9d",
          2796 => x"cf",
          2797 => x"0d",
          2798 => x"0d",
          2799 => x"56",
          2800 => x"26",
          2801 => x"52",
          2802 => x"29",
          2803 => x"87",
          2804 => x"51",
          2805 => x"82",
          2806 => x"52",
          2807 => x"c3",
          2808 => x"a8",
          2809 => x"53",
          2810 => x"9d",
          2811 => x"bb",
          2812 => x"3d",
          2813 => x"3d",
          2814 => x"84",
          2815 => x"05",
          2816 => x"80",
          2817 => x"70",
          2818 => x"25",
          2819 => x"59",
          2820 => x"87",
          2821 => x"38",
          2822 => x"76",
          2823 => x"ff",
          2824 => x"93",
          2825 => x"82",
          2826 => x"76",
          2827 => x"70",
          2828 => x"fe",
          2829 => x"b5",
          2830 => x"82",
          2831 => x"b9",
          2832 => x"a8",
          2833 => x"98",
          2834 => x"b5",
          2835 => x"96",
          2836 => x"54",
          2837 => x"77",
          2838 => x"81",
          2839 => x"82",
          2840 => x"57",
          2841 => x"08",
          2842 => x"55",
          2843 => x"89",
          2844 => x"75",
          2845 => x"d7",
          2846 => x"d8",
          2847 => x"8b",
          2848 => x"30",
          2849 => x"80",
          2850 => x"70",
          2851 => x"06",
          2852 => x"56",
          2853 => x"90",
          2854 => x"f8",
          2855 => x"98",
          2856 => x"78",
          2857 => x"3f",
          2858 => x"82",
          2859 => x"96",
          2860 => x"f8",
          2861 => x"02",
          2862 => x"05",
          2863 => x"ff",
          2864 => x"7b",
          2865 => x"fe",
          2866 => x"b5",
          2867 => x"38",
          2868 => x"88",
          2869 => x"2e",
          2870 => x"39",
          2871 => x"55",
          2872 => x"b5",
          2873 => x"52",
          2874 => x"2d",
          2875 => x"08",
          2876 => x"78",
          2877 => x"b5",
          2878 => x"3d",
          2879 => x"3d",
          2880 => x"63",
          2881 => x"80",
          2882 => x"73",
          2883 => x"41",
          2884 => x"5e",
          2885 => x"52",
          2886 => x"51",
          2887 => x"3f",
          2888 => x"51",
          2889 => x"80",
          2890 => x"27",
          2891 => x"7b",
          2892 => x"38",
          2893 => x"a6",
          2894 => x"39",
          2895 => x"72",
          2896 => x"38",
          2897 => x"82",
          2898 => x"ff",
          2899 => x"88",
          2900 => x"98",
          2901 => x"3f",
          2902 => x"80",
          2903 => x"18",
          2904 => x"27",
          2905 => x"08",
          2906 => x"80",
          2907 => x"e6",
          2908 => x"82",
          2909 => x"e0",
          2910 => x"15",
          2911 => x"74",
          2912 => x"7a",
          2913 => x"72",
          2914 => x"9e",
          2915 => x"b8",
          2916 => x"39",
          2917 => x"51",
          2918 => x"81",
          2919 => x"cc",
          2920 => x"a0",
          2921 => x"3f",
          2922 => x"82",
          2923 => x"df",
          2924 => x"55",
          2925 => x"80",
          2926 => x"18",
          2927 => x"53",
          2928 => x"7a",
          2929 => x"81",
          2930 => x"9f",
          2931 => x"38",
          2932 => x"73",
          2933 => x"ff",
          2934 => x"72",
          2935 => x"38",
          2936 => x"26",
          2937 => x"cc",
          2938 => x"73",
          2939 => x"82",
          2940 => x"52",
          2941 => x"da",
          2942 => x"55",
          2943 => x"82",
          2944 => x"de",
          2945 => x"18",
          2946 => x"58",
          2947 => x"82",
          2948 => x"98",
          2949 => x"2c",
          2950 => x"a0",
          2951 => x"06",
          2952 => x"aa",
          2953 => x"a8",
          2954 => x"70",
          2955 => x"a0",
          2956 => x"72",
          2957 => x"30",
          2958 => x"73",
          2959 => x"51",
          2960 => x"57",
          2961 => x"73",
          2962 => x"76",
          2963 => x"81",
          2964 => x"80",
          2965 => x"7c",
          2966 => x"78",
          2967 => x"38",
          2968 => x"82",
          2969 => x"8f",
          2970 => x"fc",
          2971 => x"9b",
          2972 => x"9e",
          2973 => x"9e",
          2974 => x"ff",
          2975 => x"82",
          2976 => x"51",
          2977 => x"82",
          2978 => x"82",
          2979 => x"82",
          2980 => x"52",
          2981 => x"51",
          2982 => x"3f",
          2983 => x"84",
          2984 => x"3f",
          2985 => x"04",
          2986 => x"87",
          2987 => x"08",
          2988 => x"3f",
          2989 => x"83",
          2990 => x"f4",
          2991 => x"3f",
          2992 => x"f7",
          2993 => x"2a",
          2994 => x"51",
          2995 => x"2e",
          2996 => x"51",
          2997 => x"82",
          2998 => x"98",
          2999 => x"51",
          3000 => x"72",
          3001 => x"81",
          3002 => x"71",
          3003 => x"38",
          3004 => x"c7",
          3005 => x"a0",
          3006 => x"3f",
          3007 => x"bb",
          3008 => x"2a",
          3009 => x"51",
          3010 => x"2e",
          3011 => x"51",
          3012 => x"82",
          3013 => x"98",
          3014 => x"51",
          3015 => x"72",
          3016 => x"81",
          3017 => x"71",
          3018 => x"38",
          3019 => x"8b",
          3020 => x"c4",
          3021 => x"3f",
          3022 => x"ff",
          3023 => x"2a",
          3024 => x"51",
          3025 => x"2e",
          3026 => x"51",
          3027 => x"82",
          3028 => x"98",
          3029 => x"51",
          3030 => x"72",
          3031 => x"81",
          3032 => x"71",
          3033 => x"38",
          3034 => x"cf",
          3035 => x"ec",
          3036 => x"3f",
          3037 => x"c3",
          3038 => x"2a",
          3039 => x"51",
          3040 => x"2e",
          3041 => x"51",
          3042 => x"82",
          3043 => x"97",
          3044 => x"51",
          3045 => x"72",
          3046 => x"81",
          3047 => x"71",
          3048 => x"38",
          3049 => x"93",
          3050 => x"94",
          3051 => x"3f",
          3052 => x"87",
          3053 => x"3f",
          3054 => x"04",
          3055 => x"77",
          3056 => x"a3",
          3057 => x"55",
          3058 => x"52",
          3059 => x"b6",
          3060 => x"82",
          3061 => x"54",
          3062 => x"81",
          3063 => x"d4",
          3064 => x"a8",
          3065 => x"a9",
          3066 => x"a8",
          3067 => x"82",
          3068 => x"07",
          3069 => x"71",
          3070 => x"54",
          3071 => x"82",
          3072 => x"0b",
          3073 => x"a4",
          3074 => x"81",
          3075 => x"06",
          3076 => x"cc",
          3077 => x"52",
          3078 => x"b1",
          3079 => x"b5",
          3080 => x"2e",
          3081 => x"b5",
          3082 => x"da",
          3083 => x"39",
          3084 => x"51",
          3085 => x"3f",
          3086 => x"0b",
          3087 => x"34",
          3088 => x"b0",
          3089 => x"73",
          3090 => x"81",
          3091 => x"82",
          3092 => x"74",
          3093 => x"a9",
          3094 => x"0b",
          3095 => x"0c",
          3096 => x"04",
          3097 => x"80",
          3098 => x"cc",
          3099 => x"5e",
          3100 => x"51",
          3101 => x"3f",
          3102 => x"08",
          3103 => x"5a",
          3104 => x"09",
          3105 => x"38",
          3106 => x"83",
          3107 => x"ec",
          3108 => x"e7",
          3109 => x"53",
          3110 => x"b6",
          3111 => x"f5",
          3112 => x"b5",
          3113 => x"2e",
          3114 => x"a0",
          3115 => x"95",
          3116 => x"40",
          3117 => x"a8",
          3118 => x"3f",
          3119 => x"47",
          3120 => x"52",
          3121 => x"f4",
          3122 => x"ff",
          3123 => x"f3",
          3124 => x"b5",
          3125 => x"2b",
          3126 => x"51",
          3127 => x"c2",
          3128 => x"38",
          3129 => x"24",
          3130 => x"bd",
          3131 => x"38",
          3132 => x"90",
          3133 => x"2e",
          3134 => x"79",
          3135 => x"da",
          3136 => x"39",
          3137 => x"2e",
          3138 => x"79",
          3139 => x"85",
          3140 => x"bf",
          3141 => x"38",
          3142 => x"79",
          3143 => x"89",
          3144 => x"80",
          3145 => x"38",
          3146 => x"2e",
          3147 => x"79",
          3148 => x"89",
          3149 => x"8b",
          3150 => x"83",
          3151 => x"38",
          3152 => x"24",
          3153 => x"81",
          3154 => x"d7",
          3155 => x"39",
          3156 => x"2e",
          3157 => x"89",
          3158 => x"3d",
          3159 => x"53",
          3160 => x"51",
          3161 => x"82",
          3162 => x"80",
          3163 => x"38",
          3164 => x"fc",
          3165 => x"84",
          3166 => x"b6",
          3167 => x"a8",
          3168 => x"fe",
          3169 => x"3d",
          3170 => x"53",
          3171 => x"51",
          3172 => x"82",
          3173 => x"86",
          3174 => x"a8",
          3175 => x"a1",
          3176 => x"df",
          3177 => x"5d",
          3178 => x"27",
          3179 => x"62",
          3180 => x"70",
          3181 => x"0c",
          3182 => x"f5",
          3183 => x"39",
          3184 => x"80",
          3185 => x"84",
          3186 => x"e6",
          3187 => x"a8",
          3188 => x"fd",
          3189 => x"3d",
          3190 => x"53",
          3191 => x"51",
          3192 => x"82",
          3193 => x"80",
          3194 => x"38",
          3195 => x"f8",
          3196 => x"84",
          3197 => x"ba",
          3198 => x"a8",
          3199 => x"fd",
          3200 => x"a1",
          3201 => x"fb",
          3202 => x"7a",
          3203 => x"88",
          3204 => x"7a",
          3205 => x"5c",
          3206 => x"62",
          3207 => x"eb",
          3208 => x"ff",
          3209 => x"ff",
          3210 => x"d1",
          3211 => x"b5",
          3212 => x"2e",
          3213 => x"b5",
          3214 => x"11",
          3215 => x"05",
          3216 => x"3f",
          3217 => x"08",
          3218 => x"e9",
          3219 => x"fe",
          3220 => x"ff",
          3221 => x"d0",
          3222 => x"b5",
          3223 => x"2e",
          3224 => x"82",
          3225 => x"d6",
          3226 => x"5b",
          3227 => x"a8",
          3228 => x"33",
          3229 => x"5b",
          3230 => x"2e",
          3231 => x"55",
          3232 => x"33",
          3233 => x"82",
          3234 => x"ff",
          3235 => x"81",
          3236 => x"05",
          3237 => x"39",
          3238 => x"51",
          3239 => x"b5",
          3240 => x"11",
          3241 => x"05",
          3242 => x"3f",
          3243 => x"08",
          3244 => x"82",
          3245 => x"5a",
          3246 => x"89",
          3247 => x"cc",
          3248 => x"cd",
          3249 => x"95",
          3250 => x"80",
          3251 => x"82",
          3252 => x"45",
          3253 => x"b4",
          3254 => x"79",
          3255 => x"38",
          3256 => x"08",
          3257 => x"82",
          3258 => x"5a",
          3259 => x"88",
          3260 => x"e4",
          3261 => x"39",
          3262 => x"33",
          3263 => x"2e",
          3264 => x"b3",
          3265 => x"89",
          3266 => x"fc",
          3267 => x"05",
          3268 => x"fe",
          3269 => x"ff",
          3270 => x"cf",
          3271 => x"b5",
          3272 => x"de",
          3273 => x"94",
          3274 => x"80",
          3275 => x"82",
          3276 => x"44",
          3277 => x"82",
          3278 => x"5a",
          3279 => x"88",
          3280 => x"d8",
          3281 => x"39",
          3282 => x"33",
          3283 => x"2e",
          3284 => x"b3",
          3285 => x"aa",
          3286 => x"97",
          3287 => x"80",
          3288 => x"82",
          3289 => x"44",
          3290 => x"b4",
          3291 => x"79",
          3292 => x"38",
          3293 => x"08",
          3294 => x"82",
          3295 => x"88",
          3296 => x"3d",
          3297 => x"53",
          3298 => x"51",
          3299 => x"82",
          3300 => x"80",
          3301 => x"80",
          3302 => x"7b",
          3303 => x"38",
          3304 => x"90",
          3305 => x"70",
          3306 => x"2a",
          3307 => x"51",
          3308 => x"79",
          3309 => x"38",
          3310 => x"83",
          3311 => x"82",
          3312 => x"d3",
          3313 => x"55",
          3314 => x"53",
          3315 => x"51",
          3316 => x"82",
          3317 => x"86",
          3318 => x"3d",
          3319 => x"53",
          3320 => x"51",
          3321 => x"82",
          3322 => x"80",
          3323 => x"38",
          3324 => x"fc",
          3325 => x"84",
          3326 => x"b6",
          3327 => x"a8",
          3328 => x"a4",
          3329 => x"02",
          3330 => x"33",
          3331 => x"81",
          3332 => x"3d",
          3333 => x"53",
          3334 => x"51",
          3335 => x"82",
          3336 => x"e1",
          3337 => x"39",
          3338 => x"54",
          3339 => x"90",
          3340 => x"a2",
          3341 => x"52",
          3342 => x"c0",
          3343 => x"7a",
          3344 => x"ae",
          3345 => x"38",
          3346 => x"9f",
          3347 => x"fe",
          3348 => x"ff",
          3349 => x"cc",
          3350 => x"b5",
          3351 => x"2e",
          3352 => x"5a",
          3353 => x"05",
          3354 => x"64",
          3355 => x"ff",
          3356 => x"a2",
          3357 => x"8b",
          3358 => x"39",
          3359 => x"f4",
          3360 => x"84",
          3361 => x"a3",
          3362 => x"a8",
          3363 => x"f8",
          3364 => x"3d",
          3365 => x"53",
          3366 => x"51",
          3367 => x"82",
          3368 => x"80",
          3369 => x"61",
          3370 => x"c2",
          3371 => x"70",
          3372 => x"23",
          3373 => x"3d",
          3374 => x"53",
          3375 => x"51",
          3376 => x"82",
          3377 => x"df",
          3378 => x"39",
          3379 => x"54",
          3380 => x"a4",
          3381 => x"fe",
          3382 => x"52",
          3383 => x"9c",
          3384 => x"7a",
          3385 => x"ae",
          3386 => x"38",
          3387 => x"87",
          3388 => x"05",
          3389 => x"b5",
          3390 => x"11",
          3391 => x"05",
          3392 => x"3f",
          3393 => x"08",
          3394 => x"38",
          3395 => x"80",
          3396 => x"7a",
          3397 => x"5c",
          3398 => x"ff",
          3399 => x"a2",
          3400 => x"df",
          3401 => x"39",
          3402 => x"f4",
          3403 => x"84",
          3404 => x"f7",
          3405 => x"a8",
          3406 => x"f6",
          3407 => x"3d",
          3408 => x"53",
          3409 => x"51",
          3410 => x"82",
          3411 => x"80",
          3412 => x"61",
          3413 => x"5a",
          3414 => x"42",
          3415 => x"f0",
          3416 => x"84",
          3417 => x"c3",
          3418 => x"a8",
          3419 => x"f6",
          3420 => x"70",
          3421 => x"82",
          3422 => x"ff",
          3423 => x"80",
          3424 => x"51",
          3425 => x"7a",
          3426 => x"5a",
          3427 => x"f6",
          3428 => x"7a",
          3429 => x"b5",
          3430 => x"11",
          3431 => x"05",
          3432 => x"3f",
          3433 => x"08",
          3434 => x"38",
          3435 => x"0c",
          3436 => x"05",
          3437 => x"39",
          3438 => x"51",
          3439 => x"ff",
          3440 => x"3d",
          3441 => x"53",
          3442 => x"51",
          3443 => x"82",
          3444 => x"80",
          3445 => x"38",
          3446 => x"a2",
          3447 => x"a7",
          3448 => x"5a",
          3449 => x"3d",
          3450 => x"53",
          3451 => x"51",
          3452 => x"82",
          3453 => x"80",
          3454 => x"38",
          3455 => x"a2",
          3456 => x"a7",
          3457 => x"5a",
          3458 => x"b5",
          3459 => x"2e",
          3460 => x"82",
          3461 => x"52",
          3462 => x"51",
          3463 => x"3f",
          3464 => x"82",
          3465 => x"ce",
          3466 => x"a7",
          3467 => x"85",
          3468 => x"ac",
          3469 => x"3f",
          3470 => x"a8",
          3471 => x"3f",
          3472 => x"7a",
          3473 => x"5a",
          3474 => x"f4",
          3475 => x"7e",
          3476 => x"80",
          3477 => x"38",
          3478 => x"84",
          3479 => x"d3",
          3480 => x"a8",
          3481 => x"5c",
          3482 => x"b2",
          3483 => x"24",
          3484 => x"81",
          3485 => x"80",
          3486 => x"83",
          3487 => x"80",
          3488 => x"a3",
          3489 => x"55",
          3490 => x"54",
          3491 => x"a3",
          3492 => x"3d",
          3493 => x"51",
          3494 => x"3f",
          3495 => x"a3",
          3496 => x"3d",
          3497 => x"51",
          3498 => x"3f",
          3499 => x"55",
          3500 => x"54",
          3501 => x"a3",
          3502 => x"3d",
          3503 => x"51",
          3504 => x"3f",
          3505 => x"54",
          3506 => x"a3",
          3507 => x"3d",
          3508 => x"51",
          3509 => x"3f",
          3510 => x"59",
          3511 => x"58",
          3512 => x"57",
          3513 => x"55",
          3514 => x"d0",
          3515 => x"d0",
          3516 => x"3d",
          3517 => x"51",
          3518 => x"82",
          3519 => x"82",
          3520 => x"09",
          3521 => x"72",
          3522 => x"51",
          3523 => x"80",
          3524 => x"26",
          3525 => x"5b",
          3526 => x"5a",
          3527 => x"8d",
          3528 => x"70",
          3529 => x"5d",
          3530 => x"bc",
          3531 => x"32",
          3532 => x"07",
          3533 => x"38",
          3534 => x"09",
          3535 => x"f5",
          3536 => x"ec",
          3537 => x"3f",
          3538 => x"f5",
          3539 => x"0b",
          3540 => x"34",
          3541 => x"8c",
          3542 => x"55",
          3543 => x"52",
          3544 => x"bf",
          3545 => x"a8",
          3546 => x"75",
          3547 => x"87",
          3548 => x"73",
          3549 => x"3f",
          3550 => x"a8",
          3551 => x"0c",
          3552 => x"9c",
          3553 => x"55",
          3554 => x"52",
          3555 => x"93",
          3556 => x"a8",
          3557 => x"75",
          3558 => x"87",
          3559 => x"73",
          3560 => x"3f",
          3561 => x"a8",
          3562 => x"0c",
          3563 => x"0b",
          3564 => x"84",
          3565 => x"83",
          3566 => x"94",
          3567 => x"a3",
          3568 => x"bf",
          3569 => x"d3",
          3570 => x"bf",
          3571 => x"84",
          3572 => x"34",
          3573 => x"3d",
          3574 => x"cc",
          3575 => x"c4",
          3576 => x"3f",
          3577 => x"51",
          3578 => x"82",
          3579 => x"cb",
          3580 => x"a4",
          3581 => x"8b",
          3582 => x"a8",
          3583 => x"3f",
          3584 => x"e7",
          3585 => x"3f",
          3586 => x"3d",
          3587 => x"83",
          3588 => x"2b",
          3589 => x"3f",
          3590 => x"08",
          3591 => x"72",
          3592 => x"54",
          3593 => x"25",
          3594 => x"82",
          3595 => x"84",
          3596 => x"fc",
          3597 => x"70",
          3598 => x"80",
          3599 => x"72",
          3600 => x"8a",
          3601 => x"51",
          3602 => x"09",
          3603 => x"38",
          3604 => x"f1",
          3605 => x"51",
          3606 => x"09",
          3607 => x"38",
          3608 => x"81",
          3609 => x"73",
          3610 => x"81",
          3611 => x"84",
          3612 => x"52",
          3613 => x"52",
          3614 => x"2e",
          3615 => x"54",
          3616 => x"9d",
          3617 => x"38",
          3618 => x"12",
          3619 => x"33",
          3620 => x"a0",
          3621 => x"81",
          3622 => x"2e",
          3623 => x"ea",
          3624 => x"33",
          3625 => x"a0",
          3626 => x"06",
          3627 => x"54",
          3628 => x"70",
          3629 => x"25",
          3630 => x"51",
          3631 => x"2e",
          3632 => x"72",
          3633 => x"54",
          3634 => x"0c",
          3635 => x"82",
          3636 => x"86",
          3637 => x"fc",
          3638 => x"53",
          3639 => x"2e",
          3640 => x"3d",
          3641 => x"72",
          3642 => x"bf",
          3643 => x"a8",
          3644 => x"80",
          3645 => x"74",
          3646 => x"b5",
          3647 => x"3d",
          3648 => x"3d",
          3649 => x"11",
          3650 => x"52",
          3651 => x"70",
          3652 => x"98",
          3653 => x"33",
          3654 => x"82",
          3655 => x"26",
          3656 => x"84",
          3657 => x"83",
          3658 => x"26",
          3659 => x"85",
          3660 => x"84",
          3661 => x"26",
          3662 => x"86",
          3663 => x"85",
          3664 => x"26",
          3665 => x"88",
          3666 => x"86",
          3667 => x"e7",
          3668 => x"38",
          3669 => x"54",
          3670 => x"87",
          3671 => x"cc",
          3672 => x"87",
          3673 => x"0c",
          3674 => x"c0",
          3675 => x"82",
          3676 => x"c0",
          3677 => x"83",
          3678 => x"c0",
          3679 => x"84",
          3680 => x"c0",
          3681 => x"85",
          3682 => x"c0",
          3683 => x"86",
          3684 => x"c0",
          3685 => x"74",
          3686 => x"a4",
          3687 => x"c0",
          3688 => x"80",
          3689 => x"98",
          3690 => x"52",
          3691 => x"a8",
          3692 => x"0d",
          3693 => x"0d",
          3694 => x"c0",
          3695 => x"81",
          3696 => x"c0",
          3697 => x"5e",
          3698 => x"87",
          3699 => x"08",
          3700 => x"1c",
          3701 => x"98",
          3702 => x"79",
          3703 => x"87",
          3704 => x"08",
          3705 => x"1c",
          3706 => x"98",
          3707 => x"79",
          3708 => x"87",
          3709 => x"08",
          3710 => x"1c",
          3711 => x"98",
          3712 => x"7b",
          3713 => x"87",
          3714 => x"08",
          3715 => x"1c",
          3716 => x"0c",
          3717 => x"ff",
          3718 => x"83",
          3719 => x"58",
          3720 => x"57",
          3721 => x"56",
          3722 => x"55",
          3723 => x"54",
          3724 => x"53",
          3725 => x"ff",
          3726 => x"a4",
          3727 => x"9f",
          3728 => x"3d",
          3729 => x"3d",
          3730 => x"05",
          3731 => x"c8",
          3732 => x"ff",
          3733 => x"55",
          3734 => x"84",
          3735 => x"2e",
          3736 => x"c0",
          3737 => x"70",
          3738 => x"2a",
          3739 => x"53",
          3740 => x"80",
          3741 => x"71",
          3742 => x"81",
          3743 => x"70",
          3744 => x"81",
          3745 => x"06",
          3746 => x"80",
          3747 => x"71",
          3748 => x"81",
          3749 => x"70",
          3750 => x"73",
          3751 => x"51",
          3752 => x"80",
          3753 => x"2e",
          3754 => x"c0",
          3755 => x"74",
          3756 => x"82",
          3757 => x"87",
          3758 => x"ff",
          3759 => x"8f",
          3760 => x"30",
          3761 => x"51",
          3762 => x"82",
          3763 => x"83",
          3764 => x"f9",
          3765 => x"a7",
          3766 => x"77",
          3767 => x"81",
          3768 => x"7a",
          3769 => x"eb",
          3770 => x"c8",
          3771 => x"ff",
          3772 => x"87",
          3773 => x"53",
          3774 => x"86",
          3775 => x"94",
          3776 => x"08",
          3777 => x"70",
          3778 => x"56",
          3779 => x"2e",
          3780 => x"91",
          3781 => x"06",
          3782 => x"d7",
          3783 => x"32",
          3784 => x"51",
          3785 => x"2e",
          3786 => x"93",
          3787 => x"06",
          3788 => x"ff",
          3789 => x"81",
          3790 => x"87",
          3791 => x"54",
          3792 => x"86",
          3793 => x"94",
          3794 => x"74",
          3795 => x"82",
          3796 => x"89",
          3797 => x"f9",
          3798 => x"54",
          3799 => x"70",
          3800 => x"53",
          3801 => x"77",
          3802 => x"38",
          3803 => x"06",
          3804 => x"b3",
          3805 => x"81",
          3806 => x"57",
          3807 => x"c0",
          3808 => x"75",
          3809 => x"38",
          3810 => x"94",
          3811 => x"70",
          3812 => x"81",
          3813 => x"52",
          3814 => x"8c",
          3815 => x"2a",
          3816 => x"51",
          3817 => x"38",
          3818 => x"70",
          3819 => x"51",
          3820 => x"8d",
          3821 => x"2a",
          3822 => x"51",
          3823 => x"be",
          3824 => x"ff",
          3825 => x"c0",
          3826 => x"70",
          3827 => x"38",
          3828 => x"90",
          3829 => x"0c",
          3830 => x"33",
          3831 => x"06",
          3832 => x"70",
          3833 => x"76",
          3834 => x"0c",
          3835 => x"04",
          3836 => x"82",
          3837 => x"70",
          3838 => x"54",
          3839 => x"94",
          3840 => x"80",
          3841 => x"87",
          3842 => x"51",
          3843 => x"82",
          3844 => x"06",
          3845 => x"70",
          3846 => x"38",
          3847 => x"06",
          3848 => x"94",
          3849 => x"80",
          3850 => x"87",
          3851 => x"52",
          3852 => x"81",
          3853 => x"b5",
          3854 => x"84",
          3855 => x"ff",
          3856 => x"b5",
          3857 => x"ff",
          3858 => x"a8",
          3859 => x"3d",
          3860 => x"c8",
          3861 => x"ff",
          3862 => x"87",
          3863 => x"52",
          3864 => x"86",
          3865 => x"94",
          3866 => x"08",
          3867 => x"70",
          3868 => x"51",
          3869 => x"70",
          3870 => x"38",
          3871 => x"06",
          3872 => x"94",
          3873 => x"80",
          3874 => x"87",
          3875 => x"52",
          3876 => x"98",
          3877 => x"2c",
          3878 => x"71",
          3879 => x"0c",
          3880 => x"04",
          3881 => x"87",
          3882 => x"08",
          3883 => x"8a",
          3884 => x"70",
          3885 => x"b4",
          3886 => x"9e",
          3887 => x"b3",
          3888 => x"c0",
          3889 => x"82",
          3890 => x"87",
          3891 => x"08",
          3892 => x"0c",
          3893 => x"98",
          3894 => x"d8",
          3895 => x"9e",
          3896 => x"b3",
          3897 => x"c0",
          3898 => x"82",
          3899 => x"87",
          3900 => x"08",
          3901 => x"0c",
          3902 => x"b0",
          3903 => x"e8",
          3904 => x"9e",
          3905 => x"b3",
          3906 => x"c0",
          3907 => x"82",
          3908 => x"87",
          3909 => x"08",
          3910 => x"0c",
          3911 => x"c0",
          3912 => x"f8",
          3913 => x"9e",
          3914 => x"b3",
          3915 => x"c0",
          3916 => x"51",
          3917 => x"80",
          3918 => x"9e",
          3919 => x"b4",
          3920 => x"c0",
          3921 => x"82",
          3922 => x"87",
          3923 => x"08",
          3924 => x"0c",
          3925 => x"b4",
          3926 => x"0b",
          3927 => x"90",
          3928 => x"80",
          3929 => x"52",
          3930 => x"2e",
          3931 => x"52",
          3932 => x"91",
          3933 => x"87",
          3934 => x"08",
          3935 => x"0a",
          3936 => x"52",
          3937 => x"83",
          3938 => x"71",
          3939 => x"34",
          3940 => x"c0",
          3941 => x"70",
          3942 => x"06",
          3943 => x"70",
          3944 => x"38",
          3945 => x"82",
          3946 => x"80",
          3947 => x"9e",
          3948 => x"88",
          3949 => x"51",
          3950 => x"80",
          3951 => x"81",
          3952 => x"b4",
          3953 => x"0b",
          3954 => x"90",
          3955 => x"80",
          3956 => x"52",
          3957 => x"2e",
          3958 => x"52",
          3959 => x"95",
          3960 => x"87",
          3961 => x"08",
          3962 => x"80",
          3963 => x"52",
          3964 => x"83",
          3965 => x"71",
          3966 => x"34",
          3967 => x"c0",
          3968 => x"70",
          3969 => x"06",
          3970 => x"70",
          3971 => x"38",
          3972 => x"82",
          3973 => x"80",
          3974 => x"9e",
          3975 => x"82",
          3976 => x"51",
          3977 => x"80",
          3978 => x"81",
          3979 => x"b4",
          3980 => x"0b",
          3981 => x"90",
          3982 => x"80",
          3983 => x"52",
          3984 => x"2e",
          3985 => x"52",
          3986 => x"99",
          3987 => x"87",
          3988 => x"08",
          3989 => x"80",
          3990 => x"52",
          3991 => x"83",
          3992 => x"71",
          3993 => x"34",
          3994 => x"c0",
          3995 => x"70",
          3996 => x"51",
          3997 => x"80",
          3998 => x"81",
          3999 => x"b4",
          4000 => x"c0",
          4001 => x"70",
          4002 => x"70",
          4003 => x"51",
          4004 => x"b4",
          4005 => x"0b",
          4006 => x"90",
          4007 => x"80",
          4008 => x"52",
          4009 => x"83",
          4010 => x"71",
          4011 => x"34",
          4012 => x"90",
          4013 => x"f0",
          4014 => x"2a",
          4015 => x"70",
          4016 => x"34",
          4017 => x"c0",
          4018 => x"70",
          4019 => x"52",
          4020 => x"2e",
          4021 => x"52",
          4022 => x"9f",
          4023 => x"9e",
          4024 => x"87",
          4025 => x"70",
          4026 => x"34",
          4027 => x"04",
          4028 => x"82",
          4029 => x"ff",
          4030 => x"82",
          4031 => x"54",
          4032 => x"89",
          4033 => x"f4",
          4034 => x"f7",
          4035 => x"88",
          4036 => x"ef",
          4037 => x"92",
          4038 => x"80",
          4039 => x"82",
          4040 => x"82",
          4041 => x"11",
          4042 => x"a5",
          4043 => x"95",
          4044 => x"b4",
          4045 => x"73",
          4046 => x"38",
          4047 => x"08",
          4048 => x"08",
          4049 => x"82",
          4050 => x"ff",
          4051 => x"82",
          4052 => x"54",
          4053 => x"94",
          4054 => x"cc",
          4055 => x"d0",
          4056 => x"52",
          4057 => x"51",
          4058 => x"3f",
          4059 => x"33",
          4060 => x"2e",
          4061 => x"b3",
          4062 => x"b3",
          4063 => x"54",
          4064 => x"f4",
          4065 => x"ce",
          4066 => x"96",
          4067 => x"80",
          4068 => x"82",
          4069 => x"82",
          4070 => x"11",
          4071 => x"a6",
          4072 => x"94",
          4073 => x"b4",
          4074 => x"73",
          4075 => x"38",
          4076 => x"33",
          4077 => x"ac",
          4078 => x"9a",
          4079 => x"9f",
          4080 => x"80",
          4081 => x"82",
          4082 => x"52",
          4083 => x"51",
          4084 => x"3f",
          4085 => x"33",
          4086 => x"2e",
          4087 => x"b4",
          4088 => x"82",
          4089 => x"ff",
          4090 => x"82",
          4091 => x"54",
          4092 => x"89",
          4093 => x"8c",
          4094 => x"87",
          4095 => x"93",
          4096 => x"80",
          4097 => x"82",
          4098 => x"ff",
          4099 => x"82",
          4100 => x"54",
          4101 => x"89",
          4102 => x"ac",
          4103 => x"e3",
          4104 => x"99",
          4105 => x"80",
          4106 => x"82",
          4107 => x"ff",
          4108 => x"82",
          4109 => x"54",
          4110 => x"89",
          4111 => x"c4",
          4112 => x"bf",
          4113 => x"d0",
          4114 => x"b7",
          4115 => x"f4",
          4116 => x"a7",
          4117 => x"92",
          4118 => x"b3",
          4119 => x"82",
          4120 => x"ff",
          4121 => x"82",
          4122 => x"52",
          4123 => x"51",
          4124 => x"3f",
          4125 => x"51",
          4126 => x"3f",
          4127 => x"22",
          4128 => x"dc",
          4129 => x"ce",
          4130 => x"84",
          4131 => x"84",
          4132 => x"51",
          4133 => x"82",
          4134 => x"bd",
          4135 => x"76",
          4136 => x"54",
          4137 => x"08",
          4138 => x"84",
          4139 => x"a6",
          4140 => x"97",
          4141 => x"80",
          4142 => x"82",
          4143 => x"56",
          4144 => x"52",
          4145 => x"db",
          4146 => x"a8",
          4147 => x"c0",
          4148 => x"31",
          4149 => x"b5",
          4150 => x"82",
          4151 => x"ff",
          4152 => x"82",
          4153 => x"54",
          4154 => x"a9",
          4155 => x"8c",
          4156 => x"84",
          4157 => x"51",
          4158 => x"82",
          4159 => x"bd",
          4160 => x"76",
          4161 => x"54",
          4162 => x"08",
          4163 => x"dc",
          4164 => x"c2",
          4165 => x"f0",
          4166 => x"e7",
          4167 => x"0d",
          4168 => x"0d",
          4169 => x"33",
          4170 => x"71",
          4171 => x"38",
          4172 => x"82",
          4173 => x"52",
          4174 => x"82",
          4175 => x"9d",
          4176 => x"90",
          4177 => x"82",
          4178 => x"91",
          4179 => x"a0",
          4180 => x"82",
          4181 => x"85",
          4182 => x"ac",
          4183 => x"a3",
          4184 => x"0d",
          4185 => x"80",
          4186 => x"0b",
          4187 => x"84",
          4188 => x"b4",
          4189 => x"c0",
          4190 => x"04",
          4191 => x"76",
          4192 => x"98",
          4193 => x"2b",
          4194 => x"72",
          4195 => x"82",
          4196 => x"51",
          4197 => x"80",
          4198 => x"b8",
          4199 => x"53",
          4200 => x"9c",
          4201 => x"b4",
          4202 => x"02",
          4203 => x"05",
          4204 => x"52",
          4205 => x"72",
          4206 => x"06",
          4207 => x"53",
          4208 => x"a8",
          4209 => x"0d",
          4210 => x"0d",
          4211 => x"05",
          4212 => x"71",
          4213 => x"53",
          4214 => x"a2",
          4215 => x"ff",
          4216 => x"a0",
          4217 => x"bd",
          4218 => x"ff",
          4219 => x"72",
          4220 => x"52",
          4221 => x"71",
          4222 => x"52",
          4223 => x"51",
          4224 => x"3f",
          4225 => x"86",
          4226 => x"f6",
          4227 => x"02",
          4228 => x"05",
          4229 => x"05",
          4230 => x"82",
          4231 => x"70",
          4232 => x"b4",
          4233 => x"08",
          4234 => x"5a",
          4235 => x"80",
          4236 => x"74",
          4237 => x"3f",
          4238 => x"33",
          4239 => x"82",
          4240 => x"81",
          4241 => x"58",
          4242 => x"b3",
          4243 => x"a8",
          4244 => x"82",
          4245 => x"70",
          4246 => x"b4",
          4247 => x"08",
          4248 => x"74",
          4249 => x"38",
          4250 => x"52",
          4251 => x"95",
          4252 => x"80",
          4253 => x"55",
          4254 => x"80",
          4255 => x"ff",
          4256 => x"75",
          4257 => x"80",
          4258 => x"80",
          4259 => x"2e",
          4260 => x"b4",
          4261 => x"75",
          4262 => x"38",
          4263 => x"33",
          4264 => x"38",
          4265 => x"05",
          4266 => x"78",
          4267 => x"80",
          4268 => x"82",
          4269 => x"52",
          4270 => x"8e",
          4271 => x"b4",
          4272 => x"80",
          4273 => x"8c",
          4274 => x"fd",
          4275 => x"b4",
          4276 => x"54",
          4277 => x"71",
          4278 => x"38",
          4279 => x"89",
          4280 => x"0c",
          4281 => x"14",
          4282 => x"80",
          4283 => x"80",
          4284 => x"80",
          4285 => x"fc",
          4286 => x"80",
          4287 => x"71",
          4288 => x"fe",
          4289 => x"fc",
          4290 => x"dd",
          4291 => x"82",
          4292 => x"85",
          4293 => x"dc",
          4294 => x"57",
          4295 => x"b4",
          4296 => x"80",
          4297 => x"82",
          4298 => x"80",
          4299 => x"b4",
          4300 => x"80",
          4301 => x"3d",
          4302 => x"81",
          4303 => x"82",
          4304 => x"80",
          4305 => x"75",
          4306 => x"3f",
          4307 => x"08",
          4308 => x"82",
          4309 => x"25",
          4310 => x"b5",
          4311 => x"05",
          4312 => x"55",
          4313 => x"75",
          4314 => x"81",
          4315 => x"a8",
          4316 => x"8c",
          4317 => x"ff",
          4318 => x"06",
          4319 => x"a6",
          4320 => x"d9",
          4321 => x"3d",
          4322 => x"08",
          4323 => x"70",
          4324 => x"52",
          4325 => x"08",
          4326 => x"f5",
          4327 => x"a8",
          4328 => x"38",
          4329 => x"b4",
          4330 => x"55",
          4331 => x"8b",
          4332 => x"56",
          4333 => x"3f",
          4334 => x"08",
          4335 => x"38",
          4336 => x"bf",
          4337 => x"b5",
          4338 => x"18",
          4339 => x"0b",
          4340 => x"08",
          4341 => x"82",
          4342 => x"ff",
          4343 => x"55",
          4344 => x"34",
          4345 => x"30",
          4346 => x"9f",
          4347 => x"55",
          4348 => x"85",
          4349 => x"ac",
          4350 => x"fc",
          4351 => x"08",
          4352 => x"e1",
          4353 => x"b5",
          4354 => x"2e",
          4355 => x"ad",
          4356 => x"b2",
          4357 => x"77",
          4358 => x"06",
          4359 => x"52",
          4360 => x"bf",
          4361 => x"51",
          4362 => x"3f",
          4363 => x"54",
          4364 => x"08",
          4365 => x"58",
          4366 => x"a8",
          4367 => x"0d",
          4368 => x"0d",
          4369 => x"5c",
          4370 => x"57",
          4371 => x"73",
          4372 => x"81",
          4373 => x"78",
          4374 => x"56",
          4375 => x"98",
          4376 => x"70",
          4377 => x"33",
          4378 => x"73",
          4379 => x"81",
          4380 => x"75",
          4381 => x"38",
          4382 => x"88",
          4383 => x"84",
          4384 => x"52",
          4385 => x"9d",
          4386 => x"a8",
          4387 => x"52",
          4388 => x"c1",
          4389 => x"b5",
          4390 => x"c6",
          4391 => x"33",
          4392 => x"2e",
          4393 => x"82",
          4394 => x"b6",
          4395 => x"3f",
          4396 => x"1a",
          4397 => x"fc",
          4398 => x"05",
          4399 => x"f2",
          4400 => x"a8",
          4401 => x"9a",
          4402 => x"53",
          4403 => x"51",
          4404 => x"82",
          4405 => x"81",
          4406 => x"74",
          4407 => x"54",
          4408 => x"14",
          4409 => x"06",
          4410 => x"74",
          4411 => x"38",
          4412 => x"82",
          4413 => x"8c",
          4414 => x"d3",
          4415 => x"3d",
          4416 => x"08",
          4417 => x"59",
          4418 => x"0b",
          4419 => x"82",
          4420 => x"82",
          4421 => x"55",
          4422 => x"cb",
          4423 => x"b4",
          4424 => x"55",
          4425 => x"81",
          4426 => x"2e",
          4427 => x"81",
          4428 => x"55",
          4429 => x"2e",
          4430 => x"a8",
          4431 => x"3f",
          4432 => x"08",
          4433 => x"0c",
          4434 => x"08",
          4435 => x"92",
          4436 => x"76",
          4437 => x"a8",
          4438 => x"cc",
          4439 => x"b5",
          4440 => x"2e",
          4441 => x"ad",
          4442 => x"b0",
          4443 => x"f7",
          4444 => x"a8",
          4445 => x"b4",
          4446 => x"80",
          4447 => x"3d",
          4448 => x"81",
          4449 => x"82",
          4450 => x"56",
          4451 => x"08",
          4452 => x"81",
          4453 => x"38",
          4454 => x"08",
          4455 => x"85",
          4456 => x"a8",
          4457 => x"0b",
          4458 => x"08",
          4459 => x"82",
          4460 => x"ff",
          4461 => x"55",
          4462 => x"34",
          4463 => x"81",
          4464 => x"75",
          4465 => x"3f",
          4466 => x"81",
          4467 => x"54",
          4468 => x"83",
          4469 => x"74",
          4470 => x"81",
          4471 => x"38",
          4472 => x"82",
          4473 => x"76",
          4474 => x"b4",
          4475 => x"2e",
          4476 => x"d7",
          4477 => x"5d",
          4478 => x"82",
          4479 => x"98",
          4480 => x"2c",
          4481 => x"ff",
          4482 => x"78",
          4483 => x"82",
          4484 => x"70",
          4485 => x"98",
          4486 => x"d0",
          4487 => x"2b",
          4488 => x"71",
          4489 => x"70",
          4490 => x"aa",
          4491 => x"08",
          4492 => x"51",
          4493 => x"59",
          4494 => x"5d",
          4495 => x"73",
          4496 => x"e9",
          4497 => x"27",
          4498 => x"81",
          4499 => x"81",
          4500 => x"70",
          4501 => x"55",
          4502 => x"80",
          4503 => x"53",
          4504 => x"51",
          4505 => x"82",
          4506 => x"81",
          4507 => x"73",
          4508 => x"38",
          4509 => x"d0",
          4510 => x"b1",
          4511 => x"80",
          4512 => x"80",
          4513 => x"98",
          4514 => x"ff",
          4515 => x"55",
          4516 => x"97",
          4517 => x"74",
          4518 => x"f5",
          4519 => x"b5",
          4520 => x"ff",
          4521 => x"cc",
          4522 => x"80",
          4523 => x"2e",
          4524 => x"81",
          4525 => x"82",
          4526 => x"74",
          4527 => x"98",
          4528 => x"d0",
          4529 => x"2b",
          4530 => x"70",
          4531 => x"82",
          4532 => x"b8",
          4533 => x"51",
          4534 => x"58",
          4535 => x"77",
          4536 => x"06",
          4537 => x"82",
          4538 => x"08",
          4539 => x"0b",
          4540 => x"34",
          4541 => x"cc",
          4542 => x"39",
          4543 => x"d4",
          4544 => x"cc",
          4545 => x"af",
          4546 => x"7d",
          4547 => x"73",
          4548 => x"e1",
          4549 => x"29",
          4550 => x"05",
          4551 => x"04",
          4552 => x"33",
          4553 => x"2e",
          4554 => x"82",
          4555 => x"55",
          4556 => x"ab",
          4557 => x"2b",
          4558 => x"51",
          4559 => x"24",
          4560 => x"1a",
          4561 => x"81",
          4562 => x"81",
          4563 => x"81",
          4564 => x"70",
          4565 => x"cc",
          4566 => x"51",
          4567 => x"82",
          4568 => x"81",
          4569 => x"74",
          4570 => x"34",
          4571 => x"ae",
          4572 => x"34",
          4573 => x"33",
          4574 => x"25",
          4575 => x"14",
          4576 => x"cc",
          4577 => x"cc",
          4578 => x"81",
          4579 => x"81",
          4580 => x"70",
          4581 => x"cc",
          4582 => x"51",
          4583 => x"77",
          4584 => x"74",
          4585 => x"52",
          4586 => x"f9",
          4587 => x"80",
          4588 => x"80",
          4589 => x"98",
          4590 => x"d8",
          4591 => x"55",
          4592 => x"df",
          4593 => x"dc",
          4594 => x"2b",
          4595 => x"82",
          4596 => x"5a",
          4597 => x"74",
          4598 => x"99",
          4599 => x"ff",
          4600 => x"74",
          4601 => x"29",
          4602 => x"05",
          4603 => x"82",
          4604 => x"56",
          4605 => x"75",
          4606 => x"fb",
          4607 => x"7a",
          4608 => x"81",
          4609 => x"cc",
          4610 => x"52",
          4611 => x"51",
          4612 => x"81",
          4613 => x"cc",
          4614 => x"81",
          4615 => x"55",
          4616 => x"fb",
          4617 => x"cc",
          4618 => x"05",
          4619 => x"cc",
          4620 => x"15",
          4621 => x"cc",
          4622 => x"51",
          4623 => x"3f",
          4624 => x"33",
          4625 => x"70",
          4626 => x"cc",
          4627 => x"51",
          4628 => x"74",
          4629 => x"74",
          4630 => x"14",
          4631 => x"73",
          4632 => x"ad",
          4633 => x"81",
          4634 => x"81",
          4635 => x"70",
          4636 => x"cc",
          4637 => x"51",
          4638 => x"24",
          4639 => x"51",
          4640 => x"3f",
          4641 => x"33",
          4642 => x"70",
          4643 => x"cc",
          4644 => x"51",
          4645 => x"74",
          4646 => x"38",
          4647 => x"ad",
          4648 => x"81",
          4649 => x"81",
          4650 => x"70",
          4651 => x"cc",
          4652 => x"51",
          4653 => x"25",
          4654 => x"b9",
          4655 => x"d8",
          4656 => x"54",
          4657 => x"8a",
          4658 => x"d9",
          4659 => x"d8",
          4660 => x"f6",
          4661 => x"b5",
          4662 => x"ff",
          4663 => x"96",
          4664 => x"d8",
          4665 => x"80",
          4666 => x"81",
          4667 => x"79",
          4668 => x"3f",
          4669 => x"7a",
          4670 => x"82",
          4671 => x"80",
          4672 => x"d8",
          4673 => x"b5",
          4674 => x"3d",
          4675 => x"cc",
          4676 => x"73",
          4677 => x"dd",
          4678 => x"ff",
          4679 => x"82",
          4680 => x"ff",
          4681 => x"82",
          4682 => x"73",
          4683 => x"54",
          4684 => x"cc",
          4685 => x"cc",
          4686 => x"55",
          4687 => x"f9",
          4688 => x"14",
          4689 => x"cc",
          4690 => x"98",
          4691 => x"2c",
          4692 => x"06",
          4693 => x"74",
          4694 => x"38",
          4695 => x"81",
          4696 => x"34",
          4697 => x"ff",
          4698 => x"74",
          4699 => x"29",
          4700 => x"05",
          4701 => x"82",
          4702 => x"58",
          4703 => x"75",
          4704 => x"a0",
          4705 => x"9d",
          4706 => x"dc",
          4707 => x"2b",
          4708 => x"82",
          4709 => x"57",
          4710 => x"74",
          4711 => x"d5",
          4712 => x"ff",
          4713 => x"74",
          4714 => x"29",
          4715 => x"05",
          4716 => x"82",
          4717 => x"58",
          4718 => x"75",
          4719 => x"f8",
          4720 => x"cc",
          4721 => x"81",
          4722 => x"cc",
          4723 => x"56",
          4724 => x"27",
          4725 => x"81",
          4726 => x"82",
          4727 => x"74",
          4728 => x"52",
          4729 => x"bd",
          4730 => x"dc",
          4731 => x"ff",
          4732 => x"d8",
          4733 => x"54",
          4734 => x"db",
          4735 => x"39",
          4736 => x"53",
          4737 => x"a2",
          4738 => x"bd",
          4739 => x"82",
          4740 => x"80",
          4741 => x"d8",
          4742 => x"39",
          4743 => x"82",
          4744 => x"55",
          4745 => x"a6",
          4746 => x"ff",
          4747 => x"82",
          4748 => x"82",
          4749 => x"82",
          4750 => x"81",
          4751 => x"05",
          4752 => x"79",
          4753 => x"bd",
          4754 => x"81",
          4755 => x"84",
          4756 => x"a8",
          4757 => x"08",
          4758 => x"80",
          4759 => x"74",
          4760 => x"c1",
          4761 => x"a8",
          4762 => x"d8",
          4763 => x"a8",
          4764 => x"06",
          4765 => x"74",
          4766 => x"ff",
          4767 => x"ff",
          4768 => x"fa",
          4769 => x"55",
          4770 => x"f6",
          4771 => x"51",
          4772 => x"3f",
          4773 => x"93",
          4774 => x"06",
          4775 => x"b4",
          4776 => x"74",
          4777 => x"38",
          4778 => x"b1",
          4779 => x"b5",
          4780 => x"cc",
          4781 => x"b5",
          4782 => x"ff",
          4783 => x"53",
          4784 => x"51",
          4785 => x"3f",
          4786 => x"7a",
          4787 => x"b4",
          4788 => x"08",
          4789 => x"80",
          4790 => x"74",
          4791 => x"c5",
          4792 => x"a8",
          4793 => x"d8",
          4794 => x"a8",
          4795 => x"06",
          4796 => x"74",
          4797 => x"ff",
          4798 => x"81",
          4799 => x"81",
          4800 => x"89",
          4801 => x"cc",
          4802 => x"7a",
          4803 => x"dc",
          4804 => x"d8",
          4805 => x"51",
          4806 => x"f5",
          4807 => x"cc",
          4808 => x"81",
          4809 => x"cc",
          4810 => x"56",
          4811 => x"27",
          4812 => x"81",
          4813 => x"82",
          4814 => x"74",
          4815 => x"52",
          4816 => x"e1",
          4817 => x"39",
          4818 => x"33",
          4819 => x"2e",
          4820 => x"88",
          4821 => x"cd",
          4822 => x"dc",
          4823 => x"54",
          4824 => x"dc",
          4825 => x"39",
          4826 => x"83",
          4827 => x"82",
          4828 => x"82",
          4829 => x"b5",
          4830 => x"80",
          4831 => x"83",
          4832 => x"ff",
          4833 => x"82",
          4834 => x"54",
          4835 => x"74",
          4836 => x"76",
          4837 => x"82",
          4838 => x"54",
          4839 => x"34",
          4840 => x"34",
          4841 => x"08",
          4842 => x"15",
          4843 => x"15",
          4844 => x"a0",
          4845 => x"9c",
          4846 => x"fe",
          4847 => x"70",
          4848 => x"06",
          4849 => x"58",
          4850 => x"74",
          4851 => x"73",
          4852 => x"82",
          4853 => x"70",
          4854 => x"b5",
          4855 => x"f8",
          4856 => x"55",
          4857 => x"34",
          4858 => x"34",
          4859 => x"04",
          4860 => x"73",
          4861 => x"84",
          4862 => x"38",
          4863 => x"2a",
          4864 => x"83",
          4865 => x"51",
          4866 => x"82",
          4867 => x"83",
          4868 => x"f9",
          4869 => x"a6",
          4870 => x"84",
          4871 => x"22",
          4872 => x"b5",
          4873 => x"83",
          4874 => x"74",
          4875 => x"11",
          4876 => x"12",
          4877 => x"2b",
          4878 => x"05",
          4879 => x"71",
          4880 => x"06",
          4881 => x"2a",
          4882 => x"59",
          4883 => x"57",
          4884 => x"71",
          4885 => x"81",
          4886 => x"b5",
          4887 => x"75",
          4888 => x"54",
          4889 => x"34",
          4890 => x"34",
          4891 => x"08",
          4892 => x"33",
          4893 => x"71",
          4894 => x"70",
          4895 => x"ff",
          4896 => x"52",
          4897 => x"05",
          4898 => x"ff",
          4899 => x"2a",
          4900 => x"71",
          4901 => x"72",
          4902 => x"53",
          4903 => x"34",
          4904 => x"08",
          4905 => x"76",
          4906 => x"17",
          4907 => x"0d",
          4908 => x"0d",
          4909 => x"08",
          4910 => x"9e",
          4911 => x"83",
          4912 => x"86",
          4913 => x"12",
          4914 => x"2b",
          4915 => x"07",
          4916 => x"52",
          4917 => x"05",
          4918 => x"85",
          4919 => x"88",
          4920 => x"88",
          4921 => x"56",
          4922 => x"13",
          4923 => x"13",
          4924 => x"a0",
          4925 => x"84",
          4926 => x"12",
          4927 => x"2b",
          4928 => x"07",
          4929 => x"52",
          4930 => x"12",
          4931 => x"33",
          4932 => x"07",
          4933 => x"54",
          4934 => x"70",
          4935 => x"73",
          4936 => x"82",
          4937 => x"13",
          4938 => x"12",
          4939 => x"2b",
          4940 => x"ff",
          4941 => x"88",
          4942 => x"53",
          4943 => x"73",
          4944 => x"14",
          4945 => x"0d",
          4946 => x"0d",
          4947 => x"22",
          4948 => x"08",
          4949 => x"71",
          4950 => x"81",
          4951 => x"88",
          4952 => x"88",
          4953 => x"33",
          4954 => x"71",
          4955 => x"90",
          4956 => x"5f",
          4957 => x"5a",
          4958 => x"54",
          4959 => x"80",
          4960 => x"51",
          4961 => x"82",
          4962 => x"70",
          4963 => x"81",
          4964 => x"8b",
          4965 => x"2b",
          4966 => x"70",
          4967 => x"33",
          4968 => x"07",
          4969 => x"8f",
          4970 => x"51",
          4971 => x"53",
          4972 => x"72",
          4973 => x"2a",
          4974 => x"82",
          4975 => x"83",
          4976 => x"b5",
          4977 => x"16",
          4978 => x"12",
          4979 => x"2b",
          4980 => x"07",
          4981 => x"55",
          4982 => x"33",
          4983 => x"71",
          4984 => x"70",
          4985 => x"06",
          4986 => x"57",
          4987 => x"52",
          4988 => x"71",
          4989 => x"88",
          4990 => x"fb",
          4991 => x"b5",
          4992 => x"84",
          4993 => x"22",
          4994 => x"72",
          4995 => x"33",
          4996 => x"71",
          4997 => x"83",
          4998 => x"5b",
          4999 => x"52",
          5000 => x"33",
          5001 => x"71",
          5002 => x"02",
          5003 => x"05",
          5004 => x"70",
          5005 => x"51",
          5006 => x"71",
          5007 => x"81",
          5008 => x"b5",
          5009 => x"15",
          5010 => x"12",
          5011 => x"2b",
          5012 => x"07",
          5013 => x"52",
          5014 => x"12",
          5015 => x"33",
          5016 => x"07",
          5017 => x"54",
          5018 => x"70",
          5019 => x"72",
          5020 => x"82",
          5021 => x"14",
          5022 => x"83",
          5023 => x"88",
          5024 => x"b5",
          5025 => x"54",
          5026 => x"04",
          5027 => x"7b",
          5028 => x"08",
          5029 => x"70",
          5030 => x"06",
          5031 => x"53",
          5032 => x"82",
          5033 => x"76",
          5034 => x"11",
          5035 => x"83",
          5036 => x"8b",
          5037 => x"2b",
          5038 => x"70",
          5039 => x"33",
          5040 => x"71",
          5041 => x"53",
          5042 => x"53",
          5043 => x"59",
          5044 => x"25",
          5045 => x"80",
          5046 => x"51",
          5047 => x"81",
          5048 => x"14",
          5049 => x"33",
          5050 => x"71",
          5051 => x"76",
          5052 => x"2a",
          5053 => x"58",
          5054 => x"14",
          5055 => x"ff",
          5056 => x"87",
          5057 => x"b5",
          5058 => x"19",
          5059 => x"85",
          5060 => x"88",
          5061 => x"88",
          5062 => x"5b",
          5063 => x"84",
          5064 => x"85",
          5065 => x"b5",
          5066 => x"53",
          5067 => x"14",
          5068 => x"87",
          5069 => x"b5",
          5070 => x"76",
          5071 => x"75",
          5072 => x"82",
          5073 => x"18",
          5074 => x"12",
          5075 => x"2b",
          5076 => x"80",
          5077 => x"88",
          5078 => x"55",
          5079 => x"74",
          5080 => x"15",
          5081 => x"0d",
          5082 => x"0d",
          5083 => x"b5",
          5084 => x"38",
          5085 => x"71",
          5086 => x"38",
          5087 => x"8c",
          5088 => x"0d",
          5089 => x"0d",
          5090 => x"58",
          5091 => x"82",
          5092 => x"83",
          5093 => x"82",
          5094 => x"84",
          5095 => x"12",
          5096 => x"2b",
          5097 => x"59",
          5098 => x"81",
          5099 => x"75",
          5100 => x"cb",
          5101 => x"29",
          5102 => x"81",
          5103 => x"88",
          5104 => x"81",
          5105 => x"79",
          5106 => x"ff",
          5107 => x"7f",
          5108 => x"51",
          5109 => x"77",
          5110 => x"38",
          5111 => x"85",
          5112 => x"5a",
          5113 => x"33",
          5114 => x"71",
          5115 => x"57",
          5116 => x"38",
          5117 => x"ff",
          5118 => x"7a",
          5119 => x"80",
          5120 => x"82",
          5121 => x"11",
          5122 => x"12",
          5123 => x"2b",
          5124 => x"ff",
          5125 => x"52",
          5126 => x"55",
          5127 => x"83",
          5128 => x"80",
          5129 => x"26",
          5130 => x"74",
          5131 => x"2e",
          5132 => x"77",
          5133 => x"81",
          5134 => x"75",
          5135 => x"3f",
          5136 => x"82",
          5137 => x"79",
          5138 => x"f7",
          5139 => x"b5",
          5140 => x"1c",
          5141 => x"87",
          5142 => x"8b",
          5143 => x"2b",
          5144 => x"5e",
          5145 => x"7a",
          5146 => x"ff",
          5147 => x"88",
          5148 => x"56",
          5149 => x"15",
          5150 => x"ff",
          5151 => x"85",
          5152 => x"b5",
          5153 => x"83",
          5154 => x"72",
          5155 => x"33",
          5156 => x"71",
          5157 => x"70",
          5158 => x"5b",
          5159 => x"56",
          5160 => x"19",
          5161 => x"19",
          5162 => x"a0",
          5163 => x"84",
          5164 => x"12",
          5165 => x"2b",
          5166 => x"07",
          5167 => x"55",
          5168 => x"78",
          5169 => x"76",
          5170 => x"82",
          5171 => x"70",
          5172 => x"84",
          5173 => x"12",
          5174 => x"2b",
          5175 => x"2a",
          5176 => x"52",
          5177 => x"84",
          5178 => x"85",
          5179 => x"b5",
          5180 => x"84",
          5181 => x"82",
          5182 => x"8d",
          5183 => x"fe",
          5184 => x"52",
          5185 => x"08",
          5186 => x"dc",
          5187 => x"71",
          5188 => x"38",
          5189 => x"ed",
          5190 => x"a8",
          5191 => x"82",
          5192 => x"84",
          5193 => x"ee",
          5194 => x"66",
          5195 => x"70",
          5196 => x"b5",
          5197 => x"2e",
          5198 => x"84",
          5199 => x"3f",
          5200 => x"7e",
          5201 => x"3f",
          5202 => x"08",
          5203 => x"39",
          5204 => x"7b",
          5205 => x"3f",
          5206 => x"ba",
          5207 => x"f5",
          5208 => x"b5",
          5209 => x"ff",
          5210 => x"b5",
          5211 => x"71",
          5212 => x"70",
          5213 => x"06",
          5214 => x"73",
          5215 => x"81",
          5216 => x"88",
          5217 => x"75",
          5218 => x"ff",
          5219 => x"88",
          5220 => x"73",
          5221 => x"70",
          5222 => x"33",
          5223 => x"07",
          5224 => x"53",
          5225 => x"48",
          5226 => x"54",
          5227 => x"56",
          5228 => x"80",
          5229 => x"76",
          5230 => x"06",
          5231 => x"83",
          5232 => x"42",
          5233 => x"33",
          5234 => x"71",
          5235 => x"70",
          5236 => x"70",
          5237 => x"33",
          5238 => x"71",
          5239 => x"53",
          5240 => x"56",
          5241 => x"25",
          5242 => x"75",
          5243 => x"ff",
          5244 => x"54",
          5245 => x"81",
          5246 => x"18",
          5247 => x"2e",
          5248 => x"8f",
          5249 => x"f6",
          5250 => x"83",
          5251 => x"58",
          5252 => x"7f",
          5253 => x"74",
          5254 => x"78",
          5255 => x"3f",
          5256 => x"7f",
          5257 => x"75",
          5258 => x"38",
          5259 => x"11",
          5260 => x"33",
          5261 => x"07",
          5262 => x"f4",
          5263 => x"52",
          5264 => x"b7",
          5265 => x"a8",
          5266 => x"ff",
          5267 => x"7c",
          5268 => x"2b",
          5269 => x"08",
          5270 => x"53",
          5271 => x"9f",
          5272 => x"b5",
          5273 => x"84",
          5274 => x"ff",
          5275 => x"5c",
          5276 => x"60",
          5277 => x"74",
          5278 => x"38",
          5279 => x"c9",
          5280 => x"a0",
          5281 => x"11",
          5282 => x"33",
          5283 => x"07",
          5284 => x"f4",
          5285 => x"52",
          5286 => x"df",
          5287 => x"a8",
          5288 => x"ff",
          5289 => x"7c",
          5290 => x"2b",
          5291 => x"08",
          5292 => x"53",
          5293 => x"9f",
          5294 => x"b5",
          5295 => x"84",
          5296 => x"05",
          5297 => x"73",
          5298 => x"06",
          5299 => x"7b",
          5300 => x"f9",
          5301 => x"b5",
          5302 => x"82",
          5303 => x"80",
          5304 => x"7d",
          5305 => x"82",
          5306 => x"51",
          5307 => x"3f",
          5308 => x"98",
          5309 => x"7a",
          5310 => x"38",
          5311 => x"52",
          5312 => x"8f",
          5313 => x"83",
          5314 => x"a0",
          5315 => x"05",
          5316 => x"3f",
          5317 => x"82",
          5318 => x"94",
          5319 => x"fc",
          5320 => x"77",
          5321 => x"54",
          5322 => x"82",
          5323 => x"55",
          5324 => x"08",
          5325 => x"38",
          5326 => x"52",
          5327 => x"08",
          5328 => x"c2",
          5329 => x"b5",
          5330 => x"3d",
          5331 => x"3d",
          5332 => x"05",
          5333 => x"52",
          5334 => x"87",
          5335 => x"a4",
          5336 => x"71",
          5337 => x"0c",
          5338 => x"04",
          5339 => x"02",
          5340 => x"02",
          5341 => x"05",
          5342 => x"83",
          5343 => x"26",
          5344 => x"72",
          5345 => x"c0",
          5346 => x"53",
          5347 => x"74",
          5348 => x"38",
          5349 => x"73",
          5350 => x"c0",
          5351 => x"51",
          5352 => x"85",
          5353 => x"98",
          5354 => x"52",
          5355 => x"82",
          5356 => x"70",
          5357 => x"38",
          5358 => x"8c",
          5359 => x"ec",
          5360 => x"fc",
          5361 => x"52",
          5362 => x"87",
          5363 => x"08",
          5364 => x"2e",
          5365 => x"82",
          5366 => x"34",
          5367 => x"13",
          5368 => x"82",
          5369 => x"86",
          5370 => x"f3",
          5371 => x"62",
          5372 => x"05",
          5373 => x"57",
          5374 => x"83",
          5375 => x"fe",
          5376 => x"b5",
          5377 => x"06",
          5378 => x"71",
          5379 => x"71",
          5380 => x"2b",
          5381 => x"80",
          5382 => x"92",
          5383 => x"c0",
          5384 => x"41",
          5385 => x"5a",
          5386 => x"87",
          5387 => x"0c",
          5388 => x"84",
          5389 => x"08",
          5390 => x"70",
          5391 => x"53",
          5392 => x"2e",
          5393 => x"08",
          5394 => x"70",
          5395 => x"34",
          5396 => x"80",
          5397 => x"53",
          5398 => x"2e",
          5399 => x"53",
          5400 => x"26",
          5401 => x"80",
          5402 => x"87",
          5403 => x"08",
          5404 => x"38",
          5405 => x"8c",
          5406 => x"80",
          5407 => x"78",
          5408 => x"99",
          5409 => x"0c",
          5410 => x"8c",
          5411 => x"08",
          5412 => x"51",
          5413 => x"38",
          5414 => x"8d",
          5415 => x"17",
          5416 => x"81",
          5417 => x"53",
          5418 => x"2e",
          5419 => x"fc",
          5420 => x"52",
          5421 => x"7d",
          5422 => x"ed",
          5423 => x"80",
          5424 => x"71",
          5425 => x"38",
          5426 => x"53",
          5427 => x"a8",
          5428 => x"0d",
          5429 => x"0d",
          5430 => x"02",
          5431 => x"05",
          5432 => x"58",
          5433 => x"80",
          5434 => x"fc",
          5435 => x"b5",
          5436 => x"06",
          5437 => x"71",
          5438 => x"81",
          5439 => x"38",
          5440 => x"2b",
          5441 => x"80",
          5442 => x"92",
          5443 => x"c0",
          5444 => x"40",
          5445 => x"5a",
          5446 => x"c0",
          5447 => x"76",
          5448 => x"76",
          5449 => x"75",
          5450 => x"2a",
          5451 => x"51",
          5452 => x"80",
          5453 => x"7a",
          5454 => x"5c",
          5455 => x"81",
          5456 => x"81",
          5457 => x"06",
          5458 => x"80",
          5459 => x"87",
          5460 => x"08",
          5461 => x"38",
          5462 => x"8c",
          5463 => x"80",
          5464 => x"77",
          5465 => x"99",
          5466 => x"0c",
          5467 => x"8c",
          5468 => x"08",
          5469 => x"51",
          5470 => x"38",
          5471 => x"8d",
          5472 => x"70",
          5473 => x"84",
          5474 => x"5b",
          5475 => x"2e",
          5476 => x"fc",
          5477 => x"52",
          5478 => x"7d",
          5479 => x"f8",
          5480 => x"80",
          5481 => x"71",
          5482 => x"38",
          5483 => x"53",
          5484 => x"a8",
          5485 => x"0d",
          5486 => x"0d",
          5487 => x"05",
          5488 => x"02",
          5489 => x"05",
          5490 => x"54",
          5491 => x"fe",
          5492 => x"a8",
          5493 => x"53",
          5494 => x"80",
          5495 => x"0b",
          5496 => x"8c",
          5497 => x"71",
          5498 => x"dc",
          5499 => x"24",
          5500 => x"84",
          5501 => x"92",
          5502 => x"54",
          5503 => x"8d",
          5504 => x"39",
          5505 => x"80",
          5506 => x"cb",
          5507 => x"70",
          5508 => x"81",
          5509 => x"52",
          5510 => x"8a",
          5511 => x"98",
          5512 => x"71",
          5513 => x"c0",
          5514 => x"52",
          5515 => x"81",
          5516 => x"c0",
          5517 => x"53",
          5518 => x"82",
          5519 => x"71",
          5520 => x"39",
          5521 => x"39",
          5522 => x"77",
          5523 => x"81",
          5524 => x"72",
          5525 => x"84",
          5526 => x"73",
          5527 => x"0c",
          5528 => x"04",
          5529 => x"74",
          5530 => x"71",
          5531 => x"2b",
          5532 => x"a8",
          5533 => x"84",
          5534 => x"fd",
          5535 => x"83",
          5536 => x"12",
          5537 => x"2b",
          5538 => x"07",
          5539 => x"70",
          5540 => x"2b",
          5541 => x"07",
          5542 => x"0c",
          5543 => x"56",
          5544 => x"3d",
          5545 => x"3d",
          5546 => x"84",
          5547 => x"22",
          5548 => x"72",
          5549 => x"54",
          5550 => x"2a",
          5551 => x"34",
          5552 => x"04",
          5553 => x"73",
          5554 => x"70",
          5555 => x"05",
          5556 => x"88",
          5557 => x"72",
          5558 => x"54",
          5559 => x"2a",
          5560 => x"70",
          5561 => x"34",
          5562 => x"51",
          5563 => x"83",
          5564 => x"fe",
          5565 => x"75",
          5566 => x"51",
          5567 => x"92",
          5568 => x"81",
          5569 => x"73",
          5570 => x"55",
          5571 => x"51",
          5572 => x"3d",
          5573 => x"3d",
          5574 => x"76",
          5575 => x"72",
          5576 => x"05",
          5577 => x"11",
          5578 => x"38",
          5579 => x"04",
          5580 => x"78",
          5581 => x"56",
          5582 => x"81",
          5583 => x"74",
          5584 => x"56",
          5585 => x"31",
          5586 => x"52",
          5587 => x"80",
          5588 => x"71",
          5589 => x"38",
          5590 => x"a8",
          5591 => x"0d",
          5592 => x"0d",
          5593 => x"51",
          5594 => x"73",
          5595 => x"81",
          5596 => x"33",
          5597 => x"38",
          5598 => x"b5",
          5599 => x"3d",
          5600 => x"0b",
          5601 => x"0c",
          5602 => x"82",
          5603 => x"04",
          5604 => x"7b",
          5605 => x"83",
          5606 => x"5a",
          5607 => x"80",
          5608 => x"54",
          5609 => x"53",
          5610 => x"53",
          5611 => x"52",
          5612 => x"3f",
          5613 => x"08",
          5614 => x"81",
          5615 => x"82",
          5616 => x"83",
          5617 => x"16",
          5618 => x"18",
          5619 => x"18",
          5620 => x"58",
          5621 => x"9f",
          5622 => x"33",
          5623 => x"2e",
          5624 => x"93",
          5625 => x"76",
          5626 => x"52",
          5627 => x"51",
          5628 => x"83",
          5629 => x"79",
          5630 => x"0c",
          5631 => x"04",
          5632 => x"78",
          5633 => x"80",
          5634 => x"17",
          5635 => x"38",
          5636 => x"fc",
          5637 => x"a8",
          5638 => x"b5",
          5639 => x"38",
          5640 => x"53",
          5641 => x"81",
          5642 => x"f7",
          5643 => x"b5",
          5644 => x"2e",
          5645 => x"55",
          5646 => x"b0",
          5647 => x"82",
          5648 => x"88",
          5649 => x"f8",
          5650 => x"70",
          5651 => x"c0",
          5652 => x"a8",
          5653 => x"b5",
          5654 => x"91",
          5655 => x"55",
          5656 => x"09",
          5657 => x"f0",
          5658 => x"33",
          5659 => x"2e",
          5660 => x"80",
          5661 => x"80",
          5662 => x"a8",
          5663 => x"17",
          5664 => x"fd",
          5665 => x"d4",
          5666 => x"b2",
          5667 => x"96",
          5668 => x"85",
          5669 => x"75",
          5670 => x"3f",
          5671 => x"e4",
          5672 => x"98",
          5673 => x"9c",
          5674 => x"08",
          5675 => x"17",
          5676 => x"3f",
          5677 => x"52",
          5678 => x"51",
          5679 => x"a0",
          5680 => x"05",
          5681 => x"0c",
          5682 => x"75",
          5683 => x"33",
          5684 => x"3f",
          5685 => x"34",
          5686 => x"52",
          5687 => x"51",
          5688 => x"82",
          5689 => x"80",
          5690 => x"81",
          5691 => x"b5",
          5692 => x"3d",
          5693 => x"3d",
          5694 => x"1a",
          5695 => x"fe",
          5696 => x"54",
          5697 => x"73",
          5698 => x"8a",
          5699 => x"71",
          5700 => x"08",
          5701 => x"75",
          5702 => x"0c",
          5703 => x"04",
          5704 => x"7a",
          5705 => x"56",
          5706 => x"77",
          5707 => x"38",
          5708 => x"08",
          5709 => x"38",
          5710 => x"54",
          5711 => x"2e",
          5712 => x"72",
          5713 => x"38",
          5714 => x"8d",
          5715 => x"39",
          5716 => x"81",
          5717 => x"b6",
          5718 => x"2a",
          5719 => x"2a",
          5720 => x"05",
          5721 => x"55",
          5722 => x"82",
          5723 => x"81",
          5724 => x"83",
          5725 => x"b4",
          5726 => x"17",
          5727 => x"a4",
          5728 => x"55",
          5729 => x"57",
          5730 => x"3f",
          5731 => x"08",
          5732 => x"74",
          5733 => x"14",
          5734 => x"70",
          5735 => x"07",
          5736 => x"71",
          5737 => x"52",
          5738 => x"72",
          5739 => x"75",
          5740 => x"58",
          5741 => x"76",
          5742 => x"15",
          5743 => x"73",
          5744 => x"3f",
          5745 => x"08",
          5746 => x"76",
          5747 => x"06",
          5748 => x"05",
          5749 => x"3f",
          5750 => x"08",
          5751 => x"06",
          5752 => x"76",
          5753 => x"15",
          5754 => x"73",
          5755 => x"3f",
          5756 => x"08",
          5757 => x"82",
          5758 => x"06",
          5759 => x"05",
          5760 => x"3f",
          5761 => x"08",
          5762 => x"58",
          5763 => x"58",
          5764 => x"a8",
          5765 => x"0d",
          5766 => x"0d",
          5767 => x"5a",
          5768 => x"59",
          5769 => x"82",
          5770 => x"98",
          5771 => x"82",
          5772 => x"33",
          5773 => x"2e",
          5774 => x"72",
          5775 => x"38",
          5776 => x"8d",
          5777 => x"39",
          5778 => x"81",
          5779 => x"f7",
          5780 => x"2a",
          5781 => x"2a",
          5782 => x"05",
          5783 => x"55",
          5784 => x"82",
          5785 => x"59",
          5786 => x"08",
          5787 => x"74",
          5788 => x"16",
          5789 => x"16",
          5790 => x"59",
          5791 => x"53",
          5792 => x"8f",
          5793 => x"2b",
          5794 => x"74",
          5795 => x"71",
          5796 => x"72",
          5797 => x"0b",
          5798 => x"74",
          5799 => x"17",
          5800 => x"75",
          5801 => x"3f",
          5802 => x"08",
          5803 => x"a8",
          5804 => x"38",
          5805 => x"06",
          5806 => x"78",
          5807 => x"54",
          5808 => x"77",
          5809 => x"33",
          5810 => x"71",
          5811 => x"51",
          5812 => x"34",
          5813 => x"76",
          5814 => x"17",
          5815 => x"75",
          5816 => x"3f",
          5817 => x"08",
          5818 => x"a8",
          5819 => x"38",
          5820 => x"ff",
          5821 => x"10",
          5822 => x"76",
          5823 => x"51",
          5824 => x"be",
          5825 => x"2a",
          5826 => x"05",
          5827 => x"f9",
          5828 => x"b5",
          5829 => x"82",
          5830 => x"ab",
          5831 => x"0a",
          5832 => x"2b",
          5833 => x"70",
          5834 => x"70",
          5835 => x"54",
          5836 => x"82",
          5837 => x"8f",
          5838 => x"07",
          5839 => x"f7",
          5840 => x"0b",
          5841 => x"78",
          5842 => x"0c",
          5843 => x"04",
          5844 => x"7a",
          5845 => x"08",
          5846 => x"59",
          5847 => x"a4",
          5848 => x"17",
          5849 => x"38",
          5850 => x"aa",
          5851 => x"73",
          5852 => x"fd",
          5853 => x"b5",
          5854 => x"82",
          5855 => x"80",
          5856 => x"39",
          5857 => x"eb",
          5858 => x"80",
          5859 => x"b5",
          5860 => x"80",
          5861 => x"52",
          5862 => x"84",
          5863 => x"a8",
          5864 => x"b5",
          5865 => x"2e",
          5866 => x"82",
          5867 => x"81",
          5868 => x"82",
          5869 => x"ff",
          5870 => x"80",
          5871 => x"75",
          5872 => x"3f",
          5873 => x"08",
          5874 => x"16",
          5875 => x"90",
          5876 => x"55",
          5877 => x"27",
          5878 => x"15",
          5879 => x"84",
          5880 => x"07",
          5881 => x"17",
          5882 => x"76",
          5883 => x"a6",
          5884 => x"73",
          5885 => x"0c",
          5886 => x"04",
          5887 => x"7c",
          5888 => x"59",
          5889 => x"95",
          5890 => x"08",
          5891 => x"2e",
          5892 => x"17",
          5893 => x"b2",
          5894 => x"ae",
          5895 => x"7a",
          5896 => x"3f",
          5897 => x"82",
          5898 => x"27",
          5899 => x"82",
          5900 => x"55",
          5901 => x"08",
          5902 => x"d2",
          5903 => x"08",
          5904 => x"08",
          5905 => x"38",
          5906 => x"17",
          5907 => x"54",
          5908 => x"82",
          5909 => x"7a",
          5910 => x"06",
          5911 => x"81",
          5912 => x"17",
          5913 => x"83",
          5914 => x"75",
          5915 => x"f9",
          5916 => x"59",
          5917 => x"08",
          5918 => x"81",
          5919 => x"82",
          5920 => x"59",
          5921 => x"08",
          5922 => x"70",
          5923 => x"25",
          5924 => x"82",
          5925 => x"54",
          5926 => x"55",
          5927 => x"38",
          5928 => x"08",
          5929 => x"38",
          5930 => x"54",
          5931 => x"90",
          5932 => x"18",
          5933 => x"38",
          5934 => x"39",
          5935 => x"38",
          5936 => x"16",
          5937 => x"08",
          5938 => x"38",
          5939 => x"78",
          5940 => x"38",
          5941 => x"51",
          5942 => x"82",
          5943 => x"80",
          5944 => x"80",
          5945 => x"a8",
          5946 => x"09",
          5947 => x"38",
          5948 => x"08",
          5949 => x"a8",
          5950 => x"30",
          5951 => x"80",
          5952 => x"07",
          5953 => x"55",
          5954 => x"38",
          5955 => x"09",
          5956 => x"ae",
          5957 => x"80",
          5958 => x"53",
          5959 => x"51",
          5960 => x"82",
          5961 => x"82",
          5962 => x"30",
          5963 => x"a8",
          5964 => x"25",
          5965 => x"79",
          5966 => x"38",
          5967 => x"8f",
          5968 => x"79",
          5969 => x"f9",
          5970 => x"b5",
          5971 => x"74",
          5972 => x"8c",
          5973 => x"17",
          5974 => x"90",
          5975 => x"54",
          5976 => x"86",
          5977 => x"90",
          5978 => x"17",
          5979 => x"54",
          5980 => x"34",
          5981 => x"56",
          5982 => x"90",
          5983 => x"80",
          5984 => x"82",
          5985 => x"55",
          5986 => x"56",
          5987 => x"82",
          5988 => x"8c",
          5989 => x"f8",
          5990 => x"70",
          5991 => x"f0",
          5992 => x"a8",
          5993 => x"56",
          5994 => x"08",
          5995 => x"7b",
          5996 => x"f6",
          5997 => x"b5",
          5998 => x"b5",
          5999 => x"17",
          6000 => x"80",
          6001 => x"b4",
          6002 => x"57",
          6003 => x"77",
          6004 => x"81",
          6005 => x"15",
          6006 => x"78",
          6007 => x"81",
          6008 => x"53",
          6009 => x"15",
          6010 => x"e9",
          6011 => x"a8",
          6012 => x"df",
          6013 => x"22",
          6014 => x"30",
          6015 => x"70",
          6016 => x"51",
          6017 => x"82",
          6018 => x"8a",
          6019 => x"f8",
          6020 => x"7c",
          6021 => x"56",
          6022 => x"80",
          6023 => x"f1",
          6024 => x"06",
          6025 => x"e9",
          6026 => x"18",
          6027 => x"08",
          6028 => x"38",
          6029 => x"82",
          6030 => x"38",
          6031 => x"54",
          6032 => x"74",
          6033 => x"82",
          6034 => x"22",
          6035 => x"79",
          6036 => x"38",
          6037 => x"98",
          6038 => x"cd",
          6039 => x"22",
          6040 => x"54",
          6041 => x"26",
          6042 => x"52",
          6043 => x"b0",
          6044 => x"a8",
          6045 => x"b5",
          6046 => x"2e",
          6047 => x"0b",
          6048 => x"08",
          6049 => x"98",
          6050 => x"b5",
          6051 => x"85",
          6052 => x"bd",
          6053 => x"31",
          6054 => x"73",
          6055 => x"f4",
          6056 => x"b5",
          6057 => x"18",
          6058 => x"18",
          6059 => x"08",
          6060 => x"72",
          6061 => x"38",
          6062 => x"58",
          6063 => x"89",
          6064 => x"18",
          6065 => x"ff",
          6066 => x"05",
          6067 => x"80",
          6068 => x"b5",
          6069 => x"3d",
          6070 => x"3d",
          6071 => x"08",
          6072 => x"a0",
          6073 => x"54",
          6074 => x"77",
          6075 => x"80",
          6076 => x"0c",
          6077 => x"53",
          6078 => x"80",
          6079 => x"38",
          6080 => x"06",
          6081 => x"b5",
          6082 => x"98",
          6083 => x"14",
          6084 => x"92",
          6085 => x"2a",
          6086 => x"56",
          6087 => x"26",
          6088 => x"80",
          6089 => x"16",
          6090 => x"77",
          6091 => x"53",
          6092 => x"38",
          6093 => x"51",
          6094 => x"82",
          6095 => x"53",
          6096 => x"0b",
          6097 => x"08",
          6098 => x"38",
          6099 => x"b5",
          6100 => x"2e",
          6101 => x"98",
          6102 => x"b5",
          6103 => x"80",
          6104 => x"8a",
          6105 => x"15",
          6106 => x"80",
          6107 => x"14",
          6108 => x"51",
          6109 => x"82",
          6110 => x"53",
          6111 => x"b5",
          6112 => x"2e",
          6113 => x"82",
          6114 => x"a8",
          6115 => x"ba",
          6116 => x"82",
          6117 => x"ff",
          6118 => x"82",
          6119 => x"52",
          6120 => x"f3",
          6121 => x"a8",
          6122 => x"72",
          6123 => x"72",
          6124 => x"f2",
          6125 => x"b5",
          6126 => x"15",
          6127 => x"15",
          6128 => x"b4",
          6129 => x"0c",
          6130 => x"82",
          6131 => x"8a",
          6132 => x"f7",
          6133 => x"7d",
          6134 => x"5b",
          6135 => x"76",
          6136 => x"3f",
          6137 => x"08",
          6138 => x"a8",
          6139 => x"38",
          6140 => x"08",
          6141 => x"08",
          6142 => x"f0",
          6143 => x"b5",
          6144 => x"82",
          6145 => x"80",
          6146 => x"b5",
          6147 => x"18",
          6148 => x"51",
          6149 => x"81",
          6150 => x"81",
          6151 => x"81",
          6152 => x"a8",
          6153 => x"83",
          6154 => x"77",
          6155 => x"72",
          6156 => x"38",
          6157 => x"75",
          6158 => x"81",
          6159 => x"a5",
          6160 => x"a8",
          6161 => x"52",
          6162 => x"8e",
          6163 => x"a8",
          6164 => x"b5",
          6165 => x"2e",
          6166 => x"73",
          6167 => x"81",
          6168 => x"87",
          6169 => x"b5",
          6170 => x"3d",
          6171 => x"3d",
          6172 => x"11",
          6173 => x"ec",
          6174 => x"a8",
          6175 => x"ff",
          6176 => x"33",
          6177 => x"71",
          6178 => x"81",
          6179 => x"94",
          6180 => x"d0",
          6181 => x"a8",
          6182 => x"73",
          6183 => x"82",
          6184 => x"85",
          6185 => x"fc",
          6186 => x"79",
          6187 => x"ff",
          6188 => x"12",
          6189 => x"eb",
          6190 => x"70",
          6191 => x"72",
          6192 => x"81",
          6193 => x"73",
          6194 => x"94",
          6195 => x"d6",
          6196 => x"0d",
          6197 => x"0d",
          6198 => x"55",
          6199 => x"5a",
          6200 => x"08",
          6201 => x"8a",
          6202 => x"08",
          6203 => x"ee",
          6204 => x"b5",
          6205 => x"82",
          6206 => x"80",
          6207 => x"15",
          6208 => x"55",
          6209 => x"38",
          6210 => x"e6",
          6211 => x"33",
          6212 => x"70",
          6213 => x"58",
          6214 => x"86",
          6215 => x"b5",
          6216 => x"73",
          6217 => x"83",
          6218 => x"73",
          6219 => x"38",
          6220 => x"06",
          6221 => x"80",
          6222 => x"75",
          6223 => x"38",
          6224 => x"08",
          6225 => x"54",
          6226 => x"2e",
          6227 => x"83",
          6228 => x"73",
          6229 => x"38",
          6230 => x"51",
          6231 => x"82",
          6232 => x"58",
          6233 => x"08",
          6234 => x"15",
          6235 => x"38",
          6236 => x"0b",
          6237 => x"77",
          6238 => x"0c",
          6239 => x"04",
          6240 => x"77",
          6241 => x"54",
          6242 => x"51",
          6243 => x"82",
          6244 => x"55",
          6245 => x"08",
          6246 => x"14",
          6247 => x"51",
          6248 => x"82",
          6249 => x"55",
          6250 => x"08",
          6251 => x"53",
          6252 => x"08",
          6253 => x"08",
          6254 => x"3f",
          6255 => x"14",
          6256 => x"08",
          6257 => x"3f",
          6258 => x"17",
          6259 => x"b5",
          6260 => x"3d",
          6261 => x"3d",
          6262 => x"08",
          6263 => x"54",
          6264 => x"53",
          6265 => x"82",
          6266 => x"8d",
          6267 => x"08",
          6268 => x"34",
          6269 => x"15",
          6270 => x"0d",
          6271 => x"0d",
          6272 => x"57",
          6273 => x"17",
          6274 => x"08",
          6275 => x"82",
          6276 => x"89",
          6277 => x"55",
          6278 => x"14",
          6279 => x"16",
          6280 => x"71",
          6281 => x"38",
          6282 => x"09",
          6283 => x"38",
          6284 => x"73",
          6285 => x"81",
          6286 => x"ae",
          6287 => x"05",
          6288 => x"15",
          6289 => x"70",
          6290 => x"34",
          6291 => x"8a",
          6292 => x"38",
          6293 => x"05",
          6294 => x"81",
          6295 => x"17",
          6296 => x"12",
          6297 => x"34",
          6298 => x"9c",
          6299 => x"e8",
          6300 => x"b5",
          6301 => x"0c",
          6302 => x"e7",
          6303 => x"b5",
          6304 => x"17",
          6305 => x"51",
          6306 => x"82",
          6307 => x"84",
          6308 => x"3d",
          6309 => x"3d",
          6310 => x"08",
          6311 => x"61",
          6312 => x"55",
          6313 => x"2e",
          6314 => x"55",
          6315 => x"2e",
          6316 => x"80",
          6317 => x"94",
          6318 => x"1c",
          6319 => x"81",
          6320 => x"61",
          6321 => x"56",
          6322 => x"2e",
          6323 => x"83",
          6324 => x"73",
          6325 => x"70",
          6326 => x"25",
          6327 => x"51",
          6328 => x"38",
          6329 => x"0c",
          6330 => x"51",
          6331 => x"26",
          6332 => x"80",
          6333 => x"34",
          6334 => x"51",
          6335 => x"82",
          6336 => x"55",
          6337 => x"91",
          6338 => x"1d",
          6339 => x"8b",
          6340 => x"79",
          6341 => x"3f",
          6342 => x"57",
          6343 => x"55",
          6344 => x"2e",
          6345 => x"80",
          6346 => x"18",
          6347 => x"1a",
          6348 => x"70",
          6349 => x"2a",
          6350 => x"07",
          6351 => x"5a",
          6352 => x"8c",
          6353 => x"54",
          6354 => x"81",
          6355 => x"39",
          6356 => x"70",
          6357 => x"2a",
          6358 => x"75",
          6359 => x"8c",
          6360 => x"2e",
          6361 => x"a0",
          6362 => x"38",
          6363 => x"0c",
          6364 => x"76",
          6365 => x"38",
          6366 => x"b8",
          6367 => x"70",
          6368 => x"5a",
          6369 => x"76",
          6370 => x"38",
          6371 => x"70",
          6372 => x"dc",
          6373 => x"72",
          6374 => x"80",
          6375 => x"51",
          6376 => x"73",
          6377 => x"38",
          6378 => x"18",
          6379 => x"1a",
          6380 => x"55",
          6381 => x"2e",
          6382 => x"83",
          6383 => x"73",
          6384 => x"70",
          6385 => x"25",
          6386 => x"51",
          6387 => x"38",
          6388 => x"75",
          6389 => x"81",
          6390 => x"81",
          6391 => x"27",
          6392 => x"73",
          6393 => x"38",
          6394 => x"70",
          6395 => x"32",
          6396 => x"80",
          6397 => x"2a",
          6398 => x"56",
          6399 => x"81",
          6400 => x"57",
          6401 => x"f5",
          6402 => x"2b",
          6403 => x"25",
          6404 => x"80",
          6405 => x"ae",
          6406 => x"57",
          6407 => x"e6",
          6408 => x"b5",
          6409 => x"2e",
          6410 => x"18",
          6411 => x"1a",
          6412 => x"56",
          6413 => x"3f",
          6414 => x"08",
          6415 => x"e8",
          6416 => x"54",
          6417 => x"80",
          6418 => x"17",
          6419 => x"34",
          6420 => x"11",
          6421 => x"74",
          6422 => x"75",
          6423 => x"90",
          6424 => x"3f",
          6425 => x"08",
          6426 => x"9f",
          6427 => x"99",
          6428 => x"e0",
          6429 => x"ff",
          6430 => x"79",
          6431 => x"74",
          6432 => x"57",
          6433 => x"77",
          6434 => x"76",
          6435 => x"38",
          6436 => x"73",
          6437 => x"09",
          6438 => x"38",
          6439 => x"84",
          6440 => x"27",
          6441 => x"39",
          6442 => x"f2",
          6443 => x"80",
          6444 => x"54",
          6445 => x"34",
          6446 => x"58",
          6447 => x"f2",
          6448 => x"b5",
          6449 => x"82",
          6450 => x"80",
          6451 => x"1b",
          6452 => x"51",
          6453 => x"82",
          6454 => x"56",
          6455 => x"08",
          6456 => x"9c",
          6457 => x"33",
          6458 => x"80",
          6459 => x"38",
          6460 => x"bf",
          6461 => x"86",
          6462 => x"15",
          6463 => x"2a",
          6464 => x"51",
          6465 => x"92",
          6466 => x"79",
          6467 => x"e4",
          6468 => x"b5",
          6469 => x"2e",
          6470 => x"52",
          6471 => x"ba",
          6472 => x"39",
          6473 => x"33",
          6474 => x"80",
          6475 => x"74",
          6476 => x"81",
          6477 => x"38",
          6478 => x"70",
          6479 => x"82",
          6480 => x"54",
          6481 => x"96",
          6482 => x"06",
          6483 => x"2e",
          6484 => x"ff",
          6485 => x"1c",
          6486 => x"80",
          6487 => x"81",
          6488 => x"ba",
          6489 => x"b6",
          6490 => x"2a",
          6491 => x"51",
          6492 => x"38",
          6493 => x"70",
          6494 => x"81",
          6495 => x"55",
          6496 => x"e1",
          6497 => x"08",
          6498 => x"1d",
          6499 => x"7c",
          6500 => x"3f",
          6501 => x"08",
          6502 => x"fa",
          6503 => x"82",
          6504 => x"8f",
          6505 => x"f6",
          6506 => x"5b",
          6507 => x"70",
          6508 => x"59",
          6509 => x"73",
          6510 => x"c6",
          6511 => x"81",
          6512 => x"70",
          6513 => x"52",
          6514 => x"8d",
          6515 => x"38",
          6516 => x"09",
          6517 => x"a5",
          6518 => x"d0",
          6519 => x"ff",
          6520 => x"53",
          6521 => x"91",
          6522 => x"73",
          6523 => x"d0",
          6524 => x"71",
          6525 => x"f7",
          6526 => x"82",
          6527 => x"55",
          6528 => x"55",
          6529 => x"81",
          6530 => x"74",
          6531 => x"56",
          6532 => x"12",
          6533 => x"70",
          6534 => x"38",
          6535 => x"81",
          6536 => x"51",
          6537 => x"51",
          6538 => x"89",
          6539 => x"70",
          6540 => x"53",
          6541 => x"70",
          6542 => x"51",
          6543 => x"09",
          6544 => x"38",
          6545 => x"38",
          6546 => x"77",
          6547 => x"70",
          6548 => x"2a",
          6549 => x"07",
          6550 => x"51",
          6551 => x"8f",
          6552 => x"84",
          6553 => x"83",
          6554 => x"94",
          6555 => x"74",
          6556 => x"38",
          6557 => x"0c",
          6558 => x"86",
          6559 => x"f4",
          6560 => x"82",
          6561 => x"8c",
          6562 => x"fa",
          6563 => x"56",
          6564 => x"17",
          6565 => x"b0",
          6566 => x"52",
          6567 => x"e0",
          6568 => x"82",
          6569 => x"81",
          6570 => x"b2",
          6571 => x"b4",
          6572 => x"a8",
          6573 => x"ff",
          6574 => x"55",
          6575 => x"d5",
          6576 => x"06",
          6577 => x"80",
          6578 => x"33",
          6579 => x"81",
          6580 => x"81",
          6581 => x"81",
          6582 => x"eb",
          6583 => x"70",
          6584 => x"07",
          6585 => x"73",
          6586 => x"81",
          6587 => x"81",
          6588 => x"83",
          6589 => x"a0",
          6590 => x"16",
          6591 => x"3f",
          6592 => x"08",
          6593 => x"a8",
          6594 => x"9d",
          6595 => x"82",
          6596 => x"81",
          6597 => x"e0",
          6598 => x"b5",
          6599 => x"82",
          6600 => x"80",
          6601 => x"82",
          6602 => x"b5",
          6603 => x"3d",
          6604 => x"3d",
          6605 => x"84",
          6606 => x"05",
          6607 => x"80",
          6608 => x"51",
          6609 => x"82",
          6610 => x"58",
          6611 => x"0b",
          6612 => x"08",
          6613 => x"38",
          6614 => x"08",
          6615 => x"cc",
          6616 => x"08",
          6617 => x"56",
          6618 => x"86",
          6619 => x"75",
          6620 => x"fe",
          6621 => x"54",
          6622 => x"2e",
          6623 => x"14",
          6624 => x"ca",
          6625 => x"a8",
          6626 => x"06",
          6627 => x"54",
          6628 => x"38",
          6629 => x"86",
          6630 => x"82",
          6631 => x"06",
          6632 => x"56",
          6633 => x"38",
          6634 => x"80",
          6635 => x"81",
          6636 => x"52",
          6637 => x"51",
          6638 => x"82",
          6639 => x"81",
          6640 => x"81",
          6641 => x"83",
          6642 => x"87",
          6643 => x"2e",
          6644 => x"82",
          6645 => x"06",
          6646 => x"56",
          6647 => x"38",
          6648 => x"74",
          6649 => x"a3",
          6650 => x"a8",
          6651 => x"06",
          6652 => x"2e",
          6653 => x"80",
          6654 => x"3d",
          6655 => x"83",
          6656 => x"15",
          6657 => x"53",
          6658 => x"8d",
          6659 => x"15",
          6660 => x"3f",
          6661 => x"08",
          6662 => x"70",
          6663 => x"0c",
          6664 => x"16",
          6665 => x"80",
          6666 => x"80",
          6667 => x"54",
          6668 => x"84",
          6669 => x"5b",
          6670 => x"80",
          6671 => x"7a",
          6672 => x"fc",
          6673 => x"b5",
          6674 => x"ff",
          6675 => x"77",
          6676 => x"81",
          6677 => x"76",
          6678 => x"81",
          6679 => x"2e",
          6680 => x"8d",
          6681 => x"26",
          6682 => x"bf",
          6683 => x"f4",
          6684 => x"a8",
          6685 => x"ff",
          6686 => x"84",
          6687 => x"81",
          6688 => x"38",
          6689 => x"51",
          6690 => x"82",
          6691 => x"83",
          6692 => x"58",
          6693 => x"80",
          6694 => x"db",
          6695 => x"b5",
          6696 => x"77",
          6697 => x"80",
          6698 => x"82",
          6699 => x"c4",
          6700 => x"11",
          6701 => x"06",
          6702 => x"8d",
          6703 => x"26",
          6704 => x"74",
          6705 => x"78",
          6706 => x"c1",
          6707 => x"59",
          6708 => x"15",
          6709 => x"2e",
          6710 => x"13",
          6711 => x"72",
          6712 => x"38",
          6713 => x"eb",
          6714 => x"14",
          6715 => x"3f",
          6716 => x"08",
          6717 => x"a8",
          6718 => x"23",
          6719 => x"57",
          6720 => x"83",
          6721 => x"c7",
          6722 => x"d8",
          6723 => x"a8",
          6724 => x"ff",
          6725 => x"8d",
          6726 => x"14",
          6727 => x"3f",
          6728 => x"08",
          6729 => x"14",
          6730 => x"3f",
          6731 => x"08",
          6732 => x"06",
          6733 => x"72",
          6734 => x"97",
          6735 => x"22",
          6736 => x"84",
          6737 => x"5a",
          6738 => x"83",
          6739 => x"14",
          6740 => x"79",
          6741 => x"ff",
          6742 => x"b5",
          6743 => x"82",
          6744 => x"80",
          6745 => x"38",
          6746 => x"08",
          6747 => x"ff",
          6748 => x"38",
          6749 => x"83",
          6750 => x"83",
          6751 => x"74",
          6752 => x"85",
          6753 => x"89",
          6754 => x"76",
          6755 => x"c3",
          6756 => x"70",
          6757 => x"7b",
          6758 => x"73",
          6759 => x"17",
          6760 => x"ac",
          6761 => x"55",
          6762 => x"09",
          6763 => x"38",
          6764 => x"51",
          6765 => x"82",
          6766 => x"83",
          6767 => x"53",
          6768 => x"82",
          6769 => x"82",
          6770 => x"e0",
          6771 => x"ab",
          6772 => x"a8",
          6773 => x"0c",
          6774 => x"53",
          6775 => x"56",
          6776 => x"81",
          6777 => x"13",
          6778 => x"74",
          6779 => x"82",
          6780 => x"74",
          6781 => x"81",
          6782 => x"06",
          6783 => x"83",
          6784 => x"2a",
          6785 => x"72",
          6786 => x"26",
          6787 => x"ff",
          6788 => x"0c",
          6789 => x"15",
          6790 => x"0b",
          6791 => x"76",
          6792 => x"81",
          6793 => x"38",
          6794 => x"51",
          6795 => x"82",
          6796 => x"83",
          6797 => x"53",
          6798 => x"09",
          6799 => x"f9",
          6800 => x"52",
          6801 => x"b8",
          6802 => x"a8",
          6803 => x"38",
          6804 => x"08",
          6805 => x"84",
          6806 => x"d8",
          6807 => x"b5",
          6808 => x"ff",
          6809 => x"72",
          6810 => x"2e",
          6811 => x"80",
          6812 => x"14",
          6813 => x"3f",
          6814 => x"08",
          6815 => x"a4",
          6816 => x"81",
          6817 => x"84",
          6818 => x"d7",
          6819 => x"b5",
          6820 => x"8a",
          6821 => x"2e",
          6822 => x"9d",
          6823 => x"14",
          6824 => x"3f",
          6825 => x"08",
          6826 => x"84",
          6827 => x"d7",
          6828 => x"b5",
          6829 => x"15",
          6830 => x"34",
          6831 => x"22",
          6832 => x"72",
          6833 => x"23",
          6834 => x"23",
          6835 => x"15",
          6836 => x"75",
          6837 => x"0c",
          6838 => x"04",
          6839 => x"77",
          6840 => x"73",
          6841 => x"38",
          6842 => x"72",
          6843 => x"38",
          6844 => x"71",
          6845 => x"38",
          6846 => x"84",
          6847 => x"52",
          6848 => x"09",
          6849 => x"38",
          6850 => x"51",
          6851 => x"82",
          6852 => x"81",
          6853 => x"88",
          6854 => x"08",
          6855 => x"39",
          6856 => x"73",
          6857 => x"74",
          6858 => x"0c",
          6859 => x"04",
          6860 => x"02",
          6861 => x"7a",
          6862 => x"fc",
          6863 => x"f4",
          6864 => x"54",
          6865 => x"b5",
          6866 => x"bc",
          6867 => x"a8",
          6868 => x"82",
          6869 => x"70",
          6870 => x"73",
          6871 => x"38",
          6872 => x"78",
          6873 => x"2e",
          6874 => x"74",
          6875 => x"0c",
          6876 => x"80",
          6877 => x"80",
          6878 => x"70",
          6879 => x"51",
          6880 => x"82",
          6881 => x"54",
          6882 => x"a8",
          6883 => x"0d",
          6884 => x"0d",
          6885 => x"05",
          6886 => x"33",
          6887 => x"54",
          6888 => x"84",
          6889 => x"bf",
          6890 => x"98",
          6891 => x"53",
          6892 => x"05",
          6893 => x"fa",
          6894 => x"a8",
          6895 => x"b5",
          6896 => x"a4",
          6897 => x"68",
          6898 => x"70",
          6899 => x"c6",
          6900 => x"a8",
          6901 => x"b5",
          6902 => x"38",
          6903 => x"05",
          6904 => x"2b",
          6905 => x"80",
          6906 => x"86",
          6907 => x"06",
          6908 => x"2e",
          6909 => x"74",
          6910 => x"38",
          6911 => x"09",
          6912 => x"38",
          6913 => x"f8",
          6914 => x"a8",
          6915 => x"39",
          6916 => x"33",
          6917 => x"73",
          6918 => x"77",
          6919 => x"81",
          6920 => x"73",
          6921 => x"38",
          6922 => x"bc",
          6923 => x"07",
          6924 => x"b4",
          6925 => x"2a",
          6926 => x"51",
          6927 => x"2e",
          6928 => x"62",
          6929 => x"e8",
          6930 => x"b5",
          6931 => x"82",
          6932 => x"52",
          6933 => x"51",
          6934 => x"62",
          6935 => x"8b",
          6936 => x"53",
          6937 => x"51",
          6938 => x"80",
          6939 => x"05",
          6940 => x"3f",
          6941 => x"0b",
          6942 => x"75",
          6943 => x"f1",
          6944 => x"11",
          6945 => x"80",
          6946 => x"97",
          6947 => x"51",
          6948 => x"82",
          6949 => x"55",
          6950 => x"08",
          6951 => x"b7",
          6952 => x"c4",
          6953 => x"05",
          6954 => x"2a",
          6955 => x"51",
          6956 => x"80",
          6957 => x"84",
          6958 => x"39",
          6959 => x"70",
          6960 => x"54",
          6961 => x"a9",
          6962 => x"06",
          6963 => x"2e",
          6964 => x"55",
          6965 => x"73",
          6966 => x"d6",
          6967 => x"b5",
          6968 => x"ff",
          6969 => x"0c",
          6970 => x"b5",
          6971 => x"f8",
          6972 => x"2a",
          6973 => x"51",
          6974 => x"2e",
          6975 => x"80",
          6976 => x"7a",
          6977 => x"a0",
          6978 => x"a4",
          6979 => x"53",
          6980 => x"e6",
          6981 => x"b5",
          6982 => x"b5",
          6983 => x"1b",
          6984 => x"05",
          6985 => x"d3",
          6986 => x"a8",
          6987 => x"a8",
          6988 => x"0c",
          6989 => x"56",
          6990 => x"84",
          6991 => x"90",
          6992 => x"0b",
          6993 => x"80",
          6994 => x"0c",
          6995 => x"1a",
          6996 => x"2a",
          6997 => x"51",
          6998 => x"2e",
          6999 => x"82",
          7000 => x"80",
          7001 => x"38",
          7002 => x"08",
          7003 => x"8a",
          7004 => x"89",
          7005 => x"59",
          7006 => x"76",
          7007 => x"d7",
          7008 => x"b5",
          7009 => x"82",
          7010 => x"81",
          7011 => x"82",
          7012 => x"a8",
          7013 => x"09",
          7014 => x"38",
          7015 => x"78",
          7016 => x"30",
          7017 => x"80",
          7018 => x"77",
          7019 => x"38",
          7020 => x"06",
          7021 => x"c3",
          7022 => x"1a",
          7023 => x"38",
          7024 => x"06",
          7025 => x"2e",
          7026 => x"52",
          7027 => x"a6",
          7028 => x"a8",
          7029 => x"82",
          7030 => x"75",
          7031 => x"b5",
          7032 => x"9c",
          7033 => x"39",
          7034 => x"74",
          7035 => x"b5",
          7036 => x"3d",
          7037 => x"3d",
          7038 => x"65",
          7039 => x"5d",
          7040 => x"0c",
          7041 => x"05",
          7042 => x"f9",
          7043 => x"b5",
          7044 => x"82",
          7045 => x"8a",
          7046 => x"33",
          7047 => x"2e",
          7048 => x"56",
          7049 => x"90",
          7050 => x"06",
          7051 => x"74",
          7052 => x"b6",
          7053 => x"82",
          7054 => x"34",
          7055 => x"aa",
          7056 => x"91",
          7057 => x"56",
          7058 => x"8c",
          7059 => x"1a",
          7060 => x"74",
          7061 => x"38",
          7062 => x"80",
          7063 => x"38",
          7064 => x"70",
          7065 => x"56",
          7066 => x"b2",
          7067 => x"11",
          7068 => x"77",
          7069 => x"5b",
          7070 => x"38",
          7071 => x"88",
          7072 => x"8f",
          7073 => x"08",
          7074 => x"d5",
          7075 => x"b5",
          7076 => x"81",
          7077 => x"9f",
          7078 => x"2e",
          7079 => x"74",
          7080 => x"98",
          7081 => x"7e",
          7082 => x"3f",
          7083 => x"08",
          7084 => x"83",
          7085 => x"a8",
          7086 => x"89",
          7087 => x"77",
          7088 => x"d6",
          7089 => x"7f",
          7090 => x"58",
          7091 => x"75",
          7092 => x"75",
          7093 => x"77",
          7094 => x"7c",
          7095 => x"33",
          7096 => x"3f",
          7097 => x"08",
          7098 => x"7e",
          7099 => x"56",
          7100 => x"2e",
          7101 => x"16",
          7102 => x"55",
          7103 => x"94",
          7104 => x"53",
          7105 => x"b0",
          7106 => x"31",
          7107 => x"05",
          7108 => x"3f",
          7109 => x"56",
          7110 => x"9c",
          7111 => x"19",
          7112 => x"06",
          7113 => x"31",
          7114 => x"76",
          7115 => x"7b",
          7116 => x"08",
          7117 => x"d1",
          7118 => x"b5",
          7119 => x"81",
          7120 => x"94",
          7121 => x"ff",
          7122 => x"05",
          7123 => x"cf",
          7124 => x"76",
          7125 => x"17",
          7126 => x"1e",
          7127 => x"18",
          7128 => x"5e",
          7129 => x"39",
          7130 => x"82",
          7131 => x"90",
          7132 => x"f2",
          7133 => x"63",
          7134 => x"40",
          7135 => x"7e",
          7136 => x"fc",
          7137 => x"51",
          7138 => x"82",
          7139 => x"55",
          7140 => x"08",
          7141 => x"18",
          7142 => x"80",
          7143 => x"74",
          7144 => x"39",
          7145 => x"70",
          7146 => x"81",
          7147 => x"56",
          7148 => x"80",
          7149 => x"38",
          7150 => x"0b",
          7151 => x"82",
          7152 => x"39",
          7153 => x"19",
          7154 => x"83",
          7155 => x"18",
          7156 => x"56",
          7157 => x"27",
          7158 => x"09",
          7159 => x"2e",
          7160 => x"94",
          7161 => x"83",
          7162 => x"56",
          7163 => x"38",
          7164 => x"22",
          7165 => x"89",
          7166 => x"55",
          7167 => x"75",
          7168 => x"18",
          7169 => x"9c",
          7170 => x"85",
          7171 => x"08",
          7172 => x"d7",
          7173 => x"b5",
          7174 => x"82",
          7175 => x"80",
          7176 => x"38",
          7177 => x"ff",
          7178 => x"ff",
          7179 => x"38",
          7180 => x"0c",
          7181 => x"85",
          7182 => x"19",
          7183 => x"b0",
          7184 => x"19",
          7185 => x"81",
          7186 => x"74",
          7187 => x"3f",
          7188 => x"08",
          7189 => x"98",
          7190 => x"7e",
          7191 => x"3f",
          7192 => x"08",
          7193 => x"d2",
          7194 => x"a8",
          7195 => x"89",
          7196 => x"78",
          7197 => x"d5",
          7198 => x"7f",
          7199 => x"58",
          7200 => x"75",
          7201 => x"75",
          7202 => x"78",
          7203 => x"7c",
          7204 => x"33",
          7205 => x"3f",
          7206 => x"08",
          7207 => x"7e",
          7208 => x"78",
          7209 => x"74",
          7210 => x"38",
          7211 => x"b0",
          7212 => x"31",
          7213 => x"05",
          7214 => x"51",
          7215 => x"7e",
          7216 => x"83",
          7217 => x"89",
          7218 => x"db",
          7219 => x"08",
          7220 => x"26",
          7221 => x"51",
          7222 => x"82",
          7223 => x"fd",
          7224 => x"77",
          7225 => x"55",
          7226 => x"0c",
          7227 => x"83",
          7228 => x"80",
          7229 => x"55",
          7230 => x"83",
          7231 => x"9c",
          7232 => x"7e",
          7233 => x"3f",
          7234 => x"08",
          7235 => x"75",
          7236 => x"94",
          7237 => x"ff",
          7238 => x"05",
          7239 => x"3f",
          7240 => x"0b",
          7241 => x"7b",
          7242 => x"08",
          7243 => x"76",
          7244 => x"08",
          7245 => x"1c",
          7246 => x"08",
          7247 => x"5c",
          7248 => x"83",
          7249 => x"74",
          7250 => x"fd",
          7251 => x"18",
          7252 => x"07",
          7253 => x"19",
          7254 => x"75",
          7255 => x"0c",
          7256 => x"04",
          7257 => x"7a",
          7258 => x"05",
          7259 => x"56",
          7260 => x"82",
          7261 => x"57",
          7262 => x"08",
          7263 => x"90",
          7264 => x"86",
          7265 => x"06",
          7266 => x"73",
          7267 => x"e9",
          7268 => x"08",
          7269 => x"cc",
          7270 => x"b5",
          7271 => x"82",
          7272 => x"80",
          7273 => x"16",
          7274 => x"33",
          7275 => x"55",
          7276 => x"34",
          7277 => x"53",
          7278 => x"08",
          7279 => x"3f",
          7280 => x"52",
          7281 => x"c9",
          7282 => x"88",
          7283 => x"96",
          7284 => x"f0",
          7285 => x"92",
          7286 => x"ca",
          7287 => x"81",
          7288 => x"34",
          7289 => x"df",
          7290 => x"a8",
          7291 => x"33",
          7292 => x"55",
          7293 => x"17",
          7294 => x"b5",
          7295 => x"3d",
          7296 => x"3d",
          7297 => x"52",
          7298 => x"3f",
          7299 => x"08",
          7300 => x"a8",
          7301 => x"86",
          7302 => x"52",
          7303 => x"bc",
          7304 => x"a8",
          7305 => x"b5",
          7306 => x"38",
          7307 => x"08",
          7308 => x"82",
          7309 => x"86",
          7310 => x"ff",
          7311 => x"3d",
          7312 => x"3f",
          7313 => x"0b",
          7314 => x"08",
          7315 => x"82",
          7316 => x"82",
          7317 => x"80",
          7318 => x"b5",
          7319 => x"3d",
          7320 => x"3d",
          7321 => x"93",
          7322 => x"52",
          7323 => x"e9",
          7324 => x"b5",
          7325 => x"82",
          7326 => x"80",
          7327 => x"58",
          7328 => x"3d",
          7329 => x"e0",
          7330 => x"b5",
          7331 => x"82",
          7332 => x"bc",
          7333 => x"c7",
          7334 => x"98",
          7335 => x"73",
          7336 => x"38",
          7337 => x"12",
          7338 => x"39",
          7339 => x"33",
          7340 => x"70",
          7341 => x"55",
          7342 => x"2e",
          7343 => x"7f",
          7344 => x"54",
          7345 => x"82",
          7346 => x"94",
          7347 => x"39",
          7348 => x"08",
          7349 => x"81",
          7350 => x"85",
          7351 => x"b5",
          7352 => x"3d",
          7353 => x"3d",
          7354 => x"5b",
          7355 => x"34",
          7356 => x"3d",
          7357 => x"52",
          7358 => x"e8",
          7359 => x"b5",
          7360 => x"82",
          7361 => x"82",
          7362 => x"43",
          7363 => x"11",
          7364 => x"58",
          7365 => x"80",
          7366 => x"38",
          7367 => x"3d",
          7368 => x"d5",
          7369 => x"b5",
          7370 => x"82",
          7371 => x"82",
          7372 => x"52",
          7373 => x"c8",
          7374 => x"a8",
          7375 => x"b5",
          7376 => x"c1",
          7377 => x"7b",
          7378 => x"3f",
          7379 => x"08",
          7380 => x"74",
          7381 => x"3f",
          7382 => x"08",
          7383 => x"a8",
          7384 => x"38",
          7385 => x"51",
          7386 => x"82",
          7387 => x"57",
          7388 => x"08",
          7389 => x"52",
          7390 => x"f2",
          7391 => x"b5",
          7392 => x"a6",
          7393 => x"74",
          7394 => x"3f",
          7395 => x"08",
          7396 => x"a8",
          7397 => x"cc",
          7398 => x"2e",
          7399 => x"86",
          7400 => x"81",
          7401 => x"81",
          7402 => x"3d",
          7403 => x"52",
          7404 => x"c9",
          7405 => x"3d",
          7406 => x"11",
          7407 => x"5a",
          7408 => x"2e",
          7409 => x"b9",
          7410 => x"16",
          7411 => x"33",
          7412 => x"73",
          7413 => x"16",
          7414 => x"26",
          7415 => x"75",
          7416 => x"38",
          7417 => x"05",
          7418 => x"6f",
          7419 => x"ff",
          7420 => x"55",
          7421 => x"74",
          7422 => x"38",
          7423 => x"11",
          7424 => x"74",
          7425 => x"39",
          7426 => x"09",
          7427 => x"38",
          7428 => x"11",
          7429 => x"74",
          7430 => x"82",
          7431 => x"70",
          7432 => x"ae",
          7433 => x"08",
          7434 => x"5c",
          7435 => x"73",
          7436 => x"38",
          7437 => x"1a",
          7438 => x"55",
          7439 => x"38",
          7440 => x"73",
          7441 => x"38",
          7442 => x"76",
          7443 => x"74",
          7444 => x"33",
          7445 => x"05",
          7446 => x"15",
          7447 => x"ba",
          7448 => x"05",
          7449 => x"ff",
          7450 => x"06",
          7451 => x"57",
          7452 => x"18",
          7453 => x"54",
          7454 => x"70",
          7455 => x"34",
          7456 => x"ee",
          7457 => x"34",
          7458 => x"a8",
          7459 => x"0d",
          7460 => x"0d",
          7461 => x"3d",
          7462 => x"71",
          7463 => x"ec",
          7464 => x"b5",
          7465 => x"82",
          7466 => x"82",
          7467 => x"15",
          7468 => x"82",
          7469 => x"15",
          7470 => x"76",
          7471 => x"90",
          7472 => x"81",
          7473 => x"06",
          7474 => x"72",
          7475 => x"56",
          7476 => x"54",
          7477 => x"17",
          7478 => x"78",
          7479 => x"38",
          7480 => x"22",
          7481 => x"59",
          7482 => x"78",
          7483 => x"76",
          7484 => x"51",
          7485 => x"3f",
          7486 => x"08",
          7487 => x"54",
          7488 => x"53",
          7489 => x"3f",
          7490 => x"08",
          7491 => x"38",
          7492 => x"75",
          7493 => x"18",
          7494 => x"31",
          7495 => x"57",
          7496 => x"b1",
          7497 => x"08",
          7498 => x"38",
          7499 => x"51",
          7500 => x"82",
          7501 => x"54",
          7502 => x"08",
          7503 => x"9a",
          7504 => x"a8",
          7505 => x"81",
          7506 => x"b5",
          7507 => x"16",
          7508 => x"16",
          7509 => x"2e",
          7510 => x"76",
          7511 => x"dc",
          7512 => x"31",
          7513 => x"18",
          7514 => x"90",
          7515 => x"81",
          7516 => x"06",
          7517 => x"56",
          7518 => x"9a",
          7519 => x"74",
          7520 => x"3f",
          7521 => x"08",
          7522 => x"a8",
          7523 => x"82",
          7524 => x"56",
          7525 => x"52",
          7526 => x"84",
          7527 => x"a8",
          7528 => x"ff",
          7529 => x"81",
          7530 => x"38",
          7531 => x"98",
          7532 => x"a6",
          7533 => x"16",
          7534 => x"39",
          7535 => x"16",
          7536 => x"75",
          7537 => x"53",
          7538 => x"aa",
          7539 => x"79",
          7540 => x"3f",
          7541 => x"08",
          7542 => x"0b",
          7543 => x"82",
          7544 => x"39",
          7545 => x"16",
          7546 => x"bb",
          7547 => x"2a",
          7548 => x"08",
          7549 => x"15",
          7550 => x"15",
          7551 => x"90",
          7552 => x"16",
          7553 => x"33",
          7554 => x"53",
          7555 => x"34",
          7556 => x"06",
          7557 => x"2e",
          7558 => x"9c",
          7559 => x"85",
          7560 => x"16",
          7561 => x"72",
          7562 => x"0c",
          7563 => x"04",
          7564 => x"79",
          7565 => x"75",
          7566 => x"8a",
          7567 => x"89",
          7568 => x"52",
          7569 => x"05",
          7570 => x"3f",
          7571 => x"08",
          7572 => x"a8",
          7573 => x"38",
          7574 => x"7a",
          7575 => x"d8",
          7576 => x"b5",
          7577 => x"82",
          7578 => x"80",
          7579 => x"16",
          7580 => x"2b",
          7581 => x"74",
          7582 => x"86",
          7583 => x"84",
          7584 => x"06",
          7585 => x"73",
          7586 => x"38",
          7587 => x"52",
          7588 => x"da",
          7589 => x"a8",
          7590 => x"0c",
          7591 => x"14",
          7592 => x"23",
          7593 => x"51",
          7594 => x"82",
          7595 => x"55",
          7596 => x"09",
          7597 => x"38",
          7598 => x"39",
          7599 => x"84",
          7600 => x"0c",
          7601 => x"82",
          7602 => x"89",
          7603 => x"fc",
          7604 => x"87",
          7605 => x"53",
          7606 => x"e7",
          7607 => x"b5",
          7608 => x"38",
          7609 => x"08",
          7610 => x"3d",
          7611 => x"3d",
          7612 => x"89",
          7613 => x"54",
          7614 => x"54",
          7615 => x"82",
          7616 => x"53",
          7617 => x"08",
          7618 => x"74",
          7619 => x"b5",
          7620 => x"73",
          7621 => x"3f",
          7622 => x"08",
          7623 => x"39",
          7624 => x"08",
          7625 => x"d3",
          7626 => x"b5",
          7627 => x"82",
          7628 => x"84",
          7629 => x"06",
          7630 => x"53",
          7631 => x"b5",
          7632 => x"38",
          7633 => x"51",
          7634 => x"72",
          7635 => x"cf",
          7636 => x"b5",
          7637 => x"32",
          7638 => x"72",
          7639 => x"70",
          7640 => x"08",
          7641 => x"54",
          7642 => x"b5",
          7643 => x"3d",
          7644 => x"3d",
          7645 => x"80",
          7646 => x"70",
          7647 => x"52",
          7648 => x"3f",
          7649 => x"08",
          7650 => x"a8",
          7651 => x"64",
          7652 => x"d6",
          7653 => x"b5",
          7654 => x"82",
          7655 => x"a0",
          7656 => x"cb",
          7657 => x"98",
          7658 => x"73",
          7659 => x"38",
          7660 => x"39",
          7661 => x"88",
          7662 => x"75",
          7663 => x"3f",
          7664 => x"a8",
          7665 => x"0d",
          7666 => x"0d",
          7667 => x"5c",
          7668 => x"3d",
          7669 => x"93",
          7670 => x"d6",
          7671 => x"a8",
          7672 => x"b5",
          7673 => x"80",
          7674 => x"0c",
          7675 => x"11",
          7676 => x"90",
          7677 => x"56",
          7678 => x"74",
          7679 => x"75",
          7680 => x"e4",
          7681 => x"81",
          7682 => x"5b",
          7683 => x"82",
          7684 => x"75",
          7685 => x"73",
          7686 => x"81",
          7687 => x"82",
          7688 => x"76",
          7689 => x"f0",
          7690 => x"f4",
          7691 => x"a8",
          7692 => x"d1",
          7693 => x"a8",
          7694 => x"ce",
          7695 => x"a8",
          7696 => x"82",
          7697 => x"07",
          7698 => x"05",
          7699 => x"53",
          7700 => x"98",
          7701 => x"26",
          7702 => x"f9",
          7703 => x"08",
          7704 => x"08",
          7705 => x"98",
          7706 => x"81",
          7707 => x"58",
          7708 => x"3f",
          7709 => x"08",
          7710 => x"a8",
          7711 => x"38",
          7712 => x"77",
          7713 => x"5d",
          7714 => x"74",
          7715 => x"81",
          7716 => x"b4",
          7717 => x"bb",
          7718 => x"b5",
          7719 => x"ff",
          7720 => x"30",
          7721 => x"1b",
          7722 => x"5b",
          7723 => x"39",
          7724 => x"ff",
          7725 => x"82",
          7726 => x"f0",
          7727 => x"30",
          7728 => x"1b",
          7729 => x"5b",
          7730 => x"83",
          7731 => x"58",
          7732 => x"92",
          7733 => x"0c",
          7734 => x"12",
          7735 => x"33",
          7736 => x"54",
          7737 => x"34",
          7738 => x"a8",
          7739 => x"0d",
          7740 => x"0d",
          7741 => x"fc",
          7742 => x"52",
          7743 => x"3f",
          7744 => x"08",
          7745 => x"a8",
          7746 => x"38",
          7747 => x"56",
          7748 => x"38",
          7749 => x"70",
          7750 => x"81",
          7751 => x"55",
          7752 => x"80",
          7753 => x"38",
          7754 => x"54",
          7755 => x"08",
          7756 => x"38",
          7757 => x"82",
          7758 => x"53",
          7759 => x"52",
          7760 => x"8c",
          7761 => x"a8",
          7762 => x"19",
          7763 => x"c9",
          7764 => x"08",
          7765 => x"ff",
          7766 => x"82",
          7767 => x"ff",
          7768 => x"06",
          7769 => x"56",
          7770 => x"08",
          7771 => x"81",
          7772 => x"82",
          7773 => x"75",
          7774 => x"54",
          7775 => x"08",
          7776 => x"27",
          7777 => x"17",
          7778 => x"b5",
          7779 => x"76",
          7780 => x"3f",
          7781 => x"08",
          7782 => x"08",
          7783 => x"90",
          7784 => x"c0",
          7785 => x"90",
          7786 => x"80",
          7787 => x"75",
          7788 => x"75",
          7789 => x"b5",
          7790 => x"3d",
          7791 => x"3d",
          7792 => x"a0",
          7793 => x"05",
          7794 => x"51",
          7795 => x"82",
          7796 => x"55",
          7797 => x"08",
          7798 => x"78",
          7799 => x"08",
          7800 => x"70",
          7801 => x"ae",
          7802 => x"a8",
          7803 => x"b5",
          7804 => x"db",
          7805 => x"fb",
          7806 => x"85",
          7807 => x"06",
          7808 => x"86",
          7809 => x"c7",
          7810 => x"2b",
          7811 => x"24",
          7812 => x"02",
          7813 => x"33",
          7814 => x"58",
          7815 => x"76",
          7816 => x"6b",
          7817 => x"cc",
          7818 => x"b5",
          7819 => x"84",
          7820 => x"06",
          7821 => x"73",
          7822 => x"d4",
          7823 => x"82",
          7824 => x"94",
          7825 => x"81",
          7826 => x"5a",
          7827 => x"08",
          7828 => x"8a",
          7829 => x"54",
          7830 => x"82",
          7831 => x"55",
          7832 => x"08",
          7833 => x"82",
          7834 => x"52",
          7835 => x"e5",
          7836 => x"a8",
          7837 => x"b5",
          7838 => x"38",
          7839 => x"cf",
          7840 => x"a8",
          7841 => x"88",
          7842 => x"a8",
          7843 => x"38",
          7844 => x"c2",
          7845 => x"a8",
          7846 => x"a8",
          7847 => x"82",
          7848 => x"07",
          7849 => x"55",
          7850 => x"2e",
          7851 => x"80",
          7852 => x"80",
          7853 => x"77",
          7854 => x"3f",
          7855 => x"08",
          7856 => x"38",
          7857 => x"ba",
          7858 => x"b5",
          7859 => x"74",
          7860 => x"0c",
          7861 => x"04",
          7862 => x"82",
          7863 => x"c0",
          7864 => x"3d",
          7865 => x"3f",
          7866 => x"08",
          7867 => x"a8",
          7868 => x"38",
          7869 => x"52",
          7870 => x"52",
          7871 => x"3f",
          7872 => x"08",
          7873 => x"a8",
          7874 => x"88",
          7875 => x"39",
          7876 => x"08",
          7877 => x"81",
          7878 => x"38",
          7879 => x"05",
          7880 => x"2a",
          7881 => x"55",
          7882 => x"81",
          7883 => x"5a",
          7884 => x"3d",
          7885 => x"c1",
          7886 => x"b5",
          7887 => x"55",
          7888 => x"a8",
          7889 => x"87",
          7890 => x"a8",
          7891 => x"09",
          7892 => x"38",
          7893 => x"b5",
          7894 => x"2e",
          7895 => x"86",
          7896 => x"81",
          7897 => x"81",
          7898 => x"b5",
          7899 => x"78",
          7900 => x"3f",
          7901 => x"08",
          7902 => x"a8",
          7903 => x"38",
          7904 => x"52",
          7905 => x"ff",
          7906 => x"78",
          7907 => x"b4",
          7908 => x"54",
          7909 => x"15",
          7910 => x"b2",
          7911 => x"ca",
          7912 => x"b6",
          7913 => x"53",
          7914 => x"53",
          7915 => x"3f",
          7916 => x"b4",
          7917 => x"d4",
          7918 => x"b6",
          7919 => x"54",
          7920 => x"d5",
          7921 => x"53",
          7922 => x"11",
          7923 => x"d7",
          7924 => x"81",
          7925 => x"34",
          7926 => x"a4",
          7927 => x"a8",
          7928 => x"b5",
          7929 => x"38",
          7930 => x"0a",
          7931 => x"05",
          7932 => x"d0",
          7933 => x"64",
          7934 => x"c9",
          7935 => x"54",
          7936 => x"15",
          7937 => x"81",
          7938 => x"34",
          7939 => x"b8",
          7940 => x"b5",
          7941 => x"8b",
          7942 => x"75",
          7943 => x"ff",
          7944 => x"73",
          7945 => x"0c",
          7946 => x"04",
          7947 => x"a9",
          7948 => x"51",
          7949 => x"82",
          7950 => x"ff",
          7951 => x"a9",
          7952 => x"ee",
          7953 => x"a8",
          7954 => x"b5",
          7955 => x"d3",
          7956 => x"a9",
          7957 => x"9d",
          7958 => x"58",
          7959 => x"82",
          7960 => x"55",
          7961 => x"08",
          7962 => x"02",
          7963 => x"33",
          7964 => x"54",
          7965 => x"82",
          7966 => x"53",
          7967 => x"52",
          7968 => x"88",
          7969 => x"b4",
          7970 => x"53",
          7971 => x"3d",
          7972 => x"ff",
          7973 => x"aa",
          7974 => x"73",
          7975 => x"3f",
          7976 => x"08",
          7977 => x"a8",
          7978 => x"63",
          7979 => x"81",
          7980 => x"65",
          7981 => x"2e",
          7982 => x"55",
          7983 => x"82",
          7984 => x"84",
          7985 => x"06",
          7986 => x"73",
          7987 => x"3f",
          7988 => x"08",
          7989 => x"a8",
          7990 => x"38",
          7991 => x"53",
          7992 => x"95",
          7993 => x"16",
          7994 => x"87",
          7995 => x"05",
          7996 => x"34",
          7997 => x"70",
          7998 => x"81",
          7999 => x"55",
          8000 => x"74",
          8001 => x"73",
          8002 => x"78",
          8003 => x"83",
          8004 => x"16",
          8005 => x"2a",
          8006 => x"51",
          8007 => x"80",
          8008 => x"38",
          8009 => x"80",
          8010 => x"52",
          8011 => x"be",
          8012 => x"a8",
          8013 => x"51",
          8014 => x"3f",
          8015 => x"b5",
          8016 => x"2e",
          8017 => x"82",
          8018 => x"52",
          8019 => x"b5",
          8020 => x"b5",
          8021 => x"80",
          8022 => x"58",
          8023 => x"a8",
          8024 => x"38",
          8025 => x"54",
          8026 => x"09",
          8027 => x"38",
          8028 => x"52",
          8029 => x"af",
          8030 => x"81",
          8031 => x"34",
          8032 => x"b5",
          8033 => x"38",
          8034 => x"ca",
          8035 => x"a8",
          8036 => x"b5",
          8037 => x"38",
          8038 => x"b5",
          8039 => x"b5",
          8040 => x"74",
          8041 => x"0c",
          8042 => x"04",
          8043 => x"02",
          8044 => x"33",
          8045 => x"80",
          8046 => x"57",
          8047 => x"95",
          8048 => x"52",
          8049 => x"d2",
          8050 => x"b5",
          8051 => x"82",
          8052 => x"80",
          8053 => x"5a",
          8054 => x"3d",
          8055 => x"c9",
          8056 => x"b5",
          8057 => x"82",
          8058 => x"b8",
          8059 => x"cf",
          8060 => x"a0",
          8061 => x"55",
          8062 => x"75",
          8063 => x"71",
          8064 => x"33",
          8065 => x"74",
          8066 => x"57",
          8067 => x"8b",
          8068 => x"54",
          8069 => x"15",
          8070 => x"ff",
          8071 => x"82",
          8072 => x"55",
          8073 => x"a8",
          8074 => x"0d",
          8075 => x"0d",
          8076 => x"53",
          8077 => x"05",
          8078 => x"51",
          8079 => x"82",
          8080 => x"55",
          8081 => x"08",
          8082 => x"76",
          8083 => x"93",
          8084 => x"51",
          8085 => x"82",
          8086 => x"55",
          8087 => x"08",
          8088 => x"80",
          8089 => x"81",
          8090 => x"86",
          8091 => x"38",
          8092 => x"86",
          8093 => x"90",
          8094 => x"54",
          8095 => x"ff",
          8096 => x"76",
          8097 => x"83",
          8098 => x"51",
          8099 => x"3f",
          8100 => x"08",
          8101 => x"b5",
          8102 => x"3d",
          8103 => x"3d",
          8104 => x"5c",
          8105 => x"98",
          8106 => x"52",
          8107 => x"d1",
          8108 => x"b5",
          8109 => x"b5",
          8110 => x"70",
          8111 => x"08",
          8112 => x"51",
          8113 => x"80",
          8114 => x"38",
          8115 => x"06",
          8116 => x"80",
          8117 => x"38",
          8118 => x"5f",
          8119 => x"3d",
          8120 => x"ff",
          8121 => x"82",
          8122 => x"57",
          8123 => x"08",
          8124 => x"74",
          8125 => x"c3",
          8126 => x"b5",
          8127 => x"82",
          8128 => x"bf",
          8129 => x"a8",
          8130 => x"a8",
          8131 => x"59",
          8132 => x"81",
          8133 => x"56",
          8134 => x"33",
          8135 => x"16",
          8136 => x"27",
          8137 => x"56",
          8138 => x"80",
          8139 => x"80",
          8140 => x"ff",
          8141 => x"70",
          8142 => x"56",
          8143 => x"e8",
          8144 => x"76",
          8145 => x"81",
          8146 => x"80",
          8147 => x"57",
          8148 => x"78",
          8149 => x"51",
          8150 => x"2e",
          8151 => x"73",
          8152 => x"38",
          8153 => x"08",
          8154 => x"b1",
          8155 => x"b5",
          8156 => x"82",
          8157 => x"a7",
          8158 => x"33",
          8159 => x"c3",
          8160 => x"2e",
          8161 => x"e4",
          8162 => x"2e",
          8163 => x"56",
          8164 => x"05",
          8165 => x"e3",
          8166 => x"a8",
          8167 => x"76",
          8168 => x"0c",
          8169 => x"04",
          8170 => x"82",
          8171 => x"ff",
          8172 => x"9d",
          8173 => x"fa",
          8174 => x"a8",
          8175 => x"a8",
          8176 => x"82",
          8177 => x"83",
          8178 => x"53",
          8179 => x"3d",
          8180 => x"ff",
          8181 => x"73",
          8182 => x"70",
          8183 => x"52",
          8184 => x"9f",
          8185 => x"bc",
          8186 => x"74",
          8187 => x"6d",
          8188 => x"70",
          8189 => x"af",
          8190 => x"b5",
          8191 => x"2e",
          8192 => x"70",
          8193 => x"57",
          8194 => x"fd",
          8195 => x"a8",
          8196 => x"8d",
          8197 => x"2b",
          8198 => x"81",
          8199 => x"86",
          8200 => x"a8",
          8201 => x"9f",
          8202 => x"ff",
          8203 => x"54",
          8204 => x"8a",
          8205 => x"70",
          8206 => x"06",
          8207 => x"ff",
          8208 => x"38",
          8209 => x"15",
          8210 => x"80",
          8211 => x"74",
          8212 => x"f0",
          8213 => x"89",
          8214 => x"a8",
          8215 => x"81",
          8216 => x"88",
          8217 => x"26",
          8218 => x"39",
          8219 => x"86",
          8220 => x"81",
          8221 => x"ff",
          8222 => x"38",
          8223 => x"54",
          8224 => x"81",
          8225 => x"81",
          8226 => x"78",
          8227 => x"5a",
          8228 => x"6d",
          8229 => x"81",
          8230 => x"57",
          8231 => x"9f",
          8232 => x"38",
          8233 => x"54",
          8234 => x"81",
          8235 => x"b1",
          8236 => x"2e",
          8237 => x"a7",
          8238 => x"15",
          8239 => x"54",
          8240 => x"09",
          8241 => x"38",
          8242 => x"76",
          8243 => x"41",
          8244 => x"52",
          8245 => x"52",
          8246 => x"b3",
          8247 => x"a8",
          8248 => x"b5",
          8249 => x"f7",
          8250 => x"74",
          8251 => x"e5",
          8252 => x"a8",
          8253 => x"b5",
          8254 => x"38",
          8255 => x"38",
          8256 => x"74",
          8257 => x"39",
          8258 => x"08",
          8259 => x"81",
          8260 => x"38",
          8261 => x"74",
          8262 => x"38",
          8263 => x"51",
          8264 => x"3f",
          8265 => x"08",
          8266 => x"a8",
          8267 => x"a0",
          8268 => x"a8",
          8269 => x"51",
          8270 => x"3f",
          8271 => x"0b",
          8272 => x"8b",
          8273 => x"67",
          8274 => x"a7",
          8275 => x"81",
          8276 => x"34",
          8277 => x"ad",
          8278 => x"b5",
          8279 => x"73",
          8280 => x"b5",
          8281 => x"3d",
          8282 => x"3d",
          8283 => x"02",
          8284 => x"cb",
          8285 => x"3d",
          8286 => x"72",
          8287 => x"5a",
          8288 => x"82",
          8289 => x"58",
          8290 => x"08",
          8291 => x"91",
          8292 => x"77",
          8293 => x"7c",
          8294 => x"38",
          8295 => x"59",
          8296 => x"90",
          8297 => x"81",
          8298 => x"06",
          8299 => x"73",
          8300 => x"54",
          8301 => x"82",
          8302 => x"39",
          8303 => x"8b",
          8304 => x"11",
          8305 => x"2b",
          8306 => x"54",
          8307 => x"fe",
          8308 => x"ff",
          8309 => x"70",
          8310 => x"07",
          8311 => x"b5",
          8312 => x"8c",
          8313 => x"40",
          8314 => x"55",
          8315 => x"88",
          8316 => x"08",
          8317 => x"38",
          8318 => x"77",
          8319 => x"56",
          8320 => x"51",
          8321 => x"3f",
          8322 => x"55",
          8323 => x"08",
          8324 => x"38",
          8325 => x"b5",
          8326 => x"2e",
          8327 => x"82",
          8328 => x"ff",
          8329 => x"38",
          8330 => x"08",
          8331 => x"16",
          8332 => x"2e",
          8333 => x"87",
          8334 => x"74",
          8335 => x"74",
          8336 => x"81",
          8337 => x"38",
          8338 => x"ff",
          8339 => x"2e",
          8340 => x"7b",
          8341 => x"80",
          8342 => x"81",
          8343 => x"81",
          8344 => x"06",
          8345 => x"56",
          8346 => x"52",
          8347 => x"af",
          8348 => x"b5",
          8349 => x"82",
          8350 => x"80",
          8351 => x"81",
          8352 => x"56",
          8353 => x"d3",
          8354 => x"ff",
          8355 => x"7c",
          8356 => x"55",
          8357 => x"b3",
          8358 => x"1b",
          8359 => x"1b",
          8360 => x"33",
          8361 => x"54",
          8362 => x"34",
          8363 => x"fe",
          8364 => x"08",
          8365 => x"74",
          8366 => x"75",
          8367 => x"16",
          8368 => x"33",
          8369 => x"73",
          8370 => x"77",
          8371 => x"b5",
          8372 => x"3d",
          8373 => x"3d",
          8374 => x"02",
          8375 => x"eb",
          8376 => x"3d",
          8377 => x"59",
          8378 => x"8b",
          8379 => x"82",
          8380 => x"24",
          8381 => x"82",
          8382 => x"84",
          8383 => x"e0",
          8384 => x"51",
          8385 => x"2e",
          8386 => x"75",
          8387 => x"a8",
          8388 => x"06",
          8389 => x"7e",
          8390 => x"d0",
          8391 => x"a8",
          8392 => x"06",
          8393 => x"56",
          8394 => x"74",
          8395 => x"76",
          8396 => x"81",
          8397 => x"8a",
          8398 => x"b2",
          8399 => x"fc",
          8400 => x"52",
          8401 => x"a4",
          8402 => x"b5",
          8403 => x"38",
          8404 => x"80",
          8405 => x"74",
          8406 => x"26",
          8407 => x"15",
          8408 => x"74",
          8409 => x"38",
          8410 => x"80",
          8411 => x"84",
          8412 => x"92",
          8413 => x"80",
          8414 => x"38",
          8415 => x"06",
          8416 => x"2e",
          8417 => x"56",
          8418 => x"78",
          8419 => x"89",
          8420 => x"2b",
          8421 => x"43",
          8422 => x"38",
          8423 => x"30",
          8424 => x"77",
          8425 => x"91",
          8426 => x"c2",
          8427 => x"f8",
          8428 => x"52",
          8429 => x"a4",
          8430 => x"56",
          8431 => x"08",
          8432 => x"77",
          8433 => x"77",
          8434 => x"a8",
          8435 => x"45",
          8436 => x"bf",
          8437 => x"8e",
          8438 => x"26",
          8439 => x"74",
          8440 => x"48",
          8441 => x"75",
          8442 => x"38",
          8443 => x"81",
          8444 => x"fa",
          8445 => x"2a",
          8446 => x"56",
          8447 => x"2e",
          8448 => x"87",
          8449 => x"82",
          8450 => x"38",
          8451 => x"55",
          8452 => x"83",
          8453 => x"81",
          8454 => x"56",
          8455 => x"80",
          8456 => x"38",
          8457 => x"83",
          8458 => x"06",
          8459 => x"78",
          8460 => x"91",
          8461 => x"0b",
          8462 => x"22",
          8463 => x"80",
          8464 => x"74",
          8465 => x"38",
          8466 => x"56",
          8467 => x"17",
          8468 => x"57",
          8469 => x"2e",
          8470 => x"75",
          8471 => x"79",
          8472 => x"fe",
          8473 => x"82",
          8474 => x"84",
          8475 => x"05",
          8476 => x"5e",
          8477 => x"80",
          8478 => x"a8",
          8479 => x"8a",
          8480 => x"fd",
          8481 => x"75",
          8482 => x"38",
          8483 => x"78",
          8484 => x"8c",
          8485 => x"0b",
          8486 => x"22",
          8487 => x"80",
          8488 => x"74",
          8489 => x"38",
          8490 => x"56",
          8491 => x"17",
          8492 => x"57",
          8493 => x"2e",
          8494 => x"75",
          8495 => x"79",
          8496 => x"fe",
          8497 => x"82",
          8498 => x"10",
          8499 => x"82",
          8500 => x"9f",
          8501 => x"38",
          8502 => x"b5",
          8503 => x"82",
          8504 => x"05",
          8505 => x"2a",
          8506 => x"56",
          8507 => x"17",
          8508 => x"81",
          8509 => x"60",
          8510 => x"65",
          8511 => x"12",
          8512 => x"30",
          8513 => x"74",
          8514 => x"59",
          8515 => x"7d",
          8516 => x"81",
          8517 => x"76",
          8518 => x"41",
          8519 => x"76",
          8520 => x"90",
          8521 => x"62",
          8522 => x"51",
          8523 => x"26",
          8524 => x"75",
          8525 => x"31",
          8526 => x"65",
          8527 => x"fe",
          8528 => x"82",
          8529 => x"58",
          8530 => x"09",
          8531 => x"38",
          8532 => x"08",
          8533 => x"26",
          8534 => x"78",
          8535 => x"79",
          8536 => x"78",
          8537 => x"86",
          8538 => x"82",
          8539 => x"06",
          8540 => x"83",
          8541 => x"82",
          8542 => x"27",
          8543 => x"8f",
          8544 => x"55",
          8545 => x"26",
          8546 => x"59",
          8547 => x"62",
          8548 => x"74",
          8549 => x"38",
          8550 => x"88",
          8551 => x"a8",
          8552 => x"26",
          8553 => x"86",
          8554 => x"1a",
          8555 => x"79",
          8556 => x"38",
          8557 => x"80",
          8558 => x"2e",
          8559 => x"83",
          8560 => x"9f",
          8561 => x"8b",
          8562 => x"06",
          8563 => x"74",
          8564 => x"84",
          8565 => x"52",
          8566 => x"a2",
          8567 => x"53",
          8568 => x"52",
          8569 => x"a2",
          8570 => x"80",
          8571 => x"51",
          8572 => x"3f",
          8573 => x"34",
          8574 => x"ff",
          8575 => x"1b",
          8576 => x"a2",
          8577 => x"90",
          8578 => x"83",
          8579 => x"70",
          8580 => x"80",
          8581 => x"55",
          8582 => x"ff",
          8583 => x"66",
          8584 => x"ff",
          8585 => x"38",
          8586 => x"ff",
          8587 => x"1b",
          8588 => x"f2",
          8589 => x"74",
          8590 => x"51",
          8591 => x"3f",
          8592 => x"1c",
          8593 => x"98",
          8594 => x"a0",
          8595 => x"ff",
          8596 => x"51",
          8597 => x"3f",
          8598 => x"1b",
          8599 => x"e4",
          8600 => x"2e",
          8601 => x"80",
          8602 => x"88",
          8603 => x"80",
          8604 => x"ff",
          8605 => x"7c",
          8606 => x"51",
          8607 => x"3f",
          8608 => x"1b",
          8609 => x"bc",
          8610 => x"b0",
          8611 => x"a0",
          8612 => x"52",
          8613 => x"ff",
          8614 => x"ff",
          8615 => x"c0",
          8616 => x"0b",
          8617 => x"34",
          8618 => x"ae",
          8619 => x"c7",
          8620 => x"39",
          8621 => x"0a",
          8622 => x"51",
          8623 => x"3f",
          8624 => x"ff",
          8625 => x"1b",
          8626 => x"da",
          8627 => x"0b",
          8628 => x"a9",
          8629 => x"34",
          8630 => x"ae",
          8631 => x"1b",
          8632 => x"8f",
          8633 => x"d5",
          8634 => x"1b",
          8635 => x"ff",
          8636 => x"81",
          8637 => x"7a",
          8638 => x"ff",
          8639 => x"81",
          8640 => x"a8",
          8641 => x"38",
          8642 => x"09",
          8643 => x"ee",
          8644 => x"60",
          8645 => x"7a",
          8646 => x"ff",
          8647 => x"84",
          8648 => x"52",
          8649 => x"9f",
          8650 => x"8b",
          8651 => x"52",
          8652 => x"9f",
          8653 => x"8a",
          8654 => x"52",
          8655 => x"51",
          8656 => x"3f",
          8657 => x"83",
          8658 => x"ff",
          8659 => x"82",
          8660 => x"1b",
          8661 => x"ec",
          8662 => x"d5",
          8663 => x"ff",
          8664 => x"75",
          8665 => x"05",
          8666 => x"7e",
          8667 => x"e5",
          8668 => x"60",
          8669 => x"52",
          8670 => x"9a",
          8671 => x"53",
          8672 => x"51",
          8673 => x"3f",
          8674 => x"58",
          8675 => x"09",
          8676 => x"38",
          8677 => x"51",
          8678 => x"3f",
          8679 => x"1b",
          8680 => x"a0",
          8681 => x"52",
          8682 => x"91",
          8683 => x"ff",
          8684 => x"81",
          8685 => x"f8",
          8686 => x"7a",
          8687 => x"84",
          8688 => x"61",
          8689 => x"26",
          8690 => x"57",
          8691 => x"53",
          8692 => x"51",
          8693 => x"3f",
          8694 => x"08",
          8695 => x"84",
          8696 => x"b5",
          8697 => x"7a",
          8698 => x"aa",
          8699 => x"75",
          8700 => x"56",
          8701 => x"81",
          8702 => x"80",
          8703 => x"38",
          8704 => x"83",
          8705 => x"63",
          8706 => x"74",
          8707 => x"38",
          8708 => x"54",
          8709 => x"52",
          8710 => x"99",
          8711 => x"b5",
          8712 => x"c1",
          8713 => x"75",
          8714 => x"56",
          8715 => x"8c",
          8716 => x"2e",
          8717 => x"56",
          8718 => x"ff",
          8719 => x"84",
          8720 => x"2e",
          8721 => x"56",
          8722 => x"58",
          8723 => x"38",
          8724 => x"77",
          8725 => x"ff",
          8726 => x"82",
          8727 => x"78",
          8728 => x"c2",
          8729 => x"1b",
          8730 => x"34",
          8731 => x"16",
          8732 => x"82",
          8733 => x"83",
          8734 => x"84",
          8735 => x"67",
          8736 => x"fd",
          8737 => x"51",
          8738 => x"3f",
          8739 => x"16",
          8740 => x"a8",
          8741 => x"bf",
          8742 => x"86",
          8743 => x"b5",
          8744 => x"16",
          8745 => x"83",
          8746 => x"ff",
          8747 => x"66",
          8748 => x"1b",
          8749 => x"8c",
          8750 => x"77",
          8751 => x"7e",
          8752 => x"91",
          8753 => x"82",
          8754 => x"a2",
          8755 => x"80",
          8756 => x"ff",
          8757 => x"81",
          8758 => x"a8",
          8759 => x"89",
          8760 => x"8a",
          8761 => x"86",
          8762 => x"a8",
          8763 => x"82",
          8764 => x"99",
          8765 => x"f5",
          8766 => x"60",
          8767 => x"79",
          8768 => x"5a",
          8769 => x"78",
          8770 => x"8d",
          8771 => x"55",
          8772 => x"fc",
          8773 => x"51",
          8774 => x"7a",
          8775 => x"81",
          8776 => x"8c",
          8777 => x"74",
          8778 => x"38",
          8779 => x"81",
          8780 => x"81",
          8781 => x"8a",
          8782 => x"06",
          8783 => x"76",
          8784 => x"76",
          8785 => x"55",
          8786 => x"a8",
          8787 => x"0d",
          8788 => x"0d",
          8789 => x"05",
          8790 => x"59",
          8791 => x"2e",
          8792 => x"87",
          8793 => x"76",
          8794 => x"84",
          8795 => x"80",
          8796 => x"38",
          8797 => x"77",
          8798 => x"56",
          8799 => x"34",
          8800 => x"bb",
          8801 => x"38",
          8802 => x"05",
          8803 => x"8c",
          8804 => x"08",
          8805 => x"3f",
          8806 => x"70",
          8807 => x"07",
          8808 => x"30",
          8809 => x"56",
          8810 => x"0c",
          8811 => x"18",
          8812 => x"0d",
          8813 => x"0d",
          8814 => x"08",
          8815 => x"75",
          8816 => x"89",
          8817 => x"54",
          8818 => x"16",
          8819 => x"51",
          8820 => x"82",
          8821 => x"91",
          8822 => x"08",
          8823 => x"81",
          8824 => x"88",
          8825 => x"83",
          8826 => x"74",
          8827 => x"0c",
          8828 => x"04",
          8829 => x"75",
          8830 => x"53",
          8831 => x"51",
          8832 => x"3f",
          8833 => x"85",
          8834 => x"ea",
          8835 => x"80",
          8836 => x"6a",
          8837 => x"70",
          8838 => x"d8",
          8839 => x"72",
          8840 => x"3f",
          8841 => x"8d",
          8842 => x"0d",
          8843 => x"00",
          8844 => x"ff",
          8845 => x"ff",
          8846 => x"ff",
          8847 => x"00",
          8848 => x"a8",
          8849 => x"2c",
          8850 => x"33",
          8851 => x"3a",
          8852 => x"41",
          8853 => x"48",
          8854 => x"4f",
          8855 => x"56",
          8856 => x"5d",
          8857 => x"64",
          8858 => x"6b",
          8859 => x"72",
          8860 => x"78",
          8861 => x"7e",
          8862 => x"84",
          8863 => x"8a",
          8864 => x"90",
          8865 => x"96",
          8866 => x"9c",
          8867 => x"a2",
          8868 => x"3b",
          8869 => x"41",
          8870 => x"47",
          8871 => x"4d",
          8872 => x"53",
          8873 => x"20",
          8874 => x"16",
          8875 => x"0e",
          8876 => x"48",
          8877 => x"fe",
          8878 => x"f5",
          8879 => x"c2",
          8880 => x"1e",
          8881 => x"00",
          8882 => x"96",
          8883 => x"1c",
          8884 => x"bd",
          8885 => x"f5",
          8886 => x"0e",
          8887 => x"32",
          8888 => x"c2",
          8889 => x"f5",
          8890 => x"f5",
          8891 => x"1c",
          8892 => x"96",
          8893 => x"1e",
          8894 => x"48",
          8895 => x"2f",
          8896 => x"18",
          8897 => x"18",
          8898 => x"5e",
          8899 => x"18",
          8900 => x"18",
          8901 => x"18",
          8902 => x"18",
          8903 => x"18",
          8904 => x"18",
          8905 => x"18",
          8906 => x"1b",
          8907 => x"18",
          8908 => x"46",
          8909 => x"76",
          8910 => x"18",
          8911 => x"18",
          8912 => x"18",
          8913 => x"18",
          8914 => x"18",
          8915 => x"18",
          8916 => x"18",
          8917 => x"18",
          8918 => x"18",
          8919 => x"18",
          8920 => x"18",
          8921 => x"18",
          8922 => x"18",
          8923 => x"18",
          8924 => x"18",
          8925 => x"18",
          8926 => x"18",
          8927 => x"18",
          8928 => x"18",
          8929 => x"18",
          8930 => x"18",
          8931 => x"18",
          8932 => x"18",
          8933 => x"18",
          8934 => x"18",
          8935 => x"18",
          8936 => x"18",
          8937 => x"18",
          8938 => x"18",
          8939 => x"18",
          8940 => x"18",
          8941 => x"18",
          8942 => x"18",
          8943 => x"18",
          8944 => x"18",
          8945 => x"18",
          8946 => x"a6",
          8947 => x"18",
          8948 => x"18",
          8949 => x"18",
          8950 => x"18",
          8951 => x"14",
          8952 => x"18",
          8953 => x"18",
          8954 => x"18",
          8955 => x"18",
          8956 => x"18",
          8957 => x"18",
          8958 => x"18",
          8959 => x"18",
          8960 => x"18",
          8961 => x"18",
          8962 => x"d6",
          8963 => x"3d",
          8964 => x"ad",
          8965 => x"ad",
          8966 => x"ad",
          8967 => x"18",
          8968 => x"3d",
          8969 => x"18",
          8970 => x"18",
          8971 => x"96",
          8972 => x"18",
          8973 => x"18",
          8974 => x"ea",
          8975 => x"f5",
          8976 => x"18",
          8977 => x"18",
          8978 => x"0f",
          8979 => x"18",
          8980 => x"1d",
          8981 => x"18",
          8982 => x"18",
          8983 => x"14",
          8984 => x"69",
          8985 => x"00",
          8986 => x"63",
          8987 => x"00",
          8988 => x"69",
          8989 => x"00",
          8990 => x"61",
          8991 => x"00",
          8992 => x"65",
          8993 => x"00",
          8994 => x"65",
          8995 => x"00",
          8996 => x"70",
          8997 => x"00",
          8998 => x"66",
          8999 => x"00",
          9000 => x"6d",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"6c",
          9010 => x"00",
          9011 => x"00",
          9012 => x"74",
          9013 => x"00",
          9014 => x"65",
          9015 => x"00",
          9016 => x"6f",
          9017 => x"00",
          9018 => x"74",
          9019 => x"00",
          9020 => x"73",
          9021 => x"00",
          9022 => x"73",
          9023 => x"00",
          9024 => x"6f",
          9025 => x"00",
          9026 => x"00",
          9027 => x"6b",
          9028 => x"72",
          9029 => x"00",
          9030 => x"65",
          9031 => x"6c",
          9032 => x"72",
          9033 => x"0a",
          9034 => x"00",
          9035 => x"6b",
          9036 => x"74",
          9037 => x"61",
          9038 => x"0a",
          9039 => x"00",
          9040 => x"66",
          9041 => x"20",
          9042 => x"6e",
          9043 => x"00",
          9044 => x"70",
          9045 => x"20",
          9046 => x"6e",
          9047 => x"00",
          9048 => x"61",
          9049 => x"20",
          9050 => x"65",
          9051 => x"65",
          9052 => x"00",
          9053 => x"65",
          9054 => x"64",
          9055 => x"65",
          9056 => x"00",
          9057 => x"65",
          9058 => x"72",
          9059 => x"79",
          9060 => x"69",
          9061 => x"2e",
          9062 => x"00",
          9063 => x"65",
          9064 => x"6e",
          9065 => x"20",
          9066 => x"61",
          9067 => x"2e",
          9068 => x"00",
          9069 => x"69",
          9070 => x"72",
          9071 => x"20",
          9072 => x"74",
          9073 => x"65",
          9074 => x"00",
          9075 => x"76",
          9076 => x"75",
          9077 => x"72",
          9078 => x"20",
          9079 => x"61",
          9080 => x"2e",
          9081 => x"00",
          9082 => x"6b",
          9083 => x"74",
          9084 => x"61",
          9085 => x"64",
          9086 => x"00",
          9087 => x"63",
          9088 => x"61",
          9089 => x"6c",
          9090 => x"69",
          9091 => x"79",
          9092 => x"6d",
          9093 => x"75",
          9094 => x"6f",
          9095 => x"69",
          9096 => x"0a",
          9097 => x"00",
          9098 => x"6d",
          9099 => x"61",
          9100 => x"74",
          9101 => x"0a",
          9102 => x"00",
          9103 => x"65",
          9104 => x"2c",
          9105 => x"65",
          9106 => x"69",
          9107 => x"63",
          9108 => x"65",
          9109 => x"64",
          9110 => x"00",
          9111 => x"65",
          9112 => x"20",
          9113 => x"6b",
          9114 => x"0a",
          9115 => x"00",
          9116 => x"75",
          9117 => x"63",
          9118 => x"74",
          9119 => x"6d",
          9120 => x"2e",
          9121 => x"00",
          9122 => x"20",
          9123 => x"79",
          9124 => x"65",
          9125 => x"69",
          9126 => x"2e",
          9127 => x"00",
          9128 => x"61",
          9129 => x"65",
          9130 => x"69",
          9131 => x"72",
          9132 => x"74",
          9133 => x"00",
          9134 => x"63",
          9135 => x"2e",
          9136 => x"00",
          9137 => x"6e",
          9138 => x"20",
          9139 => x"6f",
          9140 => x"00",
          9141 => x"75",
          9142 => x"74",
          9143 => x"25",
          9144 => x"74",
          9145 => x"75",
          9146 => x"74",
          9147 => x"73",
          9148 => x"0a",
          9149 => x"00",
          9150 => x"64",
          9151 => x"00",
          9152 => x"58",
          9153 => x"00",
          9154 => x"00",
          9155 => x"58",
          9156 => x"00",
          9157 => x"20",
          9158 => x"20",
          9159 => x"00",
          9160 => x"58",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"00",
          9165 => x"00",
          9166 => x"20",
          9167 => x"28",
          9168 => x"00",
          9169 => x"30",
          9170 => x"30",
          9171 => x"00",
          9172 => x"30",
          9173 => x"00",
          9174 => x"55",
          9175 => x"65",
          9176 => x"30",
          9177 => x"20",
          9178 => x"25",
          9179 => x"2a",
          9180 => x"00",
          9181 => x"20",
          9182 => x"65",
          9183 => x"70",
          9184 => x"61",
          9185 => x"65",
          9186 => x"00",
          9187 => x"65",
          9188 => x"6e",
          9189 => x"72",
          9190 => x"0a",
          9191 => x"00",
          9192 => x"20",
          9193 => x"65",
          9194 => x"70",
          9195 => x"00",
          9196 => x"54",
          9197 => x"44",
          9198 => x"74",
          9199 => x"75",
          9200 => x"00",
          9201 => x"54",
          9202 => x"52",
          9203 => x"74",
          9204 => x"75",
          9205 => x"00",
          9206 => x"54",
          9207 => x"58",
          9208 => x"74",
          9209 => x"75",
          9210 => x"00",
          9211 => x"54",
          9212 => x"58",
          9213 => x"74",
          9214 => x"75",
          9215 => x"00",
          9216 => x"54",
          9217 => x"58",
          9218 => x"74",
          9219 => x"75",
          9220 => x"00",
          9221 => x"54",
          9222 => x"58",
          9223 => x"74",
          9224 => x"75",
          9225 => x"00",
          9226 => x"74",
          9227 => x"20",
          9228 => x"74",
          9229 => x"72",
          9230 => x"0a",
          9231 => x"00",
          9232 => x"62",
          9233 => x"67",
          9234 => x"6d",
          9235 => x"2e",
          9236 => x"00",
          9237 => x"6f",
          9238 => x"63",
          9239 => x"74",
          9240 => x"00",
          9241 => x"2e",
          9242 => x"00",
          9243 => x"00",
          9244 => x"6c",
          9245 => x"74",
          9246 => x"6e",
          9247 => x"61",
          9248 => x"65",
          9249 => x"20",
          9250 => x"64",
          9251 => x"20",
          9252 => x"61",
          9253 => x"69",
          9254 => x"20",
          9255 => x"75",
          9256 => x"79",
          9257 => x"00",
          9258 => x"00",
          9259 => x"61",
          9260 => x"67",
          9261 => x"2e",
          9262 => x"00",
          9263 => x"79",
          9264 => x"2e",
          9265 => x"00",
          9266 => x"70",
          9267 => x"6e",
          9268 => x"2e",
          9269 => x"00",
          9270 => x"6c",
          9271 => x"30",
          9272 => x"2d",
          9273 => x"38",
          9274 => x"25",
          9275 => x"29",
          9276 => x"00",
          9277 => x"70",
          9278 => x"6d",
          9279 => x"0a",
          9280 => x"00",
          9281 => x"6d",
          9282 => x"74",
          9283 => x"00",
          9284 => x"58",
          9285 => x"32",
          9286 => x"00",
          9287 => x"0a",
          9288 => x"00",
          9289 => x"58",
          9290 => x"34",
          9291 => x"00",
          9292 => x"58",
          9293 => x"38",
          9294 => x"00",
          9295 => x"63",
          9296 => x"6e",
          9297 => x"6f",
          9298 => x"40",
          9299 => x"38",
          9300 => x"2e",
          9301 => x"00",
          9302 => x"6c",
          9303 => x"20",
          9304 => x"65",
          9305 => x"25",
          9306 => x"20",
          9307 => x"0a",
          9308 => x"00",
          9309 => x"6c",
          9310 => x"74",
          9311 => x"65",
          9312 => x"6f",
          9313 => x"28",
          9314 => x"2e",
          9315 => x"00",
          9316 => x"74",
          9317 => x"69",
          9318 => x"61",
          9319 => x"69",
          9320 => x"69",
          9321 => x"2e",
          9322 => x"00",
          9323 => x"64",
          9324 => x"62",
          9325 => x"69",
          9326 => x"2e",
          9327 => x"00",
          9328 => x"00",
          9329 => x"00",
          9330 => x"5c",
          9331 => x"25",
          9332 => x"73",
          9333 => x"00",
          9334 => x"5c",
          9335 => x"25",
          9336 => x"00",
          9337 => x"5c",
          9338 => x"00",
          9339 => x"20",
          9340 => x"6d",
          9341 => x"2e",
          9342 => x"00",
          9343 => x"4c",
          9344 => x"20",
          9345 => x"4d",
          9346 => x"49",
          9347 => x"00",
          9348 => x"4c",
          9349 => x"20",
          9350 => x"4d",
          9351 => x"49",
          9352 => x"00",
          9353 => x"6e",
          9354 => x"2e",
          9355 => x"00",
          9356 => x"62",
          9357 => x"67",
          9358 => x"74",
          9359 => x"75",
          9360 => x"2e",
          9361 => x"00",
          9362 => x"25",
          9363 => x"64",
          9364 => x"3a",
          9365 => x"25",
          9366 => x"64",
          9367 => x"00",
          9368 => x"20",
          9369 => x"66",
          9370 => x"72",
          9371 => x"6f",
          9372 => x"00",
          9373 => x"72",
          9374 => x"53",
          9375 => x"63",
          9376 => x"69",
          9377 => x"00",
          9378 => x"65",
          9379 => x"65",
          9380 => x"6d",
          9381 => x"6d",
          9382 => x"65",
          9383 => x"00",
          9384 => x"20",
          9385 => x"53",
          9386 => x"4d",
          9387 => x"25",
          9388 => x"3a",
          9389 => x"58",
          9390 => x"00",
          9391 => x"20",
          9392 => x"41",
          9393 => x"20",
          9394 => x"25",
          9395 => x"3a",
          9396 => x"58",
          9397 => x"00",
          9398 => x"20",
          9399 => x"4e",
          9400 => x"41",
          9401 => x"25",
          9402 => x"3a",
          9403 => x"58",
          9404 => x"00",
          9405 => x"20",
          9406 => x"4d",
          9407 => x"20",
          9408 => x"25",
          9409 => x"3a",
          9410 => x"58",
          9411 => x"00",
          9412 => x"20",
          9413 => x"20",
          9414 => x"20",
          9415 => x"25",
          9416 => x"3a",
          9417 => x"58",
          9418 => x"00",
          9419 => x"20",
          9420 => x"43",
          9421 => x"20",
          9422 => x"44",
          9423 => x"63",
          9424 => x"3d",
          9425 => x"64",
          9426 => x"00",
          9427 => x"20",
          9428 => x"45",
          9429 => x"20",
          9430 => x"54",
          9431 => x"72",
          9432 => x"3d",
          9433 => x"64",
          9434 => x"00",
          9435 => x"20",
          9436 => x"52",
          9437 => x"52",
          9438 => x"43",
          9439 => x"6e",
          9440 => x"3d",
          9441 => x"64",
          9442 => x"00",
          9443 => x"20",
          9444 => x"48",
          9445 => x"45",
          9446 => x"53",
          9447 => x"00",
          9448 => x"20",
          9449 => x"49",
          9450 => x"00",
          9451 => x"20",
          9452 => x"54",
          9453 => x"00",
          9454 => x"20",
          9455 => x"0a",
          9456 => x"00",
          9457 => x"20",
          9458 => x"0a",
          9459 => x"00",
          9460 => x"72",
          9461 => x"65",
          9462 => x"00",
          9463 => x"20",
          9464 => x"20",
          9465 => x"65",
          9466 => x"65",
          9467 => x"72",
          9468 => x"64",
          9469 => x"73",
          9470 => x"25",
          9471 => x"0a",
          9472 => x"00",
          9473 => x"20",
          9474 => x"20",
          9475 => x"6f",
          9476 => x"53",
          9477 => x"74",
          9478 => x"64",
          9479 => x"73",
          9480 => x"25",
          9481 => x"0a",
          9482 => x"00",
          9483 => x"20",
          9484 => x"63",
          9485 => x"74",
          9486 => x"20",
          9487 => x"72",
          9488 => x"20",
          9489 => x"20",
          9490 => x"25",
          9491 => x"0a",
          9492 => x"00",
          9493 => x"63",
          9494 => x"00",
          9495 => x"20",
          9496 => x"20",
          9497 => x"20",
          9498 => x"20",
          9499 => x"20",
          9500 => x"20",
          9501 => x"20",
          9502 => x"25",
          9503 => x"0a",
          9504 => x"00",
          9505 => x"20",
          9506 => x"74",
          9507 => x"43",
          9508 => x"6b",
          9509 => x"65",
          9510 => x"20",
          9511 => x"20",
          9512 => x"25",
          9513 => x"30",
          9514 => x"48",
          9515 => x"00",
          9516 => x"20",
          9517 => x"41",
          9518 => x"6c",
          9519 => x"20",
          9520 => x"71",
          9521 => x"20",
          9522 => x"20",
          9523 => x"25",
          9524 => x"30",
          9525 => x"48",
          9526 => x"00",
          9527 => x"20",
          9528 => x"68",
          9529 => x"65",
          9530 => x"52",
          9531 => x"43",
          9532 => x"6b",
          9533 => x"65",
          9534 => x"25",
          9535 => x"30",
          9536 => x"48",
          9537 => x"00",
          9538 => x"6c",
          9539 => x"00",
          9540 => x"69",
          9541 => x"00",
          9542 => x"78",
          9543 => x"00",
          9544 => x"00",
          9545 => x"6d",
          9546 => x"00",
          9547 => x"6e",
          9548 => x"00",
          9549 => x"90",
          9550 => x"00",
          9551 => x"02",
          9552 => x"8c",
          9553 => x"00",
          9554 => x"03",
          9555 => x"88",
          9556 => x"00",
          9557 => x"04",
          9558 => x"84",
          9559 => x"00",
          9560 => x"05",
          9561 => x"80",
          9562 => x"00",
          9563 => x"06",
          9564 => x"7c",
          9565 => x"00",
          9566 => x"07",
          9567 => x"78",
          9568 => x"00",
          9569 => x"01",
          9570 => x"74",
          9571 => x"00",
          9572 => x"08",
          9573 => x"70",
          9574 => x"00",
          9575 => x"0b",
          9576 => x"6c",
          9577 => x"00",
          9578 => x"09",
          9579 => x"68",
          9580 => x"00",
          9581 => x"0a",
          9582 => x"64",
          9583 => x"00",
          9584 => x"0d",
          9585 => x"60",
          9586 => x"00",
          9587 => x"0c",
          9588 => x"5c",
          9589 => x"00",
          9590 => x"0e",
          9591 => x"58",
          9592 => x"00",
          9593 => x"0f",
          9594 => x"54",
          9595 => x"00",
          9596 => x"0f",
          9597 => x"50",
          9598 => x"00",
          9599 => x"10",
          9600 => x"4c",
          9601 => x"00",
          9602 => x"11",
          9603 => x"48",
          9604 => x"00",
          9605 => x"12",
          9606 => x"44",
          9607 => x"00",
          9608 => x"13",
          9609 => x"40",
          9610 => x"00",
          9611 => x"14",
          9612 => x"3c",
          9613 => x"00",
          9614 => x"15",
          9615 => x"00",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"7e",
          9620 => x"7e",
          9621 => x"7e",
          9622 => x"00",
          9623 => x"7e",
          9624 => x"7e",
          9625 => x"7e",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"74",
          9638 => x"00",
          9639 => x"74",
          9640 => x"00",
          9641 => x"00",
          9642 => x"64",
          9643 => x"73",
          9644 => x"00",
          9645 => x"6c",
          9646 => x"74",
          9647 => x"65",
          9648 => x"20",
          9649 => x"20",
          9650 => x"74",
          9651 => x"20",
          9652 => x"65",
          9653 => x"20",
          9654 => x"2e",
          9655 => x"00",
          9656 => x"6e",
          9657 => x"6f",
          9658 => x"2f",
          9659 => x"61",
          9660 => x"68",
          9661 => x"6f",
          9662 => x"66",
          9663 => x"2c",
          9664 => x"73",
          9665 => x"69",
          9666 => x"00",
          9667 => x"00",
          9668 => x"2c",
          9669 => x"3d",
          9670 => x"5d",
          9671 => x"00",
          9672 => x"00",
          9673 => x"33",
          9674 => x"00",
          9675 => x"4d",
          9676 => x"53",
          9677 => x"00",
          9678 => x"4e",
          9679 => x"20",
          9680 => x"46",
          9681 => x"32",
          9682 => x"00",
          9683 => x"4e",
          9684 => x"20",
          9685 => x"46",
          9686 => x"20",
          9687 => x"00",
          9688 => x"0c",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"41",
          9693 => x"80",
          9694 => x"49",
          9695 => x"8f",
          9696 => x"4f",
          9697 => x"55",
          9698 => x"9b",
          9699 => x"9f",
          9700 => x"55",
          9701 => x"a7",
          9702 => x"ab",
          9703 => x"af",
          9704 => x"b3",
          9705 => x"b7",
          9706 => x"bb",
          9707 => x"bf",
          9708 => x"c3",
          9709 => x"c7",
          9710 => x"cb",
          9711 => x"cf",
          9712 => x"d3",
          9713 => x"d7",
          9714 => x"db",
          9715 => x"df",
          9716 => x"e3",
          9717 => x"e7",
          9718 => x"eb",
          9719 => x"ef",
          9720 => x"f3",
          9721 => x"f7",
          9722 => x"fb",
          9723 => x"ff",
          9724 => x"3b",
          9725 => x"2f",
          9726 => x"3a",
          9727 => x"7c",
          9728 => x"00",
          9729 => x"04",
          9730 => x"40",
          9731 => x"00",
          9732 => x"00",
          9733 => x"02",
          9734 => x"08",
          9735 => x"20",
          9736 => x"00",
          9737 => x"00",
          9738 => x"60",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"68",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"70",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"78",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"80",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"88",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"90",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"98",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"a0",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"a8",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"ac",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"b0",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"b4",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"b8",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"bc",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"c0",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"c4",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"cc",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"d0",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"d8",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"e0",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"e8",
          9823 => x"00",
          9824 => x"00",
          9825 => x"00",
          9826 => x"f0",
          9827 => x"00",
          9828 => x"00",
          9829 => x"00",
          9830 => x"f8",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"08",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"00",
          9844 => x"ff",
          9845 => x"00",
          9846 => x"ff",
          9847 => x"00",
          9848 => x"ff",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"ff",
          9853 => x"00",
          9854 => x"00",
          9855 => x"00",
          9856 => x"00",
          9857 => x"00",
          9858 => x"00",
          9859 => x"00",
          9860 => x"00",
          9861 => x"01",
          9862 => x"01",
          9863 => x"01",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"00",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"94",
          9890 => x"00",
          9891 => x"9c",
          9892 => x"00",
          9893 => x"a4",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b7",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"fe",
           279 => x"0b",
           280 => x"0b",
           281 => x"9c",
           282 => x"0b",
           283 => x"0b",
           284 => x"bb",
           285 => x"0b",
           286 => x"0b",
           287 => x"db",
           288 => x"0b",
           289 => x"0b",
           290 => x"fb",
           291 => x"0b",
           292 => x"0b",
           293 => x"9b",
           294 => x"0b",
           295 => x"0b",
           296 => x"bb",
           297 => x"0b",
           298 => x"0b",
           299 => x"db",
           300 => x"0b",
           301 => x"0b",
           302 => x"fb",
           303 => x"0b",
           304 => x"0b",
           305 => x"9b",
           306 => x"0b",
           307 => x"0b",
           308 => x"bb",
           309 => x"0b",
           310 => x"0b",
           311 => x"db",
           312 => x"0b",
           313 => x"0b",
           314 => x"fb",
           315 => x"0b",
           316 => x"0b",
           317 => x"9b",
           318 => x"0b",
           319 => x"0b",
           320 => x"bb",
           321 => x"0b",
           322 => x"0b",
           323 => x"db",
           324 => x"0b",
           325 => x"0b",
           326 => x"fb",
           327 => x"0b",
           328 => x"0b",
           329 => x"9b",
           330 => x"0b",
           331 => x"0b",
           332 => x"bb",
           333 => x"0b",
           334 => x"0b",
           335 => x"db",
           336 => x"0b",
           337 => x"0b",
           338 => x"fb",
           339 => x"0b",
           340 => x"0b",
           341 => x"9b",
           342 => x"0b",
           343 => x"0b",
           344 => x"bb",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"b5",
           386 => x"f4",
           387 => x"b5",
           388 => x"d0",
           389 => x"b5",
           390 => x"d2",
           391 => x"b4",
           392 => x"90",
           393 => x"b4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"82",
           400 => x"82",
           401 => x"94",
           402 => x"b5",
           403 => x"d0",
           404 => x"b5",
           405 => x"e2",
           406 => x"b4",
           407 => x"90",
           408 => x"b4",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"82",
           414 => x"82",
           415 => x"82",
           416 => x"93",
           417 => x"b5",
           418 => x"d0",
           419 => x"b5",
           420 => x"be",
           421 => x"b4",
           422 => x"90",
           423 => x"b4",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"2d",
           433 => x"08",
           434 => x"04",
           435 => x"0c",
           436 => x"2d",
           437 => x"08",
           438 => x"04",
           439 => x"0c",
           440 => x"2d",
           441 => x"08",
           442 => x"04",
           443 => x"0c",
           444 => x"2d",
           445 => x"08",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"04",
           451 => x"0c",
           452 => x"2d",
           453 => x"08",
           454 => x"04",
           455 => x"0c",
           456 => x"2d",
           457 => x"08",
           458 => x"04",
           459 => x"0c",
           460 => x"2d",
           461 => x"08",
           462 => x"04",
           463 => x"0c",
           464 => x"2d",
           465 => x"08",
           466 => x"04",
           467 => x"0c",
           468 => x"2d",
           469 => x"08",
           470 => x"04",
           471 => x"0c",
           472 => x"2d",
           473 => x"08",
           474 => x"04",
           475 => x"0c",
           476 => x"2d",
           477 => x"08",
           478 => x"04",
           479 => x"0c",
           480 => x"2d",
           481 => x"08",
           482 => x"04",
           483 => x"0c",
           484 => x"2d",
           485 => x"08",
           486 => x"04",
           487 => x"0c",
           488 => x"2d",
           489 => x"08",
           490 => x"04",
           491 => x"0c",
           492 => x"2d",
           493 => x"08",
           494 => x"04",
           495 => x"0c",
           496 => x"2d",
           497 => x"08",
           498 => x"04",
           499 => x"0c",
           500 => x"2d",
           501 => x"08",
           502 => x"04",
           503 => x"0c",
           504 => x"2d",
           505 => x"08",
           506 => x"04",
           507 => x"0c",
           508 => x"2d",
           509 => x"08",
           510 => x"04",
           511 => x"0c",
           512 => x"2d",
           513 => x"08",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"04",
           519 => x"0c",
           520 => x"2d",
           521 => x"08",
           522 => x"04",
           523 => x"0c",
           524 => x"2d",
           525 => x"08",
           526 => x"04",
           527 => x"0c",
           528 => x"2d",
           529 => x"08",
           530 => x"04",
           531 => x"0c",
           532 => x"2d",
           533 => x"08",
           534 => x"04",
           535 => x"0c",
           536 => x"2d",
           537 => x"08",
           538 => x"04",
           539 => x"0c",
           540 => x"2d",
           541 => x"08",
           542 => x"04",
           543 => x"0c",
           544 => x"2d",
           545 => x"08",
           546 => x"04",
           547 => x"0c",
           548 => x"2d",
           549 => x"08",
           550 => x"04",
           551 => x"0c",
           552 => x"2d",
           553 => x"08",
           554 => x"04",
           555 => x"0c",
           556 => x"2d",
           557 => x"08",
           558 => x"04",
           559 => x"0c",
           560 => x"2d",
           561 => x"08",
           562 => x"04",
           563 => x"0c",
           564 => x"2d",
           565 => x"08",
           566 => x"04",
           567 => x"0c",
           568 => x"2d",
           569 => x"08",
           570 => x"04",
           571 => x"0c",
           572 => x"2d",
           573 => x"08",
           574 => x"04",
           575 => x"0c",
           576 => x"2d",
           577 => x"08",
           578 => x"04",
           579 => x"0c",
           580 => x"2d",
           581 => x"08",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"04",
           587 => x"0c",
           588 => x"2d",
           589 => x"08",
           590 => x"04",
           591 => x"0c",
           592 => x"2d",
           593 => x"08",
           594 => x"04",
           595 => x"0c",
           596 => x"2d",
           597 => x"08",
           598 => x"04",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"53",
           608 => x"00",
           609 => x"06",
           610 => x"09",
           611 => x"05",
           612 => x"2b",
           613 => x"06",
           614 => x"04",
           615 => x"72",
           616 => x"05",
           617 => x"05",
           618 => x"72",
           619 => x"53",
           620 => x"51",
           621 => x"04",
           622 => x"70",
           623 => x"27",
           624 => x"71",
           625 => x"53",
           626 => x"0b",
           627 => x"8c",
           628 => x"ee",
           629 => x"82",
           630 => x"02",
           631 => x"0c",
           632 => x"82",
           633 => x"8c",
           634 => x"b5",
           635 => x"05",
           636 => x"b4",
           637 => x"08",
           638 => x"b4",
           639 => x"08",
           640 => x"fc",
           641 => x"84",
           642 => x"b5",
           643 => x"82",
           644 => x"f8",
           645 => x"b5",
           646 => x"05",
           647 => x"b5",
           648 => x"54",
           649 => x"82",
           650 => x"04",
           651 => x"08",
           652 => x"b4",
           653 => x"0d",
           654 => x"08",
           655 => x"85",
           656 => x"81",
           657 => x"06",
           658 => x"52",
           659 => x"80",
           660 => x"b4",
           661 => x"08",
           662 => x"8d",
           663 => x"82",
           664 => x"f4",
           665 => x"c4",
           666 => x"b4",
           667 => x"08",
           668 => x"b5",
           669 => x"05",
           670 => x"82",
           671 => x"f8",
           672 => x"b5",
           673 => x"05",
           674 => x"b4",
           675 => x"0c",
           676 => x"08",
           677 => x"8a",
           678 => x"38",
           679 => x"b5",
           680 => x"05",
           681 => x"e9",
           682 => x"b4",
           683 => x"08",
           684 => x"3f",
           685 => x"08",
           686 => x"b4",
           687 => x"0c",
           688 => x"b4",
           689 => x"08",
           690 => x"81",
           691 => x"80",
           692 => x"b4",
           693 => x"0c",
           694 => x"82",
           695 => x"fc",
           696 => x"b5",
           697 => x"05",
           698 => x"71",
           699 => x"b5",
           700 => x"05",
           701 => x"82",
           702 => x"8c",
           703 => x"b5",
           704 => x"05",
           705 => x"82",
           706 => x"fc",
           707 => x"80",
           708 => x"b4",
           709 => x"08",
           710 => x"34",
           711 => x"08",
           712 => x"70",
           713 => x"08",
           714 => x"52",
           715 => x"08",
           716 => x"82",
           717 => x"87",
           718 => x"b5",
           719 => x"82",
           720 => x"02",
           721 => x"0c",
           722 => x"86",
           723 => x"b4",
           724 => x"34",
           725 => x"08",
           726 => x"82",
           727 => x"e0",
           728 => x"0a",
           729 => x"b4",
           730 => x"0c",
           731 => x"08",
           732 => x"82",
           733 => x"fc",
           734 => x"b5",
           735 => x"05",
           736 => x"b5",
           737 => x"05",
           738 => x"b5",
           739 => x"05",
           740 => x"54",
           741 => x"82",
           742 => x"70",
           743 => x"08",
           744 => x"82",
           745 => x"ec",
           746 => x"b5",
           747 => x"05",
           748 => x"54",
           749 => x"82",
           750 => x"dc",
           751 => x"82",
           752 => x"54",
           753 => x"82",
           754 => x"04",
           755 => x"08",
           756 => x"b4",
           757 => x"0d",
           758 => x"08",
           759 => x"82",
           760 => x"fc",
           761 => x"b5",
           762 => x"05",
           763 => x"b5",
           764 => x"05",
           765 => x"b5",
           766 => x"05",
           767 => x"a3",
           768 => x"a8",
           769 => x"b5",
           770 => x"05",
           771 => x"b4",
           772 => x"08",
           773 => x"a8",
           774 => x"87",
           775 => x"b5",
           776 => x"82",
           777 => x"02",
           778 => x"0c",
           779 => x"80",
           780 => x"b4",
           781 => x"23",
           782 => x"08",
           783 => x"53",
           784 => x"14",
           785 => x"b4",
           786 => x"08",
           787 => x"70",
           788 => x"81",
           789 => x"06",
           790 => x"51",
           791 => x"2e",
           792 => x"0b",
           793 => x"08",
           794 => x"96",
           795 => x"b5",
           796 => x"05",
           797 => x"33",
           798 => x"b5",
           799 => x"05",
           800 => x"ff",
           801 => x"80",
           802 => x"38",
           803 => x"08",
           804 => x"81",
           805 => x"b4",
           806 => x"0c",
           807 => x"08",
           808 => x"70",
           809 => x"53",
           810 => x"95",
           811 => x"b5",
           812 => x"05",
           813 => x"73",
           814 => x"38",
           815 => x"08",
           816 => x"53",
           817 => x"81",
           818 => x"b5",
           819 => x"05",
           820 => x"b0",
           821 => x"06",
           822 => x"82",
           823 => x"e8",
           824 => x"98",
           825 => x"2c",
           826 => x"72",
           827 => x"b5",
           828 => x"05",
           829 => x"2a",
           830 => x"70",
           831 => x"51",
           832 => x"80",
           833 => x"82",
           834 => x"e4",
           835 => x"82",
           836 => x"53",
           837 => x"b4",
           838 => x"23",
           839 => x"82",
           840 => x"e8",
           841 => x"98",
           842 => x"2c",
           843 => x"2b",
           844 => x"11",
           845 => x"53",
           846 => x"72",
           847 => x"08",
           848 => x"82",
           849 => x"e8",
           850 => x"82",
           851 => x"f8",
           852 => x"15",
           853 => x"51",
           854 => x"b5",
           855 => x"05",
           856 => x"b4",
           857 => x"33",
           858 => x"70",
           859 => x"51",
           860 => x"25",
           861 => x"ff",
           862 => x"b4",
           863 => x"34",
           864 => x"08",
           865 => x"70",
           866 => x"81",
           867 => x"53",
           868 => x"38",
           869 => x"08",
           870 => x"70",
           871 => x"90",
           872 => x"2c",
           873 => x"51",
           874 => x"53",
           875 => x"b4",
           876 => x"23",
           877 => x"82",
           878 => x"e4",
           879 => x"83",
           880 => x"06",
           881 => x"72",
           882 => x"38",
           883 => x"08",
           884 => x"70",
           885 => x"98",
           886 => x"53",
           887 => x"81",
           888 => x"b4",
           889 => x"34",
           890 => x"08",
           891 => x"e0",
           892 => x"b4",
           893 => x"0c",
           894 => x"b4",
           895 => x"08",
           896 => x"92",
           897 => x"b5",
           898 => x"05",
           899 => x"2b",
           900 => x"11",
           901 => x"51",
           902 => x"04",
           903 => x"08",
           904 => x"70",
           905 => x"53",
           906 => x"b4",
           907 => x"23",
           908 => x"08",
           909 => x"70",
           910 => x"53",
           911 => x"b4",
           912 => x"23",
           913 => x"82",
           914 => x"e4",
           915 => x"81",
           916 => x"53",
           917 => x"b4",
           918 => x"23",
           919 => x"82",
           920 => x"e4",
           921 => x"80",
           922 => x"53",
           923 => x"b4",
           924 => x"23",
           925 => x"82",
           926 => x"e4",
           927 => x"88",
           928 => x"72",
           929 => x"08",
           930 => x"80",
           931 => x"b4",
           932 => x"34",
           933 => x"82",
           934 => x"e4",
           935 => x"84",
           936 => x"72",
           937 => x"08",
           938 => x"fb",
           939 => x"0b",
           940 => x"08",
           941 => x"82",
           942 => x"ec",
           943 => x"11",
           944 => x"82",
           945 => x"ec",
           946 => x"e3",
           947 => x"b4",
           948 => x"34",
           949 => x"82",
           950 => x"90",
           951 => x"b5",
           952 => x"05",
           953 => x"82",
           954 => x"90",
           955 => x"08",
           956 => x"82",
           957 => x"fc",
           958 => x"b5",
           959 => x"05",
           960 => x"51",
           961 => x"b5",
           962 => x"05",
           963 => x"39",
           964 => x"08",
           965 => x"82",
           966 => x"90",
           967 => x"05",
           968 => x"08",
           969 => x"70",
           970 => x"b4",
           971 => x"0c",
           972 => x"08",
           973 => x"70",
           974 => x"81",
           975 => x"51",
           976 => x"2e",
           977 => x"b5",
           978 => x"05",
           979 => x"2b",
           980 => x"2c",
           981 => x"b4",
           982 => x"08",
           983 => x"fa",
           984 => x"a8",
           985 => x"82",
           986 => x"f4",
           987 => x"39",
           988 => x"08",
           989 => x"51",
           990 => x"82",
           991 => x"53",
           992 => x"b4",
           993 => x"23",
           994 => x"08",
           995 => x"53",
           996 => x"08",
           997 => x"73",
           998 => x"54",
           999 => x"b4",
          1000 => x"23",
          1001 => x"82",
          1002 => x"90",
          1003 => x"b5",
          1004 => x"05",
          1005 => x"82",
          1006 => x"90",
          1007 => x"08",
          1008 => x"08",
          1009 => x"82",
          1010 => x"e4",
          1011 => x"83",
          1012 => x"06",
          1013 => x"53",
          1014 => x"ab",
          1015 => x"b4",
          1016 => x"33",
          1017 => x"53",
          1018 => x"53",
          1019 => x"08",
          1020 => x"52",
          1021 => x"3f",
          1022 => x"08",
          1023 => x"b5",
          1024 => x"05",
          1025 => x"82",
          1026 => x"fc",
          1027 => x"a7",
          1028 => x"b5",
          1029 => x"72",
          1030 => x"08",
          1031 => x"82",
          1032 => x"ec",
          1033 => x"82",
          1034 => x"f4",
          1035 => x"71",
          1036 => x"72",
          1037 => x"08",
          1038 => x"8a",
          1039 => x"b5",
          1040 => x"05",
          1041 => x"2a",
          1042 => x"51",
          1043 => x"80",
          1044 => x"82",
          1045 => x"90",
          1046 => x"b5",
          1047 => x"05",
          1048 => x"82",
          1049 => x"90",
          1050 => x"08",
          1051 => x"08",
          1052 => x"53",
          1053 => x"b5",
          1054 => x"05",
          1055 => x"b4",
          1056 => x"08",
          1057 => x"b5",
          1058 => x"05",
          1059 => x"82",
          1060 => x"dc",
          1061 => x"82",
          1062 => x"dc",
          1063 => x"b5",
          1064 => x"05",
          1065 => x"b4",
          1066 => x"08",
          1067 => x"38",
          1068 => x"08",
          1069 => x"70",
          1070 => x"53",
          1071 => x"b4",
          1072 => x"23",
          1073 => x"08",
          1074 => x"30",
          1075 => x"08",
          1076 => x"82",
          1077 => x"e4",
          1078 => x"ff",
          1079 => x"53",
          1080 => x"b4",
          1081 => x"23",
          1082 => x"88",
          1083 => x"b4",
          1084 => x"23",
          1085 => x"b5",
          1086 => x"05",
          1087 => x"c0",
          1088 => x"72",
          1089 => x"08",
          1090 => x"80",
          1091 => x"b5",
          1092 => x"05",
          1093 => x"82",
          1094 => x"f4",
          1095 => x"b5",
          1096 => x"05",
          1097 => x"2a",
          1098 => x"51",
          1099 => x"80",
          1100 => x"82",
          1101 => x"90",
          1102 => x"b5",
          1103 => x"05",
          1104 => x"82",
          1105 => x"90",
          1106 => x"08",
          1107 => x"08",
          1108 => x"53",
          1109 => x"b5",
          1110 => x"05",
          1111 => x"b4",
          1112 => x"08",
          1113 => x"b5",
          1114 => x"05",
          1115 => x"82",
          1116 => x"d8",
          1117 => x"82",
          1118 => x"d8",
          1119 => x"b5",
          1120 => x"05",
          1121 => x"b4",
          1122 => x"22",
          1123 => x"51",
          1124 => x"b5",
          1125 => x"05",
          1126 => x"b8",
          1127 => x"b4",
          1128 => x"0c",
          1129 => x"08",
          1130 => x"82",
          1131 => x"f4",
          1132 => x"b5",
          1133 => x"05",
          1134 => x"70",
          1135 => x"55",
          1136 => x"82",
          1137 => x"53",
          1138 => x"82",
          1139 => x"f0",
          1140 => x"b5",
          1141 => x"05",
          1142 => x"b4",
          1143 => x"08",
          1144 => x"53",
          1145 => x"a4",
          1146 => x"b4",
          1147 => x"08",
          1148 => x"54",
          1149 => x"08",
          1150 => x"70",
          1151 => x"51",
          1152 => x"82",
          1153 => x"d0",
          1154 => x"39",
          1155 => x"08",
          1156 => x"53",
          1157 => x"11",
          1158 => x"82",
          1159 => x"d0",
          1160 => x"b5",
          1161 => x"05",
          1162 => x"b5",
          1163 => x"05",
          1164 => x"82",
          1165 => x"f0",
          1166 => x"05",
          1167 => x"08",
          1168 => x"82",
          1169 => x"f4",
          1170 => x"53",
          1171 => x"08",
          1172 => x"52",
          1173 => x"3f",
          1174 => x"08",
          1175 => x"b4",
          1176 => x"0c",
          1177 => x"b4",
          1178 => x"08",
          1179 => x"38",
          1180 => x"82",
          1181 => x"f0",
          1182 => x"b5",
          1183 => x"72",
          1184 => x"75",
          1185 => x"72",
          1186 => x"08",
          1187 => x"82",
          1188 => x"e4",
          1189 => x"b2",
          1190 => x"72",
          1191 => x"38",
          1192 => x"08",
          1193 => x"ff",
          1194 => x"72",
          1195 => x"08",
          1196 => x"82",
          1197 => x"e4",
          1198 => x"86",
          1199 => x"06",
          1200 => x"72",
          1201 => x"e7",
          1202 => x"b4",
          1203 => x"22",
          1204 => x"82",
          1205 => x"cc",
          1206 => x"b5",
          1207 => x"05",
          1208 => x"82",
          1209 => x"cc",
          1210 => x"b5",
          1211 => x"05",
          1212 => x"72",
          1213 => x"81",
          1214 => x"82",
          1215 => x"cc",
          1216 => x"05",
          1217 => x"b5",
          1218 => x"05",
          1219 => x"82",
          1220 => x"cc",
          1221 => x"05",
          1222 => x"b5",
          1223 => x"05",
          1224 => x"b4",
          1225 => x"22",
          1226 => x"08",
          1227 => x"82",
          1228 => x"e4",
          1229 => x"83",
          1230 => x"06",
          1231 => x"72",
          1232 => x"d0",
          1233 => x"b4",
          1234 => x"33",
          1235 => x"70",
          1236 => x"b5",
          1237 => x"05",
          1238 => x"51",
          1239 => x"24",
          1240 => x"b5",
          1241 => x"05",
          1242 => x"06",
          1243 => x"82",
          1244 => x"e4",
          1245 => x"39",
          1246 => x"08",
          1247 => x"53",
          1248 => x"08",
          1249 => x"73",
          1250 => x"54",
          1251 => x"b4",
          1252 => x"34",
          1253 => x"08",
          1254 => x"70",
          1255 => x"81",
          1256 => x"53",
          1257 => x"b1",
          1258 => x"b4",
          1259 => x"33",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"82",
          1265 => x"ec",
          1266 => x"75",
          1267 => x"72",
          1268 => x"08",
          1269 => x"af",
          1270 => x"b4",
          1271 => x"33",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"82",
          1277 => x"ec",
          1278 => x"75",
          1279 => x"72",
          1280 => x"08",
          1281 => x"82",
          1282 => x"e4",
          1283 => x"83",
          1284 => x"53",
          1285 => x"82",
          1286 => x"ec",
          1287 => x"11",
          1288 => x"82",
          1289 => x"ec",
          1290 => x"90",
          1291 => x"2c",
          1292 => x"73",
          1293 => x"82",
          1294 => x"88",
          1295 => x"a0",
          1296 => x"3f",
          1297 => x"b5",
          1298 => x"05",
          1299 => x"2a",
          1300 => x"51",
          1301 => x"80",
          1302 => x"82",
          1303 => x"88",
          1304 => x"ad",
          1305 => x"3f",
          1306 => x"82",
          1307 => x"e4",
          1308 => x"84",
          1309 => x"06",
          1310 => x"72",
          1311 => x"38",
          1312 => x"08",
          1313 => x"52",
          1314 => x"c7",
          1315 => x"82",
          1316 => x"e4",
          1317 => x"85",
          1318 => x"06",
          1319 => x"72",
          1320 => x"38",
          1321 => x"08",
          1322 => x"52",
          1323 => x"a3",
          1324 => x"b4",
          1325 => x"22",
          1326 => x"70",
          1327 => x"51",
          1328 => x"2e",
          1329 => x"b5",
          1330 => x"05",
          1331 => x"51",
          1332 => x"82",
          1333 => x"f4",
          1334 => x"72",
          1335 => x"81",
          1336 => x"82",
          1337 => x"88",
          1338 => x"82",
          1339 => x"f8",
          1340 => x"94",
          1341 => x"b5",
          1342 => x"05",
          1343 => x"2a",
          1344 => x"51",
          1345 => x"80",
          1346 => x"82",
          1347 => x"ec",
          1348 => x"11",
          1349 => x"82",
          1350 => x"ec",
          1351 => x"90",
          1352 => x"2c",
          1353 => x"73",
          1354 => x"82",
          1355 => x"88",
          1356 => x"b0",
          1357 => x"3f",
          1358 => x"b5",
          1359 => x"05",
          1360 => x"2a",
          1361 => x"51",
          1362 => x"80",
          1363 => x"82",
          1364 => x"e8",
          1365 => x"11",
          1366 => x"82",
          1367 => x"e8",
          1368 => x"98",
          1369 => x"2c",
          1370 => x"73",
          1371 => x"82",
          1372 => x"88",
          1373 => x"b0",
          1374 => x"3f",
          1375 => x"b5",
          1376 => x"05",
          1377 => x"2a",
          1378 => x"51",
          1379 => x"b0",
          1380 => x"b4",
          1381 => x"22",
          1382 => x"54",
          1383 => x"b4",
          1384 => x"23",
          1385 => x"70",
          1386 => x"53",
          1387 => x"90",
          1388 => x"b4",
          1389 => x"08",
          1390 => x"93",
          1391 => x"39",
          1392 => x"08",
          1393 => x"53",
          1394 => x"2e",
          1395 => x"97",
          1396 => x"b4",
          1397 => x"08",
          1398 => x"b4",
          1399 => x"33",
          1400 => x"3f",
          1401 => x"82",
          1402 => x"f8",
          1403 => x"72",
          1404 => x"09",
          1405 => x"cb",
          1406 => x"b4",
          1407 => x"22",
          1408 => x"53",
          1409 => x"b4",
          1410 => x"23",
          1411 => x"ff",
          1412 => x"83",
          1413 => x"81",
          1414 => x"b5",
          1415 => x"05",
          1416 => x"b5",
          1417 => x"05",
          1418 => x"52",
          1419 => x"08",
          1420 => x"81",
          1421 => x"b4",
          1422 => x"0c",
          1423 => x"3f",
          1424 => x"82",
          1425 => x"f8",
          1426 => x"72",
          1427 => x"09",
          1428 => x"cb",
          1429 => x"b4",
          1430 => x"22",
          1431 => x"53",
          1432 => x"b4",
          1433 => x"23",
          1434 => x"ff",
          1435 => x"83",
          1436 => x"80",
          1437 => x"b5",
          1438 => x"05",
          1439 => x"b5",
          1440 => x"05",
          1441 => x"52",
          1442 => x"3f",
          1443 => x"08",
          1444 => x"81",
          1445 => x"b4",
          1446 => x"0c",
          1447 => x"82",
          1448 => x"f0",
          1449 => x"b5",
          1450 => x"38",
          1451 => x"08",
          1452 => x"52",
          1453 => x"08",
          1454 => x"ff",
          1455 => x"b4",
          1456 => x"0c",
          1457 => x"08",
          1458 => x"70",
          1459 => x"91",
          1460 => x"39",
          1461 => x"08",
          1462 => x"70",
          1463 => x"81",
          1464 => x"53",
          1465 => x"80",
          1466 => x"b5",
          1467 => x"05",
          1468 => x"54",
          1469 => x"b5",
          1470 => x"05",
          1471 => x"2b",
          1472 => x"51",
          1473 => x"25",
          1474 => x"b5",
          1475 => x"05",
          1476 => x"51",
          1477 => x"d2",
          1478 => x"b4",
          1479 => x"08",
          1480 => x"b4",
          1481 => x"33",
          1482 => x"3f",
          1483 => x"b5",
          1484 => x"05",
          1485 => x"39",
          1486 => x"08",
          1487 => x"53",
          1488 => x"09",
          1489 => x"38",
          1490 => x"b5",
          1491 => x"05",
          1492 => x"82",
          1493 => x"ec",
          1494 => x"0b",
          1495 => x"08",
          1496 => x"8a",
          1497 => x"b4",
          1498 => x"23",
          1499 => x"82",
          1500 => x"88",
          1501 => x"82",
          1502 => x"f8",
          1503 => x"8f",
          1504 => x"ea",
          1505 => x"b4",
          1506 => x"08",
          1507 => x"70",
          1508 => x"08",
          1509 => x"51",
          1510 => x"b4",
          1511 => x"08",
          1512 => x"0c",
          1513 => x"82",
          1514 => x"04",
          1515 => x"08",
          1516 => x"b4",
          1517 => x"0d",
          1518 => x"b5",
          1519 => x"05",
          1520 => x"b4",
          1521 => x"08",
          1522 => x"0c",
          1523 => x"08",
          1524 => x"70",
          1525 => x"72",
          1526 => x"82",
          1527 => x"f8",
          1528 => x"81",
          1529 => x"72",
          1530 => x"81",
          1531 => x"82",
          1532 => x"88",
          1533 => x"08",
          1534 => x"0c",
          1535 => x"82",
          1536 => x"f8",
          1537 => x"72",
          1538 => x"81",
          1539 => x"81",
          1540 => x"b4",
          1541 => x"34",
          1542 => x"08",
          1543 => x"70",
          1544 => x"71",
          1545 => x"51",
          1546 => x"82",
          1547 => x"f8",
          1548 => x"b5",
          1549 => x"05",
          1550 => x"b0",
          1551 => x"06",
          1552 => x"82",
          1553 => x"88",
          1554 => x"08",
          1555 => x"0c",
          1556 => x"53",
          1557 => x"b5",
          1558 => x"05",
          1559 => x"b4",
          1560 => x"33",
          1561 => x"08",
          1562 => x"82",
          1563 => x"e8",
          1564 => x"e2",
          1565 => x"82",
          1566 => x"e8",
          1567 => x"f8",
          1568 => x"80",
          1569 => x"0b",
          1570 => x"08",
          1571 => x"82",
          1572 => x"88",
          1573 => x"08",
          1574 => x"0c",
          1575 => x"53",
          1576 => x"b5",
          1577 => x"05",
          1578 => x"39",
          1579 => x"b5",
          1580 => x"05",
          1581 => x"b4",
          1582 => x"08",
          1583 => x"05",
          1584 => x"08",
          1585 => x"33",
          1586 => x"08",
          1587 => x"80",
          1588 => x"b5",
          1589 => x"05",
          1590 => x"a0",
          1591 => x"81",
          1592 => x"b4",
          1593 => x"0c",
          1594 => x"82",
          1595 => x"f8",
          1596 => x"af",
          1597 => x"38",
          1598 => x"08",
          1599 => x"53",
          1600 => x"83",
          1601 => x"80",
          1602 => x"b4",
          1603 => x"0c",
          1604 => x"88",
          1605 => x"b4",
          1606 => x"34",
          1607 => x"b5",
          1608 => x"05",
          1609 => x"73",
          1610 => x"82",
          1611 => x"f8",
          1612 => x"72",
          1613 => x"38",
          1614 => x"0b",
          1615 => x"08",
          1616 => x"82",
          1617 => x"0b",
          1618 => x"08",
          1619 => x"80",
          1620 => x"b4",
          1621 => x"0c",
          1622 => x"08",
          1623 => x"53",
          1624 => x"81",
          1625 => x"b5",
          1626 => x"05",
          1627 => x"e0",
          1628 => x"38",
          1629 => x"08",
          1630 => x"e0",
          1631 => x"72",
          1632 => x"08",
          1633 => x"82",
          1634 => x"f8",
          1635 => x"11",
          1636 => x"82",
          1637 => x"f8",
          1638 => x"b5",
          1639 => x"05",
          1640 => x"73",
          1641 => x"82",
          1642 => x"f8",
          1643 => x"11",
          1644 => x"82",
          1645 => x"f8",
          1646 => x"b5",
          1647 => x"05",
          1648 => x"89",
          1649 => x"80",
          1650 => x"b4",
          1651 => x"0c",
          1652 => x"82",
          1653 => x"f8",
          1654 => x"b5",
          1655 => x"05",
          1656 => x"72",
          1657 => x"38",
          1658 => x"b5",
          1659 => x"05",
          1660 => x"39",
          1661 => x"08",
          1662 => x"70",
          1663 => x"08",
          1664 => x"29",
          1665 => x"08",
          1666 => x"70",
          1667 => x"b4",
          1668 => x"0c",
          1669 => x"08",
          1670 => x"70",
          1671 => x"71",
          1672 => x"51",
          1673 => x"53",
          1674 => x"b5",
          1675 => x"05",
          1676 => x"39",
          1677 => x"08",
          1678 => x"53",
          1679 => x"90",
          1680 => x"b4",
          1681 => x"08",
          1682 => x"b4",
          1683 => x"0c",
          1684 => x"08",
          1685 => x"82",
          1686 => x"fc",
          1687 => x"0c",
          1688 => x"82",
          1689 => x"ec",
          1690 => x"b5",
          1691 => x"05",
          1692 => x"a8",
          1693 => x"0d",
          1694 => x"0c",
          1695 => x"b4",
          1696 => x"b5",
          1697 => x"3d",
          1698 => x"f8",
          1699 => x"b5",
          1700 => x"05",
          1701 => x"b5",
          1702 => x"05",
          1703 => x"8c",
          1704 => x"a8",
          1705 => x"b5",
          1706 => x"85",
          1707 => x"b5",
          1708 => x"82",
          1709 => x"02",
          1710 => x"0c",
          1711 => x"80",
          1712 => x"b4",
          1713 => x"34",
          1714 => x"08",
          1715 => x"53",
          1716 => x"82",
          1717 => x"88",
          1718 => x"08",
          1719 => x"33",
          1720 => x"b5",
          1721 => x"05",
          1722 => x"ff",
          1723 => x"a0",
          1724 => x"06",
          1725 => x"b5",
          1726 => x"05",
          1727 => x"81",
          1728 => x"53",
          1729 => x"b5",
          1730 => x"05",
          1731 => x"ad",
          1732 => x"06",
          1733 => x"0b",
          1734 => x"08",
          1735 => x"82",
          1736 => x"88",
          1737 => x"08",
          1738 => x"0c",
          1739 => x"53",
          1740 => x"b5",
          1741 => x"05",
          1742 => x"b4",
          1743 => x"33",
          1744 => x"2e",
          1745 => x"81",
          1746 => x"b5",
          1747 => x"05",
          1748 => x"81",
          1749 => x"70",
          1750 => x"72",
          1751 => x"b4",
          1752 => x"34",
          1753 => x"08",
          1754 => x"82",
          1755 => x"e8",
          1756 => x"b5",
          1757 => x"05",
          1758 => x"2e",
          1759 => x"b5",
          1760 => x"05",
          1761 => x"2e",
          1762 => x"cd",
          1763 => x"82",
          1764 => x"f4",
          1765 => x"b5",
          1766 => x"05",
          1767 => x"81",
          1768 => x"70",
          1769 => x"72",
          1770 => x"b4",
          1771 => x"34",
          1772 => x"82",
          1773 => x"b4",
          1774 => x"34",
          1775 => x"08",
          1776 => x"70",
          1777 => x"71",
          1778 => x"51",
          1779 => x"82",
          1780 => x"f8",
          1781 => x"fe",
          1782 => x"b4",
          1783 => x"33",
          1784 => x"26",
          1785 => x"0b",
          1786 => x"08",
          1787 => x"83",
          1788 => x"b5",
          1789 => x"05",
          1790 => x"73",
          1791 => x"82",
          1792 => x"f8",
          1793 => x"72",
          1794 => x"38",
          1795 => x"0b",
          1796 => x"08",
          1797 => x"82",
          1798 => x"0b",
          1799 => x"08",
          1800 => x"b2",
          1801 => x"b4",
          1802 => x"33",
          1803 => x"27",
          1804 => x"b5",
          1805 => x"05",
          1806 => x"b9",
          1807 => x"8d",
          1808 => x"82",
          1809 => x"ec",
          1810 => x"a5",
          1811 => x"82",
          1812 => x"f4",
          1813 => x"0b",
          1814 => x"08",
          1815 => x"82",
          1816 => x"f8",
          1817 => x"a0",
          1818 => x"cf",
          1819 => x"b4",
          1820 => x"33",
          1821 => x"73",
          1822 => x"82",
          1823 => x"f8",
          1824 => x"11",
          1825 => x"82",
          1826 => x"f8",
          1827 => x"b5",
          1828 => x"05",
          1829 => x"51",
          1830 => x"b5",
          1831 => x"05",
          1832 => x"b4",
          1833 => x"33",
          1834 => x"27",
          1835 => x"b5",
          1836 => x"05",
          1837 => x"51",
          1838 => x"b5",
          1839 => x"05",
          1840 => x"b4",
          1841 => x"33",
          1842 => x"26",
          1843 => x"0b",
          1844 => x"08",
          1845 => x"81",
          1846 => x"b5",
          1847 => x"05",
          1848 => x"b4",
          1849 => x"33",
          1850 => x"74",
          1851 => x"80",
          1852 => x"b4",
          1853 => x"0c",
          1854 => x"82",
          1855 => x"f4",
          1856 => x"82",
          1857 => x"fc",
          1858 => x"82",
          1859 => x"f8",
          1860 => x"12",
          1861 => x"08",
          1862 => x"82",
          1863 => x"88",
          1864 => x"08",
          1865 => x"0c",
          1866 => x"51",
          1867 => x"72",
          1868 => x"b4",
          1869 => x"34",
          1870 => x"82",
          1871 => x"f0",
          1872 => x"72",
          1873 => x"38",
          1874 => x"08",
          1875 => x"30",
          1876 => x"08",
          1877 => x"82",
          1878 => x"8c",
          1879 => x"b5",
          1880 => x"05",
          1881 => x"53",
          1882 => x"b5",
          1883 => x"05",
          1884 => x"b4",
          1885 => x"08",
          1886 => x"0c",
          1887 => x"82",
          1888 => x"04",
          1889 => x"08",
          1890 => x"b4",
          1891 => x"0d",
          1892 => x"b5",
          1893 => x"05",
          1894 => x"fc",
          1895 => x"33",
          1896 => x"70",
          1897 => x"81",
          1898 => x"51",
          1899 => x"80",
          1900 => x"ff",
          1901 => x"b4",
          1902 => x"0c",
          1903 => x"82",
          1904 => x"88",
          1905 => x"72",
          1906 => x"b4",
          1907 => x"08",
          1908 => x"b5",
          1909 => x"05",
          1910 => x"82",
          1911 => x"fc",
          1912 => x"81",
          1913 => x"72",
          1914 => x"38",
          1915 => x"08",
          1916 => x"08",
          1917 => x"b4",
          1918 => x"33",
          1919 => x"08",
          1920 => x"2d",
          1921 => x"08",
          1922 => x"2e",
          1923 => x"ff",
          1924 => x"b4",
          1925 => x"0c",
          1926 => x"82",
          1927 => x"82",
          1928 => x"53",
          1929 => x"90",
          1930 => x"72",
          1931 => x"a8",
          1932 => x"80",
          1933 => x"ff",
          1934 => x"b4",
          1935 => x"0c",
          1936 => x"08",
          1937 => x"70",
          1938 => x"08",
          1939 => x"53",
          1940 => x"08",
          1941 => x"82",
          1942 => x"87",
          1943 => x"b5",
          1944 => x"82",
          1945 => x"02",
          1946 => x"0c",
          1947 => x"80",
          1948 => x"b4",
          1949 => x"0c",
          1950 => x"08",
          1951 => x"85",
          1952 => x"81",
          1953 => x"32",
          1954 => x"51",
          1955 => x"53",
          1956 => x"8d",
          1957 => x"82",
          1958 => x"f4",
          1959 => x"f3",
          1960 => x"b4",
          1961 => x"08",
          1962 => x"82",
          1963 => x"88",
          1964 => x"05",
          1965 => x"08",
          1966 => x"53",
          1967 => x"b4",
          1968 => x"34",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"b5",
          1972 => x"05",
          1973 => x"b4",
          1974 => x"08",
          1975 => x"b4",
          1976 => x"33",
          1977 => x"08",
          1978 => x"2d",
          1979 => x"08",
          1980 => x"2e",
          1981 => x"ff",
          1982 => x"b4",
          1983 => x"0c",
          1984 => x"82",
          1985 => x"f8",
          1986 => x"82",
          1987 => x"f4",
          1988 => x"82",
          1989 => x"f4",
          1990 => x"b5",
          1991 => x"3d",
          1992 => x"b4",
          1993 => x"b5",
          1994 => x"82",
          1995 => x"fe",
          1996 => x"cc",
          1997 => x"82",
          1998 => x"88",
          1999 => x"93",
          2000 => x"a8",
          2001 => x"b5",
          2002 => x"84",
          2003 => x"b5",
          2004 => x"82",
          2005 => x"02",
          2006 => x"0c",
          2007 => x"82",
          2008 => x"8c",
          2009 => x"11",
          2010 => x"2a",
          2011 => x"70",
          2012 => x"51",
          2013 => x"72",
          2014 => x"38",
          2015 => x"b5",
          2016 => x"05",
          2017 => x"39",
          2018 => x"08",
          2019 => x"85",
          2020 => x"82",
          2021 => x"06",
          2022 => x"53",
          2023 => x"80",
          2024 => x"b5",
          2025 => x"05",
          2026 => x"b4",
          2027 => x"08",
          2028 => x"14",
          2029 => x"08",
          2030 => x"82",
          2031 => x"8c",
          2032 => x"08",
          2033 => x"b4",
          2034 => x"08",
          2035 => x"54",
          2036 => x"73",
          2037 => x"74",
          2038 => x"b4",
          2039 => x"08",
          2040 => x"81",
          2041 => x"0c",
          2042 => x"08",
          2043 => x"70",
          2044 => x"08",
          2045 => x"51",
          2046 => x"39",
          2047 => x"08",
          2048 => x"82",
          2049 => x"8c",
          2050 => x"82",
          2051 => x"88",
          2052 => x"81",
          2053 => x"90",
          2054 => x"54",
          2055 => x"82",
          2056 => x"53",
          2057 => x"82",
          2058 => x"8c",
          2059 => x"11",
          2060 => x"8c",
          2061 => x"b5",
          2062 => x"05",
          2063 => x"b5",
          2064 => x"05",
          2065 => x"8a",
          2066 => x"82",
          2067 => x"fc",
          2068 => x"b5",
          2069 => x"05",
          2070 => x"a8",
          2071 => x"0d",
          2072 => x"0c",
          2073 => x"b4",
          2074 => x"b5",
          2075 => x"3d",
          2076 => x"b4",
          2077 => x"08",
          2078 => x"70",
          2079 => x"81",
          2080 => x"51",
          2081 => x"2e",
          2082 => x"0b",
          2083 => x"08",
          2084 => x"83",
          2085 => x"b5",
          2086 => x"05",
          2087 => x"33",
          2088 => x"70",
          2089 => x"51",
          2090 => x"80",
          2091 => x"38",
          2092 => x"08",
          2093 => x"82",
          2094 => x"88",
          2095 => x"53",
          2096 => x"70",
          2097 => x"51",
          2098 => x"14",
          2099 => x"b4",
          2100 => x"08",
          2101 => x"81",
          2102 => x"0c",
          2103 => x"08",
          2104 => x"84",
          2105 => x"82",
          2106 => x"f8",
          2107 => x"51",
          2108 => x"39",
          2109 => x"08",
          2110 => x"85",
          2111 => x"82",
          2112 => x"06",
          2113 => x"52",
          2114 => x"80",
          2115 => x"b5",
          2116 => x"05",
          2117 => x"70",
          2118 => x"b4",
          2119 => x"0c",
          2120 => x"b5",
          2121 => x"05",
          2122 => x"82",
          2123 => x"88",
          2124 => x"b5",
          2125 => x"05",
          2126 => x"85",
          2127 => x"a0",
          2128 => x"71",
          2129 => x"ff",
          2130 => x"b4",
          2131 => x"0c",
          2132 => x"82",
          2133 => x"88",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"39",
          2137 => x"08",
          2138 => x"82",
          2139 => x"88",
          2140 => x"94",
          2141 => x"52",
          2142 => x"b5",
          2143 => x"82",
          2144 => x"fc",
          2145 => x"82",
          2146 => x"fc",
          2147 => x"25",
          2148 => x"82",
          2149 => x"88",
          2150 => x"b5",
          2151 => x"05",
          2152 => x"b4",
          2153 => x"08",
          2154 => x"82",
          2155 => x"f0",
          2156 => x"82",
          2157 => x"fc",
          2158 => x"2e",
          2159 => x"95",
          2160 => x"b4",
          2161 => x"08",
          2162 => x"71",
          2163 => x"08",
          2164 => x"93",
          2165 => x"b4",
          2166 => x"08",
          2167 => x"71",
          2168 => x"08",
          2169 => x"82",
          2170 => x"f4",
          2171 => x"82",
          2172 => x"ec",
          2173 => x"13",
          2174 => x"82",
          2175 => x"f8",
          2176 => x"39",
          2177 => x"08",
          2178 => x"8c",
          2179 => x"05",
          2180 => x"82",
          2181 => x"fc",
          2182 => x"81",
          2183 => x"82",
          2184 => x"f8",
          2185 => x"51",
          2186 => x"b4",
          2187 => x"08",
          2188 => x"0c",
          2189 => x"82",
          2190 => x"04",
          2191 => x"08",
          2192 => x"b4",
          2193 => x"0d",
          2194 => x"08",
          2195 => x"82",
          2196 => x"fc",
          2197 => x"b5",
          2198 => x"05",
          2199 => x"b4",
          2200 => x"0c",
          2201 => x"08",
          2202 => x"80",
          2203 => x"38",
          2204 => x"08",
          2205 => x"82",
          2206 => x"fc",
          2207 => x"81",
          2208 => x"b5",
          2209 => x"05",
          2210 => x"b4",
          2211 => x"08",
          2212 => x"b5",
          2213 => x"05",
          2214 => x"81",
          2215 => x"b5",
          2216 => x"05",
          2217 => x"b4",
          2218 => x"08",
          2219 => x"b4",
          2220 => x"0c",
          2221 => x"08",
          2222 => x"82",
          2223 => x"90",
          2224 => x"82",
          2225 => x"f8",
          2226 => x"b5",
          2227 => x"05",
          2228 => x"82",
          2229 => x"90",
          2230 => x"b5",
          2231 => x"05",
          2232 => x"82",
          2233 => x"90",
          2234 => x"b5",
          2235 => x"05",
          2236 => x"81",
          2237 => x"b5",
          2238 => x"05",
          2239 => x"82",
          2240 => x"fc",
          2241 => x"b5",
          2242 => x"05",
          2243 => x"82",
          2244 => x"f8",
          2245 => x"b5",
          2246 => x"05",
          2247 => x"b4",
          2248 => x"08",
          2249 => x"33",
          2250 => x"ae",
          2251 => x"b4",
          2252 => x"08",
          2253 => x"b5",
          2254 => x"05",
          2255 => x"b4",
          2256 => x"08",
          2257 => x"b5",
          2258 => x"05",
          2259 => x"b4",
          2260 => x"08",
          2261 => x"38",
          2262 => x"08",
          2263 => x"51",
          2264 => x"b5",
          2265 => x"05",
          2266 => x"82",
          2267 => x"f8",
          2268 => x"b5",
          2269 => x"05",
          2270 => x"71",
          2271 => x"b5",
          2272 => x"05",
          2273 => x"82",
          2274 => x"fc",
          2275 => x"ad",
          2276 => x"b4",
          2277 => x"08",
          2278 => x"a8",
          2279 => x"3d",
          2280 => x"b4",
          2281 => x"b5",
          2282 => x"82",
          2283 => x"fe",
          2284 => x"b5",
          2285 => x"05",
          2286 => x"b4",
          2287 => x"0c",
          2288 => x"08",
          2289 => x"52",
          2290 => x"b5",
          2291 => x"05",
          2292 => x"82",
          2293 => x"fc",
          2294 => x"81",
          2295 => x"51",
          2296 => x"83",
          2297 => x"82",
          2298 => x"fc",
          2299 => x"05",
          2300 => x"08",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"b5",
          2304 => x"05",
          2305 => x"82",
          2306 => x"51",
          2307 => x"82",
          2308 => x"04",
          2309 => x"08",
          2310 => x"b4",
          2311 => x"0d",
          2312 => x"08",
          2313 => x"82",
          2314 => x"fc",
          2315 => x"b5",
          2316 => x"05",
          2317 => x"33",
          2318 => x"08",
          2319 => x"81",
          2320 => x"b4",
          2321 => x"0c",
          2322 => x"08",
          2323 => x"53",
          2324 => x"34",
          2325 => x"08",
          2326 => x"81",
          2327 => x"b4",
          2328 => x"0c",
          2329 => x"06",
          2330 => x"2e",
          2331 => x"be",
          2332 => x"b4",
          2333 => x"08",
          2334 => x"a8",
          2335 => x"3d",
          2336 => x"b4",
          2337 => x"b5",
          2338 => x"82",
          2339 => x"fd",
          2340 => x"b5",
          2341 => x"05",
          2342 => x"b4",
          2343 => x"0c",
          2344 => x"08",
          2345 => x"82",
          2346 => x"f8",
          2347 => x"b5",
          2348 => x"05",
          2349 => x"80",
          2350 => x"b5",
          2351 => x"05",
          2352 => x"82",
          2353 => x"90",
          2354 => x"b5",
          2355 => x"05",
          2356 => x"82",
          2357 => x"90",
          2358 => x"b5",
          2359 => x"05",
          2360 => x"ba",
          2361 => x"b4",
          2362 => x"08",
          2363 => x"82",
          2364 => x"f8",
          2365 => x"05",
          2366 => x"08",
          2367 => x"82",
          2368 => x"fc",
          2369 => x"52",
          2370 => x"82",
          2371 => x"fc",
          2372 => x"05",
          2373 => x"08",
          2374 => x"ff",
          2375 => x"b5",
          2376 => x"05",
          2377 => x"b5",
          2378 => x"85",
          2379 => x"b5",
          2380 => x"82",
          2381 => x"02",
          2382 => x"0c",
          2383 => x"82",
          2384 => x"90",
          2385 => x"2e",
          2386 => x"82",
          2387 => x"8c",
          2388 => x"71",
          2389 => x"b4",
          2390 => x"08",
          2391 => x"b5",
          2392 => x"05",
          2393 => x"b4",
          2394 => x"08",
          2395 => x"81",
          2396 => x"54",
          2397 => x"71",
          2398 => x"80",
          2399 => x"b5",
          2400 => x"05",
          2401 => x"33",
          2402 => x"08",
          2403 => x"81",
          2404 => x"b4",
          2405 => x"0c",
          2406 => x"06",
          2407 => x"8d",
          2408 => x"82",
          2409 => x"fc",
          2410 => x"9b",
          2411 => x"b4",
          2412 => x"08",
          2413 => x"b5",
          2414 => x"05",
          2415 => x"b4",
          2416 => x"08",
          2417 => x"38",
          2418 => x"82",
          2419 => x"90",
          2420 => x"2e",
          2421 => x"82",
          2422 => x"88",
          2423 => x"33",
          2424 => x"8d",
          2425 => x"82",
          2426 => x"fc",
          2427 => x"d7",
          2428 => x"b4",
          2429 => x"08",
          2430 => x"b5",
          2431 => x"05",
          2432 => x"b4",
          2433 => x"08",
          2434 => x"52",
          2435 => x"81",
          2436 => x"b4",
          2437 => x"0c",
          2438 => x"b5",
          2439 => x"05",
          2440 => x"82",
          2441 => x"8c",
          2442 => x"33",
          2443 => x"70",
          2444 => x"08",
          2445 => x"53",
          2446 => x"53",
          2447 => x"0b",
          2448 => x"08",
          2449 => x"82",
          2450 => x"fc",
          2451 => x"b5",
          2452 => x"3d",
          2453 => x"b4",
          2454 => x"b5",
          2455 => x"82",
          2456 => x"fd",
          2457 => x"b5",
          2458 => x"05",
          2459 => x"b4",
          2460 => x"0c",
          2461 => x"08",
          2462 => x"8d",
          2463 => x"82",
          2464 => x"fc",
          2465 => x"ec",
          2466 => x"b4",
          2467 => x"08",
          2468 => x"82",
          2469 => x"f8",
          2470 => x"05",
          2471 => x"08",
          2472 => x"70",
          2473 => x"51",
          2474 => x"2e",
          2475 => x"b5",
          2476 => x"05",
          2477 => x"82",
          2478 => x"8c",
          2479 => x"b5",
          2480 => x"05",
          2481 => x"84",
          2482 => x"39",
          2483 => x"08",
          2484 => x"ff",
          2485 => x"b4",
          2486 => x"0c",
          2487 => x"08",
          2488 => x"82",
          2489 => x"88",
          2490 => x"70",
          2491 => x"08",
          2492 => x"51",
          2493 => x"08",
          2494 => x"82",
          2495 => x"85",
          2496 => x"b5",
          2497 => x"82",
          2498 => x"02",
          2499 => x"0c",
          2500 => x"82",
          2501 => x"88",
          2502 => x"b5",
          2503 => x"05",
          2504 => x"b4",
          2505 => x"08",
          2506 => x"d4",
          2507 => x"b4",
          2508 => x"08",
          2509 => x"b5",
          2510 => x"05",
          2511 => x"b4",
          2512 => x"08",
          2513 => x"b5",
          2514 => x"05",
          2515 => x"b4",
          2516 => x"08",
          2517 => x"38",
          2518 => x"08",
          2519 => x"51",
          2520 => x"b4",
          2521 => x"08",
          2522 => x"71",
          2523 => x"b4",
          2524 => x"08",
          2525 => x"b5",
          2526 => x"05",
          2527 => x"39",
          2528 => x"08",
          2529 => x"70",
          2530 => x"0c",
          2531 => x"0d",
          2532 => x"0c",
          2533 => x"b4",
          2534 => x"b5",
          2535 => x"3d",
          2536 => x"82",
          2537 => x"fc",
          2538 => x"b5",
          2539 => x"05",
          2540 => x"b9",
          2541 => x"b4",
          2542 => x"08",
          2543 => x"b4",
          2544 => x"0c",
          2545 => x"b5",
          2546 => x"05",
          2547 => x"b4",
          2548 => x"08",
          2549 => x"0b",
          2550 => x"08",
          2551 => x"82",
          2552 => x"f4",
          2553 => x"b5",
          2554 => x"05",
          2555 => x"b4",
          2556 => x"08",
          2557 => x"38",
          2558 => x"08",
          2559 => x"30",
          2560 => x"08",
          2561 => x"80",
          2562 => x"b4",
          2563 => x"0c",
          2564 => x"08",
          2565 => x"8a",
          2566 => x"82",
          2567 => x"f0",
          2568 => x"b5",
          2569 => x"05",
          2570 => x"b4",
          2571 => x"0c",
          2572 => x"b5",
          2573 => x"05",
          2574 => x"b5",
          2575 => x"05",
          2576 => x"c5",
          2577 => x"a8",
          2578 => x"b5",
          2579 => x"05",
          2580 => x"b5",
          2581 => x"05",
          2582 => x"90",
          2583 => x"b4",
          2584 => x"08",
          2585 => x"b4",
          2586 => x"0c",
          2587 => x"08",
          2588 => x"70",
          2589 => x"0c",
          2590 => x"0d",
          2591 => x"0c",
          2592 => x"b4",
          2593 => x"b5",
          2594 => x"3d",
          2595 => x"82",
          2596 => x"fc",
          2597 => x"b5",
          2598 => x"05",
          2599 => x"99",
          2600 => x"b4",
          2601 => x"08",
          2602 => x"b4",
          2603 => x"0c",
          2604 => x"b5",
          2605 => x"05",
          2606 => x"b4",
          2607 => x"08",
          2608 => x"38",
          2609 => x"08",
          2610 => x"30",
          2611 => x"08",
          2612 => x"81",
          2613 => x"b4",
          2614 => x"08",
          2615 => x"b4",
          2616 => x"08",
          2617 => x"3f",
          2618 => x"08",
          2619 => x"b4",
          2620 => x"0c",
          2621 => x"b4",
          2622 => x"08",
          2623 => x"38",
          2624 => x"08",
          2625 => x"30",
          2626 => x"08",
          2627 => x"82",
          2628 => x"f8",
          2629 => x"82",
          2630 => x"54",
          2631 => x"82",
          2632 => x"04",
          2633 => x"08",
          2634 => x"b4",
          2635 => x"0d",
          2636 => x"b5",
          2637 => x"05",
          2638 => x"b5",
          2639 => x"05",
          2640 => x"c5",
          2641 => x"a8",
          2642 => x"b5",
          2643 => x"85",
          2644 => x"b5",
          2645 => x"82",
          2646 => x"02",
          2647 => x"0c",
          2648 => x"81",
          2649 => x"b4",
          2650 => x"08",
          2651 => x"b4",
          2652 => x"08",
          2653 => x"82",
          2654 => x"70",
          2655 => x"0c",
          2656 => x"0d",
          2657 => x"0c",
          2658 => x"b4",
          2659 => x"b5",
          2660 => x"3d",
          2661 => x"82",
          2662 => x"fc",
          2663 => x"0b",
          2664 => x"08",
          2665 => x"82",
          2666 => x"8c",
          2667 => x"b5",
          2668 => x"05",
          2669 => x"38",
          2670 => x"08",
          2671 => x"80",
          2672 => x"80",
          2673 => x"b4",
          2674 => x"08",
          2675 => x"82",
          2676 => x"8c",
          2677 => x"82",
          2678 => x"8c",
          2679 => x"b5",
          2680 => x"05",
          2681 => x"b5",
          2682 => x"05",
          2683 => x"39",
          2684 => x"08",
          2685 => x"80",
          2686 => x"38",
          2687 => x"08",
          2688 => x"82",
          2689 => x"88",
          2690 => x"ad",
          2691 => x"b4",
          2692 => x"08",
          2693 => x"08",
          2694 => x"31",
          2695 => x"08",
          2696 => x"82",
          2697 => x"f8",
          2698 => x"b5",
          2699 => x"05",
          2700 => x"b5",
          2701 => x"05",
          2702 => x"b4",
          2703 => x"08",
          2704 => x"b5",
          2705 => x"05",
          2706 => x"b4",
          2707 => x"08",
          2708 => x"b5",
          2709 => x"05",
          2710 => x"39",
          2711 => x"08",
          2712 => x"80",
          2713 => x"82",
          2714 => x"88",
          2715 => x"82",
          2716 => x"f4",
          2717 => x"91",
          2718 => x"b4",
          2719 => x"08",
          2720 => x"b4",
          2721 => x"0c",
          2722 => x"b4",
          2723 => x"08",
          2724 => x"0c",
          2725 => x"82",
          2726 => x"04",
          2727 => x"79",
          2728 => x"56",
          2729 => x"80",
          2730 => x"38",
          2731 => x"08",
          2732 => x"3f",
          2733 => x"08",
          2734 => x"85",
          2735 => x"80",
          2736 => x"33",
          2737 => x"2e",
          2738 => x"86",
          2739 => x"55",
          2740 => x"57",
          2741 => x"82",
          2742 => x"70",
          2743 => x"f1",
          2744 => x"b5",
          2745 => x"74",
          2746 => x"51",
          2747 => x"82",
          2748 => x"8b",
          2749 => x"33",
          2750 => x"2e",
          2751 => x"81",
          2752 => x"ff",
          2753 => x"99",
          2754 => x"38",
          2755 => x"82",
          2756 => x"89",
          2757 => x"ff",
          2758 => x"52",
          2759 => x"81",
          2760 => x"84",
          2761 => x"c0",
          2762 => x"08",
          2763 => x"8c",
          2764 => x"39",
          2765 => x"51",
          2766 => x"82",
          2767 => x"80",
          2768 => x"9a",
          2769 => x"eb",
          2770 => x"d0",
          2771 => x"39",
          2772 => x"51",
          2773 => x"82",
          2774 => x"80",
          2775 => x"9b",
          2776 => x"cf",
          2777 => x"9c",
          2778 => x"39",
          2779 => x"51",
          2780 => x"82",
          2781 => x"bb",
          2782 => x"e8",
          2783 => x"82",
          2784 => x"af",
          2785 => x"a8",
          2786 => x"82",
          2787 => x"a3",
          2788 => x"dc",
          2789 => x"82",
          2790 => x"97",
          2791 => x"88",
          2792 => x"82",
          2793 => x"8b",
          2794 => x"b8",
          2795 => x"82",
          2796 => x"e3",
          2797 => x"3d",
          2798 => x"3d",
          2799 => x"56",
          2800 => x"e7",
          2801 => x"74",
          2802 => x"e8",
          2803 => x"39",
          2804 => x"74",
          2805 => x"3f",
          2806 => x"08",
          2807 => x"fa",
          2808 => x"b5",
          2809 => x"79",
          2810 => x"82",
          2811 => x"ff",
          2812 => x"87",
          2813 => x"ec",
          2814 => x"02",
          2815 => x"e3",
          2816 => x"57",
          2817 => x"30",
          2818 => x"73",
          2819 => x"59",
          2820 => x"77",
          2821 => x"83",
          2822 => x"74",
          2823 => x"81",
          2824 => x"55",
          2825 => x"81",
          2826 => x"53",
          2827 => x"3d",
          2828 => x"80",
          2829 => x"82",
          2830 => x"57",
          2831 => x"08",
          2832 => x"b5",
          2833 => x"c0",
          2834 => x"82",
          2835 => x"59",
          2836 => x"05",
          2837 => x"53",
          2838 => x"51",
          2839 => x"3f",
          2840 => x"08",
          2841 => x"a8",
          2842 => x"7a",
          2843 => x"2e",
          2844 => x"19",
          2845 => x"59",
          2846 => x"3d",
          2847 => x"81",
          2848 => x"76",
          2849 => x"07",
          2850 => x"30",
          2851 => x"72",
          2852 => x"51",
          2853 => x"2e",
          2854 => x"9d",
          2855 => x"c0",
          2856 => x"52",
          2857 => x"92",
          2858 => x"75",
          2859 => x"0c",
          2860 => x"04",
          2861 => x"7c",
          2862 => x"b7",
          2863 => x"59",
          2864 => x"53",
          2865 => x"51",
          2866 => x"82",
          2867 => x"a6",
          2868 => x"2e",
          2869 => x"81",
          2870 => x"9a",
          2871 => x"61",
          2872 => x"82",
          2873 => x"7f",
          2874 => x"78",
          2875 => x"a8",
          2876 => x"39",
          2877 => x"82",
          2878 => x"8a",
          2879 => x"f3",
          2880 => x"61",
          2881 => x"05",
          2882 => x"33",
          2883 => x"68",
          2884 => x"5c",
          2885 => x"7a",
          2886 => x"80",
          2887 => x"b7",
          2888 => x"88",
          2889 => x"3f",
          2890 => x"79",
          2891 => x"38",
          2892 => x"89",
          2893 => x"2e",
          2894 => x"c4",
          2895 => x"53",
          2896 => x"8e",
          2897 => x"52",
          2898 => x"51",
          2899 => x"3f",
          2900 => x"9e",
          2901 => x"ac",
          2902 => x"55",
          2903 => x"74",
          2904 => x"7a",
          2905 => x"72",
          2906 => x"9e",
          2907 => x"b8",
          2908 => x"39",
          2909 => x"51",
          2910 => x"84",
          2911 => x"39",
          2912 => x"72",
          2913 => x"38",
          2914 => x"82",
          2915 => x"ff",
          2916 => x"88",
          2917 => x"a8",
          2918 => x"3f",
          2919 => x"82",
          2920 => x"52",
          2921 => x"ab",
          2922 => x"39",
          2923 => x"51",
          2924 => x"80",
          2925 => x"27",
          2926 => x"74",
          2927 => x"55",
          2928 => x"72",
          2929 => x"38",
          2930 => x"53",
          2931 => x"83",
          2932 => x"75",
          2933 => x"81",
          2934 => x"53",
          2935 => x"90",
          2936 => x"fe",
          2937 => x"82",
          2938 => x"52",
          2939 => x"39",
          2940 => x"08",
          2941 => x"e2",
          2942 => x"15",
          2943 => x"39",
          2944 => x"51",
          2945 => x"78",
          2946 => x"5c",
          2947 => x"3f",
          2948 => x"08",
          2949 => x"98",
          2950 => x"76",
          2951 => x"81",
          2952 => x"9c",
          2953 => x"b5",
          2954 => x"2b",
          2955 => x"70",
          2956 => x"30",
          2957 => x"70",
          2958 => x"07",
          2959 => x"06",
          2960 => x"59",
          2961 => x"80",
          2962 => x"38",
          2963 => x"09",
          2964 => x"38",
          2965 => x"39",
          2966 => x"72",
          2967 => x"b7",
          2968 => x"72",
          2969 => x"0c",
          2970 => x"04",
          2971 => x"02",
          2972 => x"82",
          2973 => x"82",
          2974 => x"55",
          2975 => x"3f",
          2976 => x"22",
          2977 => x"3f",
          2978 => x"54",
          2979 => x"53",
          2980 => x"33",
          2981 => x"d8",
          2982 => x"bb",
          2983 => x"2e",
          2984 => x"cd",
          2985 => x"0d",
          2986 => x"0d",
          2987 => x"80",
          2988 => x"b7",
          2989 => x"98",
          2990 => x"9e",
          2991 => x"98",
          2992 => x"97",
          2993 => x"81",
          2994 => x"06",
          2995 => x"80",
          2996 => x"81",
          2997 => x"3f",
          2998 => x"51",
          2999 => x"80",
          3000 => x"3f",
          3001 => x"70",
          3002 => x"52",
          3003 => x"92",
          3004 => x"97",
          3005 => x"9f",
          3006 => x"dc",
          3007 => x"97",
          3008 => x"83",
          3009 => x"06",
          3010 => x"80",
          3011 => x"81",
          3012 => x"3f",
          3013 => x"51",
          3014 => x"80",
          3015 => x"3f",
          3016 => x"70",
          3017 => x"52",
          3018 => x"92",
          3019 => x"97",
          3020 => x"9f",
          3021 => x"a0",
          3022 => x"96",
          3023 => x"85",
          3024 => x"06",
          3025 => x"80",
          3026 => x"81",
          3027 => x"3f",
          3028 => x"51",
          3029 => x"80",
          3030 => x"3f",
          3031 => x"70",
          3032 => x"52",
          3033 => x"92",
          3034 => x"96",
          3035 => x"9f",
          3036 => x"e4",
          3037 => x"96",
          3038 => x"87",
          3039 => x"06",
          3040 => x"80",
          3041 => x"81",
          3042 => x"3f",
          3043 => x"51",
          3044 => x"80",
          3045 => x"3f",
          3046 => x"70",
          3047 => x"52",
          3048 => x"92",
          3049 => x"96",
          3050 => x"a0",
          3051 => x"a8",
          3052 => x"96",
          3053 => x"bb",
          3054 => x"0d",
          3055 => x"0d",
          3056 => x"05",
          3057 => x"70",
          3058 => x"80",
          3059 => x"ee",
          3060 => x"0b",
          3061 => x"33",
          3062 => x"38",
          3063 => x"a0",
          3064 => x"cc",
          3065 => x"f7",
          3066 => x"b5",
          3067 => x"70",
          3068 => x"08",
          3069 => x"82",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"34",
          3073 => x"b0",
          3074 => x"73",
          3075 => x"81",
          3076 => x"82",
          3077 => x"74",
          3078 => x"81",
          3079 => x"82",
          3080 => x"80",
          3081 => x"82",
          3082 => x"51",
          3083 => x"91",
          3084 => x"a8",
          3085 => x"cb",
          3086 => x"0b",
          3087 => x"a4",
          3088 => x"82",
          3089 => x"54",
          3090 => x"09",
          3091 => x"38",
          3092 => x"53",
          3093 => x"51",
          3094 => x"80",
          3095 => x"a8",
          3096 => x"0d",
          3097 => x"0d",
          3098 => x"82",
          3099 => x"40",
          3100 => x"7d",
          3101 => x"f5",
          3102 => x"a8",
          3103 => x"06",
          3104 => x"2e",
          3105 => x"a3",
          3106 => x"5a",
          3107 => x"a0",
          3108 => x"51",
          3109 => x"7d",
          3110 => x"82",
          3111 => x"80",
          3112 => x"82",
          3113 => x"7e",
          3114 => x"82",
          3115 => x"8d",
          3116 => x"70",
          3117 => x"a1",
          3118 => x"c8",
          3119 => x"70",
          3120 => x"f8",
          3121 => x"fd",
          3122 => x"3d",
          3123 => x"51",
          3124 => x"82",
          3125 => x"90",
          3126 => x"2c",
          3127 => x"80",
          3128 => x"99",
          3129 => x"c2",
          3130 => x"79",
          3131 => x"d1",
          3132 => x"24",
          3133 => x"80",
          3134 => x"38",
          3135 => x"80",
          3136 => x"c0",
          3137 => x"c0",
          3138 => x"38",
          3139 => x"24",
          3140 => x"79",
          3141 => x"8a",
          3142 => x"39",
          3143 => x"2e",
          3144 => x"79",
          3145 => x"92",
          3146 => x"c3",
          3147 => x"38",
          3148 => x"2e",
          3149 => x"8a",
          3150 => x"81",
          3151 => x"f2",
          3152 => x"83",
          3153 => x"79",
          3154 => x"89",
          3155 => x"f4",
          3156 => x"85",
          3157 => x"38",
          3158 => x"b5",
          3159 => x"11",
          3160 => x"05",
          3161 => x"3f",
          3162 => x"08",
          3163 => x"c6",
          3164 => x"fe",
          3165 => x"ff",
          3166 => x"d2",
          3167 => x"b5",
          3168 => x"2e",
          3169 => x"b5",
          3170 => x"11",
          3171 => x"05",
          3172 => x"3f",
          3173 => x"08",
          3174 => x"b5",
          3175 => x"82",
          3176 => x"d7",
          3177 => x"64",
          3178 => x"7c",
          3179 => x"38",
          3180 => x"7b",
          3181 => x"5d",
          3182 => x"26",
          3183 => x"d9",
          3184 => x"ff",
          3185 => x"ff",
          3186 => x"d1",
          3187 => x"b5",
          3188 => x"2e",
          3189 => x"b5",
          3190 => x"11",
          3191 => x"05",
          3192 => x"3f",
          3193 => x"08",
          3194 => x"ca",
          3195 => x"fe",
          3196 => x"ff",
          3197 => x"d1",
          3198 => x"b5",
          3199 => x"2e",
          3200 => x"82",
          3201 => x"d6",
          3202 => x"5b",
          3203 => x"81",
          3204 => x"5a",
          3205 => x"05",
          3206 => x"34",
          3207 => x"43",
          3208 => x"3d",
          3209 => x"53",
          3210 => x"51",
          3211 => x"82",
          3212 => x"80",
          3213 => x"38",
          3214 => x"fc",
          3215 => x"84",
          3216 => x"ef",
          3217 => x"a8",
          3218 => x"fc",
          3219 => x"3d",
          3220 => x"53",
          3221 => x"51",
          3222 => x"82",
          3223 => x"80",
          3224 => x"38",
          3225 => x"51",
          3226 => x"64",
          3227 => x"27",
          3228 => x"70",
          3229 => x"5f",
          3230 => x"7d",
          3231 => x"79",
          3232 => x"7a",
          3233 => x"52",
          3234 => x"51",
          3235 => x"3f",
          3236 => x"81",
          3237 => x"d5",
          3238 => x"f0",
          3239 => x"39",
          3240 => x"80",
          3241 => x"84",
          3242 => x"87",
          3243 => x"a8",
          3244 => x"38",
          3245 => x"33",
          3246 => x"2e",
          3247 => x"b3",
          3248 => x"80",
          3249 => x"b4",
          3250 => x"79",
          3251 => x"38",
          3252 => x"08",
          3253 => x"82",
          3254 => x"5a",
          3255 => x"88",
          3256 => x"dc",
          3257 => x"39",
          3258 => x"33",
          3259 => x"2e",
          3260 => x"b3",
          3261 => x"9a",
          3262 => x"92",
          3263 => x"80",
          3264 => x"82",
          3265 => x"45",
          3266 => x"b3",
          3267 => x"80",
          3268 => x"3d",
          3269 => x"53",
          3270 => x"51",
          3271 => x"82",
          3272 => x"80",
          3273 => x"b4",
          3274 => x"79",
          3275 => x"38",
          3276 => x"08",
          3277 => x"39",
          3278 => x"33",
          3279 => x"2e",
          3280 => x"b3",
          3281 => x"bb",
          3282 => x"96",
          3283 => x"80",
          3284 => x"82",
          3285 => x"44",
          3286 => x"b4",
          3287 => x"79",
          3288 => x"38",
          3289 => x"08",
          3290 => x"82",
          3291 => x"5a",
          3292 => x"88",
          3293 => x"f0",
          3294 => x"39",
          3295 => x"08",
          3296 => x"b5",
          3297 => x"11",
          3298 => x"05",
          3299 => x"3f",
          3300 => x"08",
          3301 => x"38",
          3302 => x"5d",
          3303 => x"83",
          3304 => x"7b",
          3305 => x"30",
          3306 => x"9f",
          3307 => x"06",
          3308 => x"5b",
          3309 => x"88",
          3310 => x"2e",
          3311 => x"43",
          3312 => x"51",
          3313 => x"a0",
          3314 => x"62",
          3315 => x"64",
          3316 => x"3f",
          3317 => x"51",
          3318 => x"b5",
          3319 => x"11",
          3320 => x"05",
          3321 => x"3f",
          3322 => x"08",
          3323 => x"c6",
          3324 => x"fe",
          3325 => x"ff",
          3326 => x"cd",
          3327 => x"b5",
          3328 => x"2e",
          3329 => x"5a",
          3330 => x"05",
          3331 => x"64",
          3332 => x"b5",
          3333 => x"11",
          3334 => x"05",
          3335 => x"3f",
          3336 => x"08",
          3337 => x"8e",
          3338 => x"33",
          3339 => x"a2",
          3340 => x"ab",
          3341 => x"f8",
          3342 => x"cc",
          3343 => x"46",
          3344 => x"79",
          3345 => x"ee",
          3346 => x"27",
          3347 => x"3d",
          3348 => x"53",
          3349 => x"51",
          3350 => x"82",
          3351 => x"80",
          3352 => x"64",
          3353 => x"cf",
          3354 => x"34",
          3355 => x"45",
          3356 => x"82",
          3357 => x"d2",
          3358 => x"ad",
          3359 => x"fe",
          3360 => x"ff",
          3361 => x"c6",
          3362 => x"b5",
          3363 => x"2e",
          3364 => x"b5",
          3365 => x"11",
          3366 => x"05",
          3367 => x"3f",
          3368 => x"08",
          3369 => x"38",
          3370 => x"80",
          3371 => x"7a",
          3372 => x"5c",
          3373 => x"b5",
          3374 => x"11",
          3375 => x"05",
          3376 => x"3f",
          3377 => x"08",
          3378 => x"ea",
          3379 => x"22",
          3380 => x"a2",
          3381 => x"a9",
          3382 => x"f8",
          3383 => x"cb",
          3384 => x"46",
          3385 => x"79",
          3386 => x"ca",
          3387 => x"26",
          3388 => x"82",
          3389 => x"39",
          3390 => x"f0",
          3391 => x"84",
          3392 => x"a8",
          3393 => x"a8",
          3394 => x"93",
          3395 => x"02",
          3396 => x"22",
          3397 => x"05",
          3398 => x"42",
          3399 => x"82",
          3400 => x"d0",
          3401 => x"a5",
          3402 => x"fe",
          3403 => x"ff",
          3404 => x"c4",
          3405 => x"b5",
          3406 => x"2e",
          3407 => x"b5",
          3408 => x"11",
          3409 => x"05",
          3410 => x"3f",
          3411 => x"08",
          3412 => x"38",
          3413 => x"0c",
          3414 => x"05",
          3415 => x"fe",
          3416 => x"ff",
          3417 => x"c4",
          3418 => x"b5",
          3419 => x"38",
          3420 => x"61",
          3421 => x"52",
          3422 => x"51",
          3423 => x"3f",
          3424 => x"7a",
          3425 => x"3f",
          3426 => x"33",
          3427 => x"2e",
          3428 => x"9f",
          3429 => x"38",
          3430 => x"f0",
          3431 => x"84",
          3432 => x"88",
          3433 => x"a8",
          3434 => x"8d",
          3435 => x"71",
          3436 => x"84",
          3437 => x"bb",
          3438 => x"9c",
          3439 => x"3f",
          3440 => x"b5",
          3441 => x"11",
          3442 => x"05",
          3443 => x"3f",
          3444 => x"08",
          3445 => x"de",
          3446 => x"82",
          3447 => x"ff",
          3448 => x"64",
          3449 => x"b5",
          3450 => x"11",
          3451 => x"05",
          3452 => x"3f",
          3453 => x"08",
          3454 => x"ba",
          3455 => x"82",
          3456 => x"ff",
          3457 => x"64",
          3458 => x"82",
          3459 => x"80",
          3460 => x"38",
          3461 => x"08",
          3462 => x"f4",
          3463 => x"b7",
          3464 => x"39",
          3465 => x"51",
          3466 => x"ff",
          3467 => x"f5",
          3468 => x"a3",
          3469 => x"cc",
          3470 => x"ff",
          3471 => x"b1",
          3472 => x"39",
          3473 => x"33",
          3474 => x"2e",
          3475 => x"7e",
          3476 => x"79",
          3477 => x"d6",
          3478 => x"ff",
          3479 => x"83",
          3480 => x"b5",
          3481 => x"81",
          3482 => x"2e",
          3483 => x"82",
          3484 => x"7b",
          3485 => x"38",
          3486 => x"7b",
          3487 => x"38",
          3488 => x"82",
          3489 => x"7c",
          3490 => x"c4",
          3491 => x"82",
          3492 => x"b5",
          3493 => x"05",
          3494 => x"a3",
          3495 => x"82",
          3496 => x"b5",
          3497 => x"05",
          3498 => x"93",
          3499 => x"7c",
          3500 => x"c4",
          3501 => x"82",
          3502 => x"b5",
          3503 => x"05",
          3504 => x"fb",
          3505 => x"7c",
          3506 => x"82",
          3507 => x"b5",
          3508 => x"05",
          3509 => x"e7",
          3510 => x"f8",
          3511 => x"cc",
          3512 => x"d8",
          3513 => x"65",
          3514 => x"82",
          3515 => x"82",
          3516 => x"b5",
          3517 => x"05",
          3518 => x"3f",
          3519 => x"08",
          3520 => x"08",
          3521 => x"70",
          3522 => x"25",
          3523 => x"40",
          3524 => x"83",
          3525 => x"81",
          3526 => x"06",
          3527 => x"2e",
          3528 => x"1c",
          3529 => x"06",
          3530 => x"fe",
          3531 => x"81",
          3532 => x"32",
          3533 => x"8a",
          3534 => x"2e",
          3535 => x"f2",
          3536 => x"a3",
          3537 => x"bc",
          3538 => x"39",
          3539 => x"80",
          3540 => x"d8",
          3541 => x"94",
          3542 => x"54",
          3543 => x"80",
          3544 => x"e3",
          3545 => x"b5",
          3546 => x"2b",
          3547 => x"53",
          3548 => x"52",
          3549 => x"ac",
          3550 => x"b5",
          3551 => x"75",
          3552 => x"94",
          3553 => x"54",
          3554 => x"80",
          3555 => x"e3",
          3556 => x"b5",
          3557 => x"2b",
          3558 => x"53",
          3559 => x"52",
          3560 => x"80",
          3561 => x"b5",
          3562 => x"75",
          3563 => x"83",
          3564 => x"94",
          3565 => x"80",
          3566 => x"c0",
          3567 => x"82",
          3568 => x"cb",
          3569 => x"f5",
          3570 => x"f8",
          3571 => x"02",
          3572 => x"05",
          3573 => x"8d",
          3574 => x"82",
          3575 => x"89",
          3576 => x"87",
          3577 => x"90",
          3578 => x"3f",
          3579 => x"51",
          3580 => x"82",
          3581 => x"cb",
          3582 => x"dd",
          3583 => x"e6",
          3584 => x"ec",
          3585 => x"dd",
          3586 => x"fe",
          3587 => x"52",
          3588 => x"88",
          3589 => x"d9",
          3590 => x"a8",
          3591 => x"06",
          3592 => x"14",
          3593 => x"80",
          3594 => x"71",
          3595 => x"0c",
          3596 => x"04",
          3597 => x"76",
          3598 => x"55",
          3599 => x"54",
          3600 => x"81",
          3601 => x"33",
          3602 => x"2e",
          3603 => x"86",
          3604 => x"53",
          3605 => x"33",
          3606 => x"2e",
          3607 => x"86",
          3608 => x"53",
          3609 => x"52",
          3610 => x"09",
          3611 => x"38",
          3612 => x"12",
          3613 => x"33",
          3614 => x"a2",
          3615 => x"81",
          3616 => x"2e",
          3617 => x"ea",
          3618 => x"81",
          3619 => x"72",
          3620 => x"70",
          3621 => x"38",
          3622 => x"80",
          3623 => x"73",
          3624 => x"72",
          3625 => x"70",
          3626 => x"81",
          3627 => x"81",
          3628 => x"32",
          3629 => x"80",
          3630 => x"51",
          3631 => x"80",
          3632 => x"80",
          3633 => x"05",
          3634 => x"75",
          3635 => x"70",
          3636 => x"0c",
          3637 => x"04",
          3638 => x"76",
          3639 => x"80",
          3640 => x"86",
          3641 => x"52",
          3642 => x"bd",
          3643 => x"b5",
          3644 => x"38",
          3645 => x"39",
          3646 => x"82",
          3647 => x"86",
          3648 => x"fc",
          3649 => x"82",
          3650 => x"05",
          3651 => x"52",
          3652 => x"81",
          3653 => x"13",
          3654 => x"51",
          3655 => x"9e",
          3656 => x"38",
          3657 => x"51",
          3658 => x"97",
          3659 => x"38",
          3660 => x"51",
          3661 => x"bb",
          3662 => x"38",
          3663 => x"51",
          3664 => x"bb",
          3665 => x"38",
          3666 => x"55",
          3667 => x"87",
          3668 => x"d9",
          3669 => x"22",
          3670 => x"73",
          3671 => x"80",
          3672 => x"0b",
          3673 => x"9c",
          3674 => x"87",
          3675 => x"0c",
          3676 => x"87",
          3677 => x"0c",
          3678 => x"87",
          3679 => x"0c",
          3680 => x"87",
          3681 => x"0c",
          3682 => x"87",
          3683 => x"0c",
          3684 => x"87",
          3685 => x"0c",
          3686 => x"98",
          3687 => x"87",
          3688 => x"0c",
          3689 => x"c0",
          3690 => x"80",
          3691 => x"b5",
          3692 => x"3d",
          3693 => x"3d",
          3694 => x"87",
          3695 => x"5d",
          3696 => x"87",
          3697 => x"08",
          3698 => x"23",
          3699 => x"b8",
          3700 => x"82",
          3701 => x"c0",
          3702 => x"5a",
          3703 => x"34",
          3704 => x"b0",
          3705 => x"84",
          3706 => x"c0",
          3707 => x"5a",
          3708 => x"34",
          3709 => x"a8",
          3710 => x"86",
          3711 => x"c0",
          3712 => x"5c",
          3713 => x"23",
          3714 => x"a0",
          3715 => x"8a",
          3716 => x"7d",
          3717 => x"ff",
          3718 => x"7b",
          3719 => x"06",
          3720 => x"33",
          3721 => x"33",
          3722 => x"33",
          3723 => x"33",
          3724 => x"33",
          3725 => x"ff",
          3726 => x"82",
          3727 => x"ff",
          3728 => x"8f",
          3729 => x"fb",
          3730 => x"9f",
          3731 => x"b3",
          3732 => x"81",
          3733 => x"55",
          3734 => x"94",
          3735 => x"80",
          3736 => x"87",
          3737 => x"51",
          3738 => x"96",
          3739 => x"06",
          3740 => x"70",
          3741 => x"38",
          3742 => x"70",
          3743 => x"51",
          3744 => x"72",
          3745 => x"81",
          3746 => x"70",
          3747 => x"38",
          3748 => x"70",
          3749 => x"51",
          3750 => x"38",
          3751 => x"06",
          3752 => x"94",
          3753 => x"80",
          3754 => x"87",
          3755 => x"52",
          3756 => x"74",
          3757 => x"0c",
          3758 => x"04",
          3759 => x"02",
          3760 => x"70",
          3761 => x"2a",
          3762 => x"70",
          3763 => x"34",
          3764 => x"04",
          3765 => x"02",
          3766 => x"58",
          3767 => x"09",
          3768 => x"38",
          3769 => x"51",
          3770 => x"b3",
          3771 => x"81",
          3772 => x"56",
          3773 => x"84",
          3774 => x"2e",
          3775 => x"c0",
          3776 => x"72",
          3777 => x"2a",
          3778 => x"55",
          3779 => x"80",
          3780 => x"73",
          3781 => x"81",
          3782 => x"72",
          3783 => x"81",
          3784 => x"06",
          3785 => x"80",
          3786 => x"73",
          3787 => x"81",
          3788 => x"72",
          3789 => x"75",
          3790 => x"53",
          3791 => x"80",
          3792 => x"2e",
          3793 => x"c0",
          3794 => x"77",
          3795 => x"0b",
          3796 => x"0c",
          3797 => x"04",
          3798 => x"79",
          3799 => x"33",
          3800 => x"06",
          3801 => x"70",
          3802 => x"fc",
          3803 => x"ff",
          3804 => x"82",
          3805 => x"70",
          3806 => x"59",
          3807 => x"87",
          3808 => x"51",
          3809 => x"86",
          3810 => x"94",
          3811 => x"08",
          3812 => x"70",
          3813 => x"54",
          3814 => x"2e",
          3815 => x"91",
          3816 => x"06",
          3817 => x"d7",
          3818 => x"32",
          3819 => x"51",
          3820 => x"2e",
          3821 => x"93",
          3822 => x"06",
          3823 => x"ff",
          3824 => x"81",
          3825 => x"87",
          3826 => x"52",
          3827 => x"86",
          3828 => x"94",
          3829 => x"72",
          3830 => x"74",
          3831 => x"ff",
          3832 => x"57",
          3833 => x"38",
          3834 => x"a8",
          3835 => x"0d",
          3836 => x"0d",
          3837 => x"33",
          3838 => x"06",
          3839 => x"c0",
          3840 => x"72",
          3841 => x"38",
          3842 => x"94",
          3843 => x"70",
          3844 => x"81",
          3845 => x"51",
          3846 => x"e2",
          3847 => x"ff",
          3848 => x"c0",
          3849 => x"70",
          3850 => x"38",
          3851 => x"90",
          3852 => x"70",
          3853 => x"82",
          3854 => x"51",
          3855 => x"04",
          3856 => x"82",
          3857 => x"81",
          3858 => x"b5",
          3859 => x"fe",
          3860 => x"b3",
          3861 => x"81",
          3862 => x"53",
          3863 => x"84",
          3864 => x"2e",
          3865 => x"c0",
          3866 => x"71",
          3867 => x"2a",
          3868 => x"51",
          3869 => x"52",
          3870 => x"a0",
          3871 => x"ff",
          3872 => x"c0",
          3873 => x"70",
          3874 => x"38",
          3875 => x"90",
          3876 => x"70",
          3877 => x"98",
          3878 => x"51",
          3879 => x"a8",
          3880 => x"0d",
          3881 => x"0d",
          3882 => x"80",
          3883 => x"2a",
          3884 => x"51",
          3885 => x"84",
          3886 => x"c0",
          3887 => x"82",
          3888 => x"87",
          3889 => x"08",
          3890 => x"0c",
          3891 => x"94",
          3892 => x"d4",
          3893 => x"9e",
          3894 => x"b3",
          3895 => x"c0",
          3896 => x"82",
          3897 => x"87",
          3898 => x"08",
          3899 => x"0c",
          3900 => x"ac",
          3901 => x"e4",
          3902 => x"9e",
          3903 => x"b3",
          3904 => x"c0",
          3905 => x"82",
          3906 => x"87",
          3907 => x"08",
          3908 => x"0c",
          3909 => x"bc",
          3910 => x"f4",
          3911 => x"9e",
          3912 => x"b3",
          3913 => x"c0",
          3914 => x"82",
          3915 => x"87",
          3916 => x"08",
          3917 => x"b4",
          3918 => x"c0",
          3919 => x"82",
          3920 => x"87",
          3921 => x"08",
          3922 => x"0c",
          3923 => x"8c",
          3924 => x"8c",
          3925 => x"82",
          3926 => x"80",
          3927 => x"9e",
          3928 => x"84",
          3929 => x"51",
          3930 => x"80",
          3931 => x"81",
          3932 => x"b4",
          3933 => x"0b",
          3934 => x"90",
          3935 => x"80",
          3936 => x"52",
          3937 => x"2e",
          3938 => x"52",
          3939 => x"92",
          3940 => x"87",
          3941 => x"08",
          3942 => x"0a",
          3943 => x"52",
          3944 => x"83",
          3945 => x"71",
          3946 => x"34",
          3947 => x"c0",
          3948 => x"70",
          3949 => x"06",
          3950 => x"70",
          3951 => x"38",
          3952 => x"82",
          3953 => x"80",
          3954 => x"9e",
          3955 => x"a0",
          3956 => x"51",
          3957 => x"80",
          3958 => x"81",
          3959 => x"b4",
          3960 => x"0b",
          3961 => x"90",
          3962 => x"80",
          3963 => x"52",
          3964 => x"2e",
          3965 => x"52",
          3966 => x"96",
          3967 => x"87",
          3968 => x"08",
          3969 => x"80",
          3970 => x"52",
          3971 => x"83",
          3972 => x"71",
          3973 => x"34",
          3974 => x"c0",
          3975 => x"70",
          3976 => x"06",
          3977 => x"70",
          3978 => x"38",
          3979 => x"82",
          3980 => x"80",
          3981 => x"9e",
          3982 => x"81",
          3983 => x"51",
          3984 => x"80",
          3985 => x"81",
          3986 => x"b4",
          3987 => x"0b",
          3988 => x"90",
          3989 => x"c0",
          3990 => x"52",
          3991 => x"2e",
          3992 => x"52",
          3993 => x"9a",
          3994 => x"87",
          3995 => x"08",
          3996 => x"06",
          3997 => x"70",
          3998 => x"38",
          3999 => x"82",
          4000 => x"87",
          4001 => x"08",
          4002 => x"06",
          4003 => x"51",
          4004 => x"82",
          4005 => x"80",
          4006 => x"9e",
          4007 => x"84",
          4008 => x"52",
          4009 => x"2e",
          4010 => x"52",
          4011 => x"9d",
          4012 => x"9e",
          4013 => x"83",
          4014 => x"84",
          4015 => x"51",
          4016 => x"9e",
          4017 => x"87",
          4018 => x"08",
          4019 => x"51",
          4020 => x"80",
          4021 => x"81",
          4022 => x"b4",
          4023 => x"c0",
          4024 => x"70",
          4025 => x"51",
          4026 => x"a0",
          4027 => x"0d",
          4028 => x"0d",
          4029 => x"51",
          4030 => x"3f",
          4031 => x"33",
          4032 => x"2e",
          4033 => x"a4",
          4034 => x"bc",
          4035 => x"a5",
          4036 => x"bc",
          4037 => x"b4",
          4038 => x"73",
          4039 => x"38",
          4040 => x"08",
          4041 => x"08",
          4042 => x"82",
          4043 => x"ff",
          4044 => x"82",
          4045 => x"54",
          4046 => x"94",
          4047 => x"e4",
          4048 => x"e8",
          4049 => x"52",
          4050 => x"51",
          4051 => x"3f",
          4052 => x"33",
          4053 => x"2e",
          4054 => x"b3",
          4055 => x"b3",
          4056 => x"54",
          4057 => x"d8",
          4058 => x"eb",
          4059 => x"95",
          4060 => x"80",
          4061 => x"82",
          4062 => x"82",
          4063 => x"11",
          4064 => x"a5",
          4065 => x"94",
          4066 => x"b4",
          4067 => x"73",
          4068 => x"38",
          4069 => x"08",
          4070 => x"08",
          4071 => x"82",
          4072 => x"ff",
          4073 => x"82",
          4074 => x"54",
          4075 => x"8e",
          4076 => x"9c",
          4077 => x"a6",
          4078 => x"94",
          4079 => x"b4",
          4080 => x"73",
          4081 => x"38",
          4082 => x"33",
          4083 => x"cc",
          4084 => x"83",
          4085 => x"9d",
          4086 => x"80",
          4087 => x"82",
          4088 => x"52",
          4089 => x"51",
          4090 => x"3f",
          4091 => x"33",
          4092 => x"2e",
          4093 => x"a7",
          4094 => x"bb",
          4095 => x"b4",
          4096 => x"73",
          4097 => x"38",
          4098 => x"51",
          4099 => x"3f",
          4100 => x"33",
          4101 => x"2e",
          4102 => x"a7",
          4103 => x"ba",
          4104 => x"b4",
          4105 => x"73",
          4106 => x"38",
          4107 => x"51",
          4108 => x"3f",
          4109 => x"33",
          4110 => x"2e",
          4111 => x"a7",
          4112 => x"ba",
          4113 => x"a7",
          4114 => x"ba",
          4115 => x"b3",
          4116 => x"82",
          4117 => x"ff",
          4118 => x"82",
          4119 => x"52",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"08",
          4123 => x"ac",
          4124 => x"e3",
          4125 => x"d4",
          4126 => x"88",
          4127 => x"80",
          4128 => x"a8",
          4129 => x"92",
          4130 => x"b4",
          4131 => x"bd",
          4132 => x"75",
          4133 => x"3f",
          4134 => x"08",
          4135 => x"29",
          4136 => x"54",
          4137 => x"a8",
          4138 => x"a9",
          4139 => x"92",
          4140 => x"b4",
          4141 => x"73",
          4142 => x"38",
          4143 => x"08",
          4144 => x"c0",
          4145 => x"d0",
          4146 => x"b5",
          4147 => x"84",
          4148 => x"71",
          4149 => x"82",
          4150 => x"52",
          4151 => x"51",
          4152 => x"3f",
          4153 => x"33",
          4154 => x"2e",
          4155 => x"b4",
          4156 => x"bd",
          4157 => x"75",
          4158 => x"3f",
          4159 => x"08",
          4160 => x"29",
          4161 => x"54",
          4162 => x"a8",
          4163 => x"a9",
          4164 => x"91",
          4165 => x"a1",
          4166 => x"b8",
          4167 => x"3d",
          4168 => x"3d",
          4169 => x"05",
          4170 => x"52",
          4171 => x"aa",
          4172 => x"29",
          4173 => x"05",
          4174 => x"04",
          4175 => x"51",
          4176 => x"aa",
          4177 => x"39",
          4178 => x"51",
          4179 => x"aa",
          4180 => x"39",
          4181 => x"51",
          4182 => x"aa",
          4183 => x"b8",
          4184 => x"3d",
          4185 => x"88",
          4186 => x"80",
          4187 => x"96",
          4188 => x"82",
          4189 => x"87",
          4190 => x"0c",
          4191 => x"0d",
          4192 => x"70",
          4193 => x"98",
          4194 => x"2c",
          4195 => x"70",
          4196 => x"53",
          4197 => x"51",
          4198 => x"aa",
          4199 => x"55",
          4200 => x"25",
          4201 => x"aa",
          4202 => x"12",
          4203 => x"97",
          4204 => x"33",
          4205 => x"70",
          4206 => x"81",
          4207 => x"81",
          4208 => x"b5",
          4209 => x"3d",
          4210 => x"3d",
          4211 => x"84",
          4212 => x"33",
          4213 => x"55",
          4214 => x"2e",
          4215 => x"51",
          4216 => x"3f",
          4217 => x"ba",
          4218 => x"51",
          4219 => x"3f",
          4220 => x"05",
          4221 => x"34",
          4222 => x"06",
          4223 => x"76",
          4224 => x"80",
          4225 => x"34",
          4226 => x"04",
          4227 => x"7c",
          4228 => x"b7",
          4229 => x"88",
          4230 => x"33",
          4231 => x"33",
          4232 => x"82",
          4233 => x"70",
          4234 => x"59",
          4235 => x"74",
          4236 => x"38",
          4237 => x"b2",
          4238 => x"80",
          4239 => x"29",
          4240 => x"05",
          4241 => x"54",
          4242 => x"9d",
          4243 => x"b5",
          4244 => x"0c",
          4245 => x"33",
          4246 => x"82",
          4247 => x"70",
          4248 => x"5a",
          4249 => x"a6",
          4250 => x"78",
          4251 => x"c4",
          4252 => x"b5",
          4253 => x"05",
          4254 => x"b5",
          4255 => x"81",
          4256 => x"93",
          4257 => x"38",
          4258 => x"b5",
          4259 => x"80",
          4260 => x"82",
          4261 => x"56",
          4262 => x"ac",
          4263 => x"f8",
          4264 => x"a4",
          4265 => x"fc",
          4266 => x"53",
          4267 => x"51",
          4268 => x"3f",
          4269 => x"08",
          4270 => x"81",
          4271 => x"82",
          4272 => x"51",
          4273 => x"3f",
          4274 => x"04",
          4275 => x"82",
          4276 => x"93",
          4277 => x"52",
          4278 => x"89",
          4279 => x"99",
          4280 => x"73",
          4281 => x"84",
          4282 => x"73",
          4283 => x"38",
          4284 => x"b5",
          4285 => x"b4",
          4286 => x"71",
          4287 => x"38",
          4288 => x"dd",
          4289 => x"b4",
          4290 => x"98",
          4291 => x"0b",
          4292 => x"0c",
          4293 => x"04",
          4294 => x"81",
          4295 => x"82",
          4296 => x"51",
          4297 => x"3f",
          4298 => x"08",
          4299 => x"82",
          4300 => x"53",
          4301 => x"88",
          4302 => x"56",
          4303 => x"3f",
          4304 => x"08",
          4305 => x"38",
          4306 => x"da",
          4307 => x"a8",
          4308 => x"0b",
          4309 => x"08",
          4310 => x"82",
          4311 => x"ff",
          4312 => x"55",
          4313 => x"34",
          4314 => x"52",
          4315 => x"ad",
          4316 => x"ff",
          4317 => x"74",
          4318 => x"81",
          4319 => x"38",
          4320 => x"04",
          4321 => x"aa",
          4322 => x"3d",
          4323 => x"81",
          4324 => x"80",
          4325 => x"fc",
          4326 => x"e1",
          4327 => x"b5",
          4328 => x"95",
          4329 => x"82",
          4330 => x"54",
          4331 => x"52",
          4332 => x"52",
          4333 => x"c0",
          4334 => x"a8",
          4335 => x"a5",
          4336 => x"ff",
          4337 => x"82",
          4338 => x"81",
          4339 => x"80",
          4340 => x"a8",
          4341 => x"38",
          4342 => x"08",
          4343 => x"17",
          4344 => x"74",
          4345 => x"70",
          4346 => x"07",
          4347 => x"55",
          4348 => x"2e",
          4349 => x"ff",
          4350 => x"b4",
          4351 => x"11",
          4352 => x"80",
          4353 => x"82",
          4354 => x"80",
          4355 => x"82",
          4356 => x"ff",
          4357 => x"78",
          4358 => x"81",
          4359 => x"75",
          4360 => x"ff",
          4361 => x"79",
          4362 => x"fa",
          4363 => x"08",
          4364 => x"a8",
          4365 => x"80",
          4366 => x"b5",
          4367 => x"3d",
          4368 => x"3d",
          4369 => x"71",
          4370 => x"33",
          4371 => x"58",
          4372 => x"09",
          4373 => x"38",
          4374 => x"05",
          4375 => x"27",
          4376 => x"17",
          4377 => x"71",
          4378 => x"55",
          4379 => x"09",
          4380 => x"38",
          4381 => x"ea",
          4382 => x"73",
          4383 => x"b5",
          4384 => x"08",
          4385 => x"be",
          4386 => x"b5",
          4387 => x"79",
          4388 => x"51",
          4389 => x"82",
          4390 => x"80",
          4391 => x"15",
          4392 => x"81",
          4393 => x"74",
          4394 => x"38",
          4395 => x"e8",
          4396 => x"81",
          4397 => x"3d",
          4398 => x"f8",
          4399 => x"ab",
          4400 => x"b5",
          4401 => x"2e",
          4402 => x"1b",
          4403 => x"77",
          4404 => x"3f",
          4405 => x"08",
          4406 => x"55",
          4407 => x"74",
          4408 => x"81",
          4409 => x"ff",
          4410 => x"82",
          4411 => x"8b",
          4412 => x"73",
          4413 => x"0c",
          4414 => x"04",
          4415 => x"b0",
          4416 => x"3d",
          4417 => x"08",
          4418 => x"80",
          4419 => x"34",
          4420 => x"33",
          4421 => x"08",
          4422 => x"81",
          4423 => x"82",
          4424 => x"55",
          4425 => x"38",
          4426 => x"80",
          4427 => x"38",
          4428 => x"06",
          4429 => x"80",
          4430 => x"38",
          4431 => x"c0",
          4432 => x"a8",
          4433 => x"fc",
          4434 => x"a8",
          4435 => x"81",
          4436 => x"53",
          4437 => x"b5",
          4438 => x"80",
          4439 => x"82",
          4440 => x"80",
          4441 => x"82",
          4442 => x"ff",
          4443 => x"80",
          4444 => x"b5",
          4445 => x"82",
          4446 => x"53",
          4447 => x"90",
          4448 => x"54",
          4449 => x"3f",
          4450 => x"08",
          4451 => x"a8",
          4452 => x"09",
          4453 => x"d0",
          4454 => x"a8",
          4455 => x"bc",
          4456 => x"b5",
          4457 => x"80",
          4458 => x"a8",
          4459 => x"38",
          4460 => x"08",
          4461 => x"17",
          4462 => x"74",
          4463 => x"74",
          4464 => x"52",
          4465 => x"c4",
          4466 => x"70",
          4467 => x"5c",
          4468 => x"27",
          4469 => x"5b",
          4470 => x"09",
          4471 => x"97",
          4472 => x"75",
          4473 => x"34",
          4474 => x"82",
          4475 => x"80",
          4476 => x"f9",
          4477 => x"3d",
          4478 => x"3f",
          4479 => x"08",
          4480 => x"98",
          4481 => x"78",
          4482 => x"38",
          4483 => x"06",
          4484 => x"33",
          4485 => x"70",
          4486 => x"cc",
          4487 => x"98",
          4488 => x"2c",
          4489 => x"05",
          4490 => x"82",
          4491 => x"70",
          4492 => x"33",
          4493 => x"51",
          4494 => x"59",
          4495 => x"56",
          4496 => x"80",
          4497 => x"74",
          4498 => x"74",
          4499 => x"29",
          4500 => x"05",
          4501 => x"51",
          4502 => x"24",
          4503 => x"76",
          4504 => x"77",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"54",
          4508 => x"d7",
          4509 => x"cc",
          4510 => x"56",
          4511 => x"81",
          4512 => x"81",
          4513 => x"70",
          4514 => x"81",
          4515 => x"51",
          4516 => x"26",
          4517 => x"53",
          4518 => x"51",
          4519 => x"82",
          4520 => x"81",
          4521 => x"73",
          4522 => x"39",
          4523 => x"80",
          4524 => x"38",
          4525 => x"74",
          4526 => x"34",
          4527 => x"70",
          4528 => x"cc",
          4529 => x"98",
          4530 => x"2c",
          4531 => x"70",
          4532 => x"aa",
          4533 => x"5e",
          4534 => x"57",
          4535 => x"74",
          4536 => x"81",
          4537 => x"38",
          4538 => x"14",
          4539 => x"80",
          4540 => x"d4",
          4541 => x"82",
          4542 => x"92",
          4543 => x"cc",
          4544 => x"82",
          4545 => x"78",
          4546 => x"75",
          4547 => x"54",
          4548 => x"fd",
          4549 => x"84",
          4550 => x"a4",
          4551 => x"08",
          4552 => x"dc",
          4553 => x"7e",
          4554 => x"38",
          4555 => x"33",
          4556 => x"27",
          4557 => x"98",
          4558 => x"2c",
          4559 => x"75",
          4560 => x"74",
          4561 => x"33",
          4562 => x"74",
          4563 => x"29",
          4564 => x"05",
          4565 => x"82",
          4566 => x"56",
          4567 => x"39",
          4568 => x"33",
          4569 => x"54",
          4570 => x"dc",
          4571 => x"54",
          4572 => x"74",
          4573 => x"d8",
          4574 => x"7e",
          4575 => x"81",
          4576 => x"82",
          4577 => x"82",
          4578 => x"70",
          4579 => x"29",
          4580 => x"05",
          4581 => x"82",
          4582 => x"5a",
          4583 => x"74",
          4584 => x"38",
          4585 => x"33",
          4586 => x"ae",
          4587 => x"81",
          4588 => x"81",
          4589 => x"70",
          4590 => x"cc",
          4591 => x"51",
          4592 => x"24",
          4593 => x"cc",
          4594 => x"98",
          4595 => x"2c",
          4596 => x"33",
          4597 => x"56",
          4598 => x"fc",
          4599 => x"51",
          4600 => x"3f",
          4601 => x"0a",
          4602 => x"0a",
          4603 => x"2c",
          4604 => x"33",
          4605 => x"73",
          4606 => x"38",
          4607 => x"83",
          4608 => x"0b",
          4609 => x"82",
          4610 => x"80",
          4611 => x"f0",
          4612 => x"3f",
          4613 => x"82",
          4614 => x"70",
          4615 => x"55",
          4616 => x"2e",
          4617 => x"82",
          4618 => x"ff",
          4619 => x"82",
          4620 => x"ff",
          4621 => x"82",
          4622 => x"88",
          4623 => x"e6",
          4624 => x"dc",
          4625 => x"2b",
          4626 => x"82",
          4627 => x"57",
          4628 => x"74",
          4629 => x"38",
          4630 => x"81",
          4631 => x"34",
          4632 => x"ff",
          4633 => x"74",
          4634 => x"29",
          4635 => x"05",
          4636 => x"82",
          4637 => x"58",
          4638 => x"75",
          4639 => x"a0",
          4640 => x"a2",
          4641 => x"dc",
          4642 => x"2b",
          4643 => x"82",
          4644 => x"57",
          4645 => x"74",
          4646 => x"da",
          4647 => x"ff",
          4648 => x"74",
          4649 => x"29",
          4650 => x"05",
          4651 => x"82",
          4652 => x"58",
          4653 => x"75",
          4654 => x"fa",
          4655 => x"cc",
          4656 => x"05",
          4657 => x"34",
          4658 => x"ac",
          4659 => x"cc",
          4660 => x"51",
          4661 => x"82",
          4662 => x"81",
          4663 => x"73",
          4664 => x"cc",
          4665 => x"73",
          4666 => x"38",
          4667 => x"52",
          4668 => x"98",
          4669 => x"80",
          4670 => x"0b",
          4671 => x"34",
          4672 => x"cc",
          4673 => x"82",
          4674 => x"af",
          4675 => x"82",
          4676 => x"54",
          4677 => x"f9",
          4678 => x"51",
          4679 => x"3f",
          4680 => x"33",
          4681 => x"73",
          4682 => x"34",
          4683 => x"06",
          4684 => x"82",
          4685 => x"82",
          4686 => x"55",
          4687 => x"2e",
          4688 => x"ff",
          4689 => x"82",
          4690 => x"74",
          4691 => x"98",
          4692 => x"ff",
          4693 => x"55",
          4694 => x"a8",
          4695 => x"54",
          4696 => x"74",
          4697 => x"51",
          4698 => x"3f",
          4699 => x"0a",
          4700 => x"0a",
          4701 => x"2c",
          4702 => x"33",
          4703 => x"75",
          4704 => x"38",
          4705 => x"ab",
          4706 => x"cc",
          4707 => x"98",
          4708 => x"2c",
          4709 => x"33",
          4710 => x"57",
          4711 => x"f8",
          4712 => x"51",
          4713 => x"3f",
          4714 => x"0a",
          4715 => x"0a",
          4716 => x"2c",
          4717 => x"33",
          4718 => x"75",
          4719 => x"38",
          4720 => x"82",
          4721 => x"70",
          4722 => x"82",
          4723 => x"59",
          4724 => x"77",
          4725 => x"38",
          4726 => x"73",
          4727 => x"34",
          4728 => x"33",
          4729 => x"aa",
          4730 => x"cc",
          4731 => x"81",
          4732 => x"cc",
          4733 => x"56",
          4734 => x"26",
          4735 => x"f6",
          4736 => x"dc",
          4737 => x"82",
          4738 => x"ef",
          4739 => x"0b",
          4740 => x"34",
          4741 => x"cc",
          4742 => x"da",
          4743 => x"38",
          4744 => x"08",
          4745 => x"2e",
          4746 => x"51",
          4747 => x"3f",
          4748 => x"08",
          4749 => x"34",
          4750 => x"08",
          4751 => x"81",
          4752 => x"52",
          4753 => x"b4",
          4754 => x"5b",
          4755 => x"7a",
          4756 => x"b4",
          4757 => x"11",
          4758 => x"74",
          4759 => x"38",
          4760 => x"b2",
          4761 => x"b5",
          4762 => x"cc",
          4763 => x"b5",
          4764 => x"ff",
          4765 => x"53",
          4766 => x"51",
          4767 => x"3f",
          4768 => x"80",
          4769 => x"08",
          4770 => x"2e",
          4771 => x"74",
          4772 => x"92",
          4773 => x"7a",
          4774 => x"81",
          4775 => x"82",
          4776 => x"55",
          4777 => x"a4",
          4778 => x"ff",
          4779 => x"82",
          4780 => x"82",
          4781 => x"82",
          4782 => x"81",
          4783 => x"05",
          4784 => x"79",
          4785 => x"be",
          4786 => x"39",
          4787 => x"82",
          4788 => x"70",
          4789 => x"74",
          4790 => x"38",
          4791 => x"b1",
          4792 => x"b5",
          4793 => x"cc",
          4794 => x"b5",
          4795 => x"ff",
          4796 => x"53",
          4797 => x"51",
          4798 => x"3f",
          4799 => x"73",
          4800 => x"5b",
          4801 => x"82",
          4802 => x"74",
          4803 => x"cc",
          4804 => x"cc",
          4805 => x"79",
          4806 => x"3f",
          4807 => x"82",
          4808 => x"70",
          4809 => x"82",
          4810 => x"59",
          4811 => x"77",
          4812 => x"38",
          4813 => x"73",
          4814 => x"34",
          4815 => x"33",
          4816 => x"a7",
          4817 => x"ae",
          4818 => x"dc",
          4819 => x"80",
          4820 => x"38",
          4821 => x"a7",
          4822 => x"cc",
          4823 => x"05",
          4824 => x"cc",
          4825 => x"8e",
          4826 => x"0d",
          4827 => x"0b",
          4828 => x"0c",
          4829 => x"82",
          4830 => x"90",
          4831 => x"52",
          4832 => x"51",
          4833 => x"3f",
          4834 => x"08",
          4835 => x"77",
          4836 => x"57",
          4837 => x"34",
          4838 => x"08",
          4839 => x"15",
          4840 => x"15",
          4841 => x"a0",
          4842 => x"86",
          4843 => x"87",
          4844 => x"b5",
          4845 => x"b5",
          4846 => x"05",
          4847 => x"07",
          4848 => x"ff",
          4849 => x"2a",
          4850 => x"56",
          4851 => x"34",
          4852 => x"34",
          4853 => x"22",
          4854 => x"82",
          4855 => x"05",
          4856 => x"55",
          4857 => x"15",
          4858 => x"15",
          4859 => x"0d",
          4860 => x"0d",
          4861 => x"51",
          4862 => x"8f",
          4863 => x"83",
          4864 => x"70",
          4865 => x"06",
          4866 => x"70",
          4867 => x"0c",
          4868 => x"04",
          4869 => x"02",
          4870 => x"02",
          4871 => x"05",
          4872 => x"82",
          4873 => x"71",
          4874 => x"11",
          4875 => x"73",
          4876 => x"81",
          4877 => x"88",
          4878 => x"a4",
          4879 => x"22",
          4880 => x"ff",
          4881 => x"88",
          4882 => x"52",
          4883 => x"5b",
          4884 => x"55",
          4885 => x"70",
          4886 => x"82",
          4887 => x"14",
          4888 => x"52",
          4889 => x"15",
          4890 => x"15",
          4891 => x"a0",
          4892 => x"70",
          4893 => x"33",
          4894 => x"07",
          4895 => x"8f",
          4896 => x"51",
          4897 => x"71",
          4898 => x"ff",
          4899 => x"88",
          4900 => x"51",
          4901 => x"34",
          4902 => x"06",
          4903 => x"12",
          4904 => x"a0",
          4905 => x"71",
          4906 => x"81",
          4907 => x"3d",
          4908 => x"3d",
          4909 => x"a0",
          4910 => x"05",
          4911 => x"70",
          4912 => x"11",
          4913 => x"87",
          4914 => x"8b",
          4915 => x"2b",
          4916 => x"59",
          4917 => x"72",
          4918 => x"33",
          4919 => x"71",
          4920 => x"70",
          4921 => x"56",
          4922 => x"84",
          4923 => x"85",
          4924 => x"b5",
          4925 => x"14",
          4926 => x"85",
          4927 => x"8b",
          4928 => x"2b",
          4929 => x"57",
          4930 => x"86",
          4931 => x"13",
          4932 => x"2b",
          4933 => x"2a",
          4934 => x"52",
          4935 => x"34",
          4936 => x"34",
          4937 => x"08",
          4938 => x"81",
          4939 => x"88",
          4940 => x"81",
          4941 => x"70",
          4942 => x"51",
          4943 => x"71",
          4944 => x"81",
          4945 => x"3d",
          4946 => x"3d",
          4947 => x"05",
          4948 => x"a0",
          4949 => x"2b",
          4950 => x"33",
          4951 => x"71",
          4952 => x"70",
          4953 => x"70",
          4954 => x"33",
          4955 => x"71",
          4956 => x"53",
          4957 => x"52",
          4958 => x"53",
          4959 => x"25",
          4960 => x"72",
          4961 => x"3f",
          4962 => x"08",
          4963 => x"33",
          4964 => x"71",
          4965 => x"83",
          4966 => x"11",
          4967 => x"12",
          4968 => x"2b",
          4969 => x"2b",
          4970 => x"06",
          4971 => x"51",
          4972 => x"53",
          4973 => x"88",
          4974 => x"72",
          4975 => x"73",
          4976 => x"82",
          4977 => x"70",
          4978 => x"81",
          4979 => x"8b",
          4980 => x"2b",
          4981 => x"57",
          4982 => x"70",
          4983 => x"33",
          4984 => x"07",
          4985 => x"ff",
          4986 => x"2a",
          4987 => x"58",
          4988 => x"34",
          4989 => x"34",
          4990 => x"04",
          4991 => x"82",
          4992 => x"02",
          4993 => x"05",
          4994 => x"2b",
          4995 => x"11",
          4996 => x"33",
          4997 => x"71",
          4998 => x"59",
          4999 => x"56",
          5000 => x"71",
          5001 => x"33",
          5002 => x"07",
          5003 => x"a2",
          5004 => x"07",
          5005 => x"53",
          5006 => x"53",
          5007 => x"70",
          5008 => x"82",
          5009 => x"70",
          5010 => x"81",
          5011 => x"8b",
          5012 => x"2b",
          5013 => x"57",
          5014 => x"82",
          5015 => x"13",
          5016 => x"2b",
          5017 => x"2a",
          5018 => x"52",
          5019 => x"34",
          5020 => x"34",
          5021 => x"08",
          5022 => x"33",
          5023 => x"71",
          5024 => x"82",
          5025 => x"52",
          5026 => x"0d",
          5027 => x"0d",
          5028 => x"a0",
          5029 => x"2a",
          5030 => x"ff",
          5031 => x"57",
          5032 => x"3f",
          5033 => x"08",
          5034 => x"71",
          5035 => x"33",
          5036 => x"71",
          5037 => x"83",
          5038 => x"11",
          5039 => x"12",
          5040 => x"2b",
          5041 => x"07",
          5042 => x"51",
          5043 => x"55",
          5044 => x"80",
          5045 => x"82",
          5046 => x"75",
          5047 => x"3f",
          5048 => x"84",
          5049 => x"15",
          5050 => x"2b",
          5051 => x"07",
          5052 => x"88",
          5053 => x"55",
          5054 => x"86",
          5055 => x"81",
          5056 => x"75",
          5057 => x"82",
          5058 => x"70",
          5059 => x"33",
          5060 => x"71",
          5061 => x"70",
          5062 => x"57",
          5063 => x"72",
          5064 => x"73",
          5065 => x"82",
          5066 => x"18",
          5067 => x"86",
          5068 => x"0b",
          5069 => x"82",
          5070 => x"53",
          5071 => x"34",
          5072 => x"34",
          5073 => x"08",
          5074 => x"81",
          5075 => x"88",
          5076 => x"82",
          5077 => x"70",
          5078 => x"51",
          5079 => x"74",
          5080 => x"81",
          5081 => x"3d",
          5082 => x"3d",
          5083 => x"82",
          5084 => x"84",
          5085 => x"3f",
          5086 => x"86",
          5087 => x"fe",
          5088 => x"3d",
          5089 => x"3d",
          5090 => x"52",
          5091 => x"3f",
          5092 => x"08",
          5093 => x"06",
          5094 => x"08",
          5095 => x"85",
          5096 => x"88",
          5097 => x"5f",
          5098 => x"5a",
          5099 => x"59",
          5100 => x"80",
          5101 => x"88",
          5102 => x"33",
          5103 => x"71",
          5104 => x"70",
          5105 => x"06",
          5106 => x"83",
          5107 => x"70",
          5108 => x"53",
          5109 => x"55",
          5110 => x"8a",
          5111 => x"2e",
          5112 => x"78",
          5113 => x"15",
          5114 => x"33",
          5115 => x"07",
          5116 => x"c2",
          5117 => x"ff",
          5118 => x"38",
          5119 => x"56",
          5120 => x"2b",
          5121 => x"08",
          5122 => x"81",
          5123 => x"88",
          5124 => x"81",
          5125 => x"51",
          5126 => x"5c",
          5127 => x"2e",
          5128 => x"55",
          5129 => x"78",
          5130 => x"38",
          5131 => x"80",
          5132 => x"38",
          5133 => x"09",
          5134 => x"38",
          5135 => x"f2",
          5136 => x"39",
          5137 => x"53",
          5138 => x"51",
          5139 => x"82",
          5140 => x"70",
          5141 => x"33",
          5142 => x"71",
          5143 => x"83",
          5144 => x"5a",
          5145 => x"05",
          5146 => x"83",
          5147 => x"70",
          5148 => x"59",
          5149 => x"84",
          5150 => x"81",
          5151 => x"76",
          5152 => x"82",
          5153 => x"75",
          5154 => x"11",
          5155 => x"11",
          5156 => x"33",
          5157 => x"07",
          5158 => x"53",
          5159 => x"5a",
          5160 => x"86",
          5161 => x"87",
          5162 => x"b5",
          5163 => x"1c",
          5164 => x"85",
          5165 => x"8b",
          5166 => x"2b",
          5167 => x"5a",
          5168 => x"54",
          5169 => x"34",
          5170 => x"34",
          5171 => x"08",
          5172 => x"1d",
          5173 => x"85",
          5174 => x"88",
          5175 => x"88",
          5176 => x"5f",
          5177 => x"73",
          5178 => x"75",
          5179 => x"82",
          5180 => x"1b",
          5181 => x"73",
          5182 => x"0c",
          5183 => x"04",
          5184 => x"74",
          5185 => x"a0",
          5186 => x"f4",
          5187 => x"53",
          5188 => x"8b",
          5189 => x"fc",
          5190 => x"b5",
          5191 => x"72",
          5192 => x"0c",
          5193 => x"04",
          5194 => x"64",
          5195 => x"80",
          5196 => x"82",
          5197 => x"60",
          5198 => x"06",
          5199 => x"a9",
          5200 => x"38",
          5201 => x"b8",
          5202 => x"a8",
          5203 => x"c7",
          5204 => x"38",
          5205 => x"92",
          5206 => x"83",
          5207 => x"51",
          5208 => x"82",
          5209 => x"83",
          5210 => x"82",
          5211 => x"7d",
          5212 => x"2a",
          5213 => x"ff",
          5214 => x"2b",
          5215 => x"33",
          5216 => x"71",
          5217 => x"70",
          5218 => x"83",
          5219 => x"70",
          5220 => x"05",
          5221 => x"1a",
          5222 => x"12",
          5223 => x"2b",
          5224 => x"2b",
          5225 => x"53",
          5226 => x"5c",
          5227 => x"5c",
          5228 => x"73",
          5229 => x"38",
          5230 => x"ff",
          5231 => x"70",
          5232 => x"06",
          5233 => x"16",
          5234 => x"33",
          5235 => x"07",
          5236 => x"1c",
          5237 => x"12",
          5238 => x"2b",
          5239 => x"07",
          5240 => x"52",
          5241 => x"80",
          5242 => x"78",
          5243 => x"83",
          5244 => x"41",
          5245 => x"27",
          5246 => x"60",
          5247 => x"7b",
          5248 => x"06",
          5249 => x"51",
          5250 => x"7a",
          5251 => x"06",
          5252 => x"39",
          5253 => x"7a",
          5254 => x"38",
          5255 => x"aa",
          5256 => x"39",
          5257 => x"7a",
          5258 => x"c8",
          5259 => x"82",
          5260 => x"12",
          5261 => x"2b",
          5262 => x"54",
          5263 => x"80",
          5264 => x"f7",
          5265 => x"b5",
          5266 => x"ff",
          5267 => x"54",
          5268 => x"83",
          5269 => x"a0",
          5270 => x"05",
          5271 => x"ff",
          5272 => x"82",
          5273 => x"14",
          5274 => x"83",
          5275 => x"59",
          5276 => x"39",
          5277 => x"7a",
          5278 => x"d4",
          5279 => x"f5",
          5280 => x"b5",
          5281 => x"82",
          5282 => x"12",
          5283 => x"2b",
          5284 => x"54",
          5285 => x"80",
          5286 => x"f6",
          5287 => x"b5",
          5288 => x"ff",
          5289 => x"54",
          5290 => x"83",
          5291 => x"a0",
          5292 => x"05",
          5293 => x"ff",
          5294 => x"82",
          5295 => x"14",
          5296 => x"62",
          5297 => x"5c",
          5298 => x"ff",
          5299 => x"39",
          5300 => x"54",
          5301 => x"82",
          5302 => x"5c",
          5303 => x"08",
          5304 => x"38",
          5305 => x"52",
          5306 => x"08",
          5307 => x"96",
          5308 => x"f7",
          5309 => x"58",
          5310 => x"99",
          5311 => x"7a",
          5312 => x"f2",
          5313 => x"19",
          5314 => x"b5",
          5315 => x"84",
          5316 => x"f9",
          5317 => x"73",
          5318 => x"0c",
          5319 => x"04",
          5320 => x"77",
          5321 => x"52",
          5322 => x"3f",
          5323 => x"08",
          5324 => x"a8",
          5325 => x"8e",
          5326 => x"80",
          5327 => x"a8",
          5328 => x"a7",
          5329 => x"82",
          5330 => x"86",
          5331 => x"ff",
          5332 => x"8f",
          5333 => x"81",
          5334 => x"26",
          5335 => x"b5",
          5336 => x"52",
          5337 => x"a8",
          5338 => x"0d",
          5339 => x"0d",
          5340 => x"33",
          5341 => x"9f",
          5342 => x"53",
          5343 => x"81",
          5344 => x"38",
          5345 => x"87",
          5346 => x"11",
          5347 => x"54",
          5348 => x"84",
          5349 => x"54",
          5350 => x"87",
          5351 => x"11",
          5352 => x"0c",
          5353 => x"c0",
          5354 => x"70",
          5355 => x"70",
          5356 => x"51",
          5357 => x"8a",
          5358 => x"98",
          5359 => x"70",
          5360 => x"08",
          5361 => x"06",
          5362 => x"38",
          5363 => x"8c",
          5364 => x"80",
          5365 => x"71",
          5366 => x"14",
          5367 => x"a4",
          5368 => x"70",
          5369 => x"0c",
          5370 => x"04",
          5371 => x"60",
          5372 => x"8c",
          5373 => x"33",
          5374 => x"5b",
          5375 => x"5a",
          5376 => x"82",
          5377 => x"81",
          5378 => x"52",
          5379 => x"38",
          5380 => x"84",
          5381 => x"92",
          5382 => x"c0",
          5383 => x"87",
          5384 => x"13",
          5385 => x"57",
          5386 => x"0b",
          5387 => x"8c",
          5388 => x"0c",
          5389 => x"75",
          5390 => x"2a",
          5391 => x"51",
          5392 => x"80",
          5393 => x"7b",
          5394 => x"7b",
          5395 => x"5d",
          5396 => x"59",
          5397 => x"06",
          5398 => x"73",
          5399 => x"81",
          5400 => x"ff",
          5401 => x"72",
          5402 => x"38",
          5403 => x"8c",
          5404 => x"c3",
          5405 => x"98",
          5406 => x"71",
          5407 => x"38",
          5408 => x"2e",
          5409 => x"76",
          5410 => x"92",
          5411 => x"72",
          5412 => x"06",
          5413 => x"f7",
          5414 => x"5a",
          5415 => x"80",
          5416 => x"70",
          5417 => x"5a",
          5418 => x"80",
          5419 => x"73",
          5420 => x"06",
          5421 => x"38",
          5422 => x"fe",
          5423 => x"fc",
          5424 => x"52",
          5425 => x"83",
          5426 => x"71",
          5427 => x"b5",
          5428 => x"3d",
          5429 => x"3d",
          5430 => x"64",
          5431 => x"bf",
          5432 => x"40",
          5433 => x"59",
          5434 => x"58",
          5435 => x"82",
          5436 => x"81",
          5437 => x"52",
          5438 => x"09",
          5439 => x"b1",
          5440 => x"84",
          5441 => x"92",
          5442 => x"c0",
          5443 => x"87",
          5444 => x"13",
          5445 => x"56",
          5446 => x"87",
          5447 => x"0c",
          5448 => x"82",
          5449 => x"58",
          5450 => x"84",
          5451 => x"06",
          5452 => x"71",
          5453 => x"38",
          5454 => x"05",
          5455 => x"0c",
          5456 => x"73",
          5457 => x"81",
          5458 => x"71",
          5459 => x"38",
          5460 => x"8c",
          5461 => x"d0",
          5462 => x"98",
          5463 => x"71",
          5464 => x"38",
          5465 => x"2e",
          5466 => x"76",
          5467 => x"92",
          5468 => x"72",
          5469 => x"06",
          5470 => x"f7",
          5471 => x"59",
          5472 => x"1a",
          5473 => x"06",
          5474 => x"59",
          5475 => x"80",
          5476 => x"73",
          5477 => x"06",
          5478 => x"38",
          5479 => x"fe",
          5480 => x"fc",
          5481 => x"52",
          5482 => x"83",
          5483 => x"71",
          5484 => x"b5",
          5485 => x"3d",
          5486 => x"3d",
          5487 => x"84",
          5488 => x"33",
          5489 => x"a7",
          5490 => x"54",
          5491 => x"fa",
          5492 => x"b5",
          5493 => x"06",
          5494 => x"72",
          5495 => x"85",
          5496 => x"98",
          5497 => x"56",
          5498 => x"80",
          5499 => x"76",
          5500 => x"74",
          5501 => x"c0",
          5502 => x"54",
          5503 => x"2e",
          5504 => x"d4",
          5505 => x"2e",
          5506 => x"80",
          5507 => x"08",
          5508 => x"70",
          5509 => x"51",
          5510 => x"2e",
          5511 => x"c0",
          5512 => x"52",
          5513 => x"87",
          5514 => x"08",
          5515 => x"38",
          5516 => x"87",
          5517 => x"14",
          5518 => x"70",
          5519 => x"52",
          5520 => x"96",
          5521 => x"92",
          5522 => x"0a",
          5523 => x"39",
          5524 => x"0c",
          5525 => x"39",
          5526 => x"54",
          5527 => x"a8",
          5528 => x"0d",
          5529 => x"0d",
          5530 => x"33",
          5531 => x"88",
          5532 => x"b5",
          5533 => x"51",
          5534 => x"04",
          5535 => x"75",
          5536 => x"82",
          5537 => x"90",
          5538 => x"2b",
          5539 => x"33",
          5540 => x"88",
          5541 => x"71",
          5542 => x"a8",
          5543 => x"54",
          5544 => x"85",
          5545 => x"ff",
          5546 => x"02",
          5547 => x"05",
          5548 => x"70",
          5549 => x"05",
          5550 => x"88",
          5551 => x"72",
          5552 => x"0d",
          5553 => x"0d",
          5554 => x"52",
          5555 => x"81",
          5556 => x"70",
          5557 => x"70",
          5558 => x"05",
          5559 => x"88",
          5560 => x"72",
          5561 => x"54",
          5562 => x"2a",
          5563 => x"34",
          5564 => x"04",
          5565 => x"76",
          5566 => x"54",
          5567 => x"2e",
          5568 => x"70",
          5569 => x"33",
          5570 => x"05",
          5571 => x"11",
          5572 => x"84",
          5573 => x"fe",
          5574 => x"77",
          5575 => x"53",
          5576 => x"81",
          5577 => x"ff",
          5578 => x"f4",
          5579 => x"0d",
          5580 => x"0d",
          5581 => x"56",
          5582 => x"70",
          5583 => x"33",
          5584 => x"05",
          5585 => x"71",
          5586 => x"56",
          5587 => x"72",
          5588 => x"38",
          5589 => x"e2",
          5590 => x"b5",
          5591 => x"3d",
          5592 => x"3d",
          5593 => x"54",
          5594 => x"71",
          5595 => x"38",
          5596 => x"70",
          5597 => x"f3",
          5598 => x"82",
          5599 => x"84",
          5600 => x"80",
          5601 => x"a8",
          5602 => x"0b",
          5603 => x"0c",
          5604 => x"0d",
          5605 => x"0b",
          5606 => x"56",
          5607 => x"2e",
          5608 => x"81",
          5609 => x"08",
          5610 => x"70",
          5611 => x"33",
          5612 => x"a2",
          5613 => x"a8",
          5614 => x"09",
          5615 => x"38",
          5616 => x"08",
          5617 => x"b0",
          5618 => x"a4",
          5619 => x"9c",
          5620 => x"56",
          5621 => x"27",
          5622 => x"16",
          5623 => x"82",
          5624 => x"06",
          5625 => x"54",
          5626 => x"78",
          5627 => x"33",
          5628 => x"3f",
          5629 => x"5a",
          5630 => x"a8",
          5631 => x"0d",
          5632 => x"0d",
          5633 => x"56",
          5634 => x"b0",
          5635 => x"af",
          5636 => x"fe",
          5637 => x"b5",
          5638 => x"82",
          5639 => x"9f",
          5640 => x"74",
          5641 => x"52",
          5642 => x"51",
          5643 => x"82",
          5644 => x"80",
          5645 => x"ff",
          5646 => x"74",
          5647 => x"76",
          5648 => x"0c",
          5649 => x"04",
          5650 => x"7a",
          5651 => x"fe",
          5652 => x"b5",
          5653 => x"82",
          5654 => x"81",
          5655 => x"33",
          5656 => x"2e",
          5657 => x"80",
          5658 => x"17",
          5659 => x"81",
          5660 => x"06",
          5661 => x"84",
          5662 => x"b5",
          5663 => x"b4",
          5664 => x"56",
          5665 => x"82",
          5666 => x"84",
          5667 => x"fc",
          5668 => x"8b",
          5669 => x"52",
          5670 => x"a9",
          5671 => x"85",
          5672 => x"84",
          5673 => x"fc",
          5674 => x"17",
          5675 => x"9c",
          5676 => x"91",
          5677 => x"08",
          5678 => x"17",
          5679 => x"3f",
          5680 => x"81",
          5681 => x"19",
          5682 => x"53",
          5683 => x"17",
          5684 => x"82",
          5685 => x"18",
          5686 => x"80",
          5687 => x"33",
          5688 => x"3f",
          5689 => x"08",
          5690 => x"38",
          5691 => x"82",
          5692 => x"8a",
          5693 => x"fb",
          5694 => x"fe",
          5695 => x"08",
          5696 => x"56",
          5697 => x"74",
          5698 => x"38",
          5699 => x"75",
          5700 => x"16",
          5701 => x"53",
          5702 => x"a8",
          5703 => x"0d",
          5704 => x"0d",
          5705 => x"08",
          5706 => x"81",
          5707 => x"df",
          5708 => x"15",
          5709 => x"d7",
          5710 => x"33",
          5711 => x"82",
          5712 => x"38",
          5713 => x"89",
          5714 => x"2e",
          5715 => x"bf",
          5716 => x"2e",
          5717 => x"81",
          5718 => x"81",
          5719 => x"89",
          5720 => x"08",
          5721 => x"52",
          5722 => x"3f",
          5723 => x"08",
          5724 => x"74",
          5725 => x"14",
          5726 => x"81",
          5727 => x"2a",
          5728 => x"05",
          5729 => x"57",
          5730 => x"f5",
          5731 => x"a8",
          5732 => x"38",
          5733 => x"06",
          5734 => x"33",
          5735 => x"78",
          5736 => x"06",
          5737 => x"5c",
          5738 => x"53",
          5739 => x"38",
          5740 => x"06",
          5741 => x"39",
          5742 => x"a4",
          5743 => x"52",
          5744 => x"bd",
          5745 => x"a8",
          5746 => x"38",
          5747 => x"fe",
          5748 => x"b4",
          5749 => x"8d",
          5750 => x"a8",
          5751 => x"ff",
          5752 => x"39",
          5753 => x"a4",
          5754 => x"52",
          5755 => x"91",
          5756 => x"a8",
          5757 => x"76",
          5758 => x"fc",
          5759 => x"b4",
          5760 => x"f8",
          5761 => x"a8",
          5762 => x"06",
          5763 => x"81",
          5764 => x"b5",
          5765 => x"3d",
          5766 => x"3d",
          5767 => x"7e",
          5768 => x"82",
          5769 => x"27",
          5770 => x"76",
          5771 => x"27",
          5772 => x"75",
          5773 => x"79",
          5774 => x"38",
          5775 => x"89",
          5776 => x"2e",
          5777 => x"80",
          5778 => x"2e",
          5779 => x"81",
          5780 => x"81",
          5781 => x"89",
          5782 => x"08",
          5783 => x"52",
          5784 => x"3f",
          5785 => x"08",
          5786 => x"a8",
          5787 => x"38",
          5788 => x"06",
          5789 => x"81",
          5790 => x"06",
          5791 => x"77",
          5792 => x"2e",
          5793 => x"84",
          5794 => x"06",
          5795 => x"06",
          5796 => x"53",
          5797 => x"81",
          5798 => x"34",
          5799 => x"a4",
          5800 => x"52",
          5801 => x"d9",
          5802 => x"a8",
          5803 => x"b5",
          5804 => x"94",
          5805 => x"ff",
          5806 => x"05",
          5807 => x"54",
          5808 => x"38",
          5809 => x"74",
          5810 => x"06",
          5811 => x"07",
          5812 => x"74",
          5813 => x"39",
          5814 => x"a4",
          5815 => x"52",
          5816 => x"9d",
          5817 => x"a8",
          5818 => x"b5",
          5819 => x"d8",
          5820 => x"ff",
          5821 => x"76",
          5822 => x"06",
          5823 => x"05",
          5824 => x"3f",
          5825 => x"87",
          5826 => x"08",
          5827 => x"51",
          5828 => x"82",
          5829 => x"59",
          5830 => x"08",
          5831 => x"f0",
          5832 => x"82",
          5833 => x"06",
          5834 => x"05",
          5835 => x"54",
          5836 => x"3f",
          5837 => x"08",
          5838 => x"74",
          5839 => x"51",
          5840 => x"81",
          5841 => x"34",
          5842 => x"a8",
          5843 => x"0d",
          5844 => x"0d",
          5845 => x"72",
          5846 => x"56",
          5847 => x"27",
          5848 => x"98",
          5849 => x"9d",
          5850 => x"2e",
          5851 => x"53",
          5852 => x"51",
          5853 => x"82",
          5854 => x"54",
          5855 => x"08",
          5856 => x"93",
          5857 => x"80",
          5858 => x"54",
          5859 => x"82",
          5860 => x"54",
          5861 => x"74",
          5862 => x"fb",
          5863 => x"b5",
          5864 => x"82",
          5865 => x"80",
          5866 => x"38",
          5867 => x"08",
          5868 => x"38",
          5869 => x"08",
          5870 => x"38",
          5871 => x"52",
          5872 => x"d6",
          5873 => x"a8",
          5874 => x"98",
          5875 => x"11",
          5876 => x"57",
          5877 => x"74",
          5878 => x"81",
          5879 => x"0c",
          5880 => x"81",
          5881 => x"84",
          5882 => x"55",
          5883 => x"ff",
          5884 => x"54",
          5885 => x"a8",
          5886 => x"0d",
          5887 => x"0d",
          5888 => x"08",
          5889 => x"79",
          5890 => x"17",
          5891 => x"80",
          5892 => x"98",
          5893 => x"26",
          5894 => x"58",
          5895 => x"52",
          5896 => x"fd",
          5897 => x"74",
          5898 => x"08",
          5899 => x"38",
          5900 => x"08",
          5901 => x"a8",
          5902 => x"82",
          5903 => x"17",
          5904 => x"a8",
          5905 => x"c7",
          5906 => x"90",
          5907 => x"56",
          5908 => x"2e",
          5909 => x"77",
          5910 => x"81",
          5911 => x"38",
          5912 => x"98",
          5913 => x"26",
          5914 => x"56",
          5915 => x"51",
          5916 => x"80",
          5917 => x"a8",
          5918 => x"09",
          5919 => x"38",
          5920 => x"08",
          5921 => x"a8",
          5922 => x"30",
          5923 => x"80",
          5924 => x"07",
          5925 => x"08",
          5926 => x"55",
          5927 => x"ef",
          5928 => x"a8",
          5929 => x"95",
          5930 => x"08",
          5931 => x"27",
          5932 => x"98",
          5933 => x"89",
          5934 => x"85",
          5935 => x"db",
          5936 => x"81",
          5937 => x"17",
          5938 => x"89",
          5939 => x"75",
          5940 => x"ac",
          5941 => x"7a",
          5942 => x"3f",
          5943 => x"08",
          5944 => x"38",
          5945 => x"b5",
          5946 => x"2e",
          5947 => x"86",
          5948 => x"a8",
          5949 => x"b5",
          5950 => x"70",
          5951 => x"07",
          5952 => x"7c",
          5953 => x"55",
          5954 => x"f8",
          5955 => x"2e",
          5956 => x"ff",
          5957 => x"55",
          5958 => x"ff",
          5959 => x"76",
          5960 => x"3f",
          5961 => x"08",
          5962 => x"08",
          5963 => x"b5",
          5964 => x"80",
          5965 => x"55",
          5966 => x"94",
          5967 => x"2e",
          5968 => x"53",
          5969 => x"51",
          5970 => x"82",
          5971 => x"55",
          5972 => x"75",
          5973 => x"98",
          5974 => x"05",
          5975 => x"56",
          5976 => x"26",
          5977 => x"15",
          5978 => x"84",
          5979 => x"07",
          5980 => x"18",
          5981 => x"ff",
          5982 => x"2e",
          5983 => x"39",
          5984 => x"39",
          5985 => x"08",
          5986 => x"81",
          5987 => x"74",
          5988 => x"0c",
          5989 => x"04",
          5990 => x"7a",
          5991 => x"f3",
          5992 => x"b5",
          5993 => x"81",
          5994 => x"a8",
          5995 => x"38",
          5996 => x"51",
          5997 => x"82",
          5998 => x"82",
          5999 => x"b0",
          6000 => x"84",
          6001 => x"52",
          6002 => x"52",
          6003 => x"3f",
          6004 => x"39",
          6005 => x"8a",
          6006 => x"75",
          6007 => x"38",
          6008 => x"19",
          6009 => x"81",
          6010 => x"ed",
          6011 => x"b5",
          6012 => x"2e",
          6013 => x"15",
          6014 => x"70",
          6015 => x"07",
          6016 => x"53",
          6017 => x"75",
          6018 => x"0c",
          6019 => x"04",
          6020 => x"7a",
          6021 => x"58",
          6022 => x"f0",
          6023 => x"80",
          6024 => x"9f",
          6025 => x"80",
          6026 => x"90",
          6027 => x"17",
          6028 => x"aa",
          6029 => x"53",
          6030 => x"88",
          6031 => x"08",
          6032 => x"38",
          6033 => x"53",
          6034 => x"17",
          6035 => x"72",
          6036 => x"fe",
          6037 => x"08",
          6038 => x"80",
          6039 => x"16",
          6040 => x"2b",
          6041 => x"75",
          6042 => x"73",
          6043 => x"f5",
          6044 => x"b5",
          6045 => x"82",
          6046 => x"ff",
          6047 => x"81",
          6048 => x"a8",
          6049 => x"38",
          6050 => x"82",
          6051 => x"26",
          6052 => x"58",
          6053 => x"73",
          6054 => x"39",
          6055 => x"51",
          6056 => x"82",
          6057 => x"98",
          6058 => x"94",
          6059 => x"17",
          6060 => x"58",
          6061 => x"9a",
          6062 => x"81",
          6063 => x"74",
          6064 => x"98",
          6065 => x"83",
          6066 => x"b4",
          6067 => x"0c",
          6068 => x"82",
          6069 => x"8a",
          6070 => x"f8",
          6071 => x"70",
          6072 => x"08",
          6073 => x"57",
          6074 => x"0a",
          6075 => x"38",
          6076 => x"15",
          6077 => x"08",
          6078 => x"72",
          6079 => x"cb",
          6080 => x"ff",
          6081 => x"81",
          6082 => x"13",
          6083 => x"94",
          6084 => x"74",
          6085 => x"85",
          6086 => x"22",
          6087 => x"73",
          6088 => x"38",
          6089 => x"8a",
          6090 => x"05",
          6091 => x"06",
          6092 => x"8a",
          6093 => x"73",
          6094 => x"3f",
          6095 => x"08",
          6096 => x"81",
          6097 => x"a8",
          6098 => x"ff",
          6099 => x"82",
          6100 => x"ff",
          6101 => x"38",
          6102 => x"82",
          6103 => x"26",
          6104 => x"7b",
          6105 => x"98",
          6106 => x"55",
          6107 => x"94",
          6108 => x"73",
          6109 => x"3f",
          6110 => x"08",
          6111 => x"82",
          6112 => x"80",
          6113 => x"38",
          6114 => x"b5",
          6115 => x"2e",
          6116 => x"55",
          6117 => x"08",
          6118 => x"38",
          6119 => x"08",
          6120 => x"fb",
          6121 => x"b5",
          6122 => x"38",
          6123 => x"0c",
          6124 => x"51",
          6125 => x"82",
          6126 => x"98",
          6127 => x"90",
          6128 => x"16",
          6129 => x"15",
          6130 => x"74",
          6131 => x"0c",
          6132 => x"04",
          6133 => x"7b",
          6134 => x"5b",
          6135 => x"52",
          6136 => x"ac",
          6137 => x"a8",
          6138 => x"b5",
          6139 => x"ec",
          6140 => x"a8",
          6141 => x"17",
          6142 => x"51",
          6143 => x"82",
          6144 => x"54",
          6145 => x"08",
          6146 => x"82",
          6147 => x"9c",
          6148 => x"33",
          6149 => x"72",
          6150 => x"09",
          6151 => x"38",
          6152 => x"b5",
          6153 => x"72",
          6154 => x"55",
          6155 => x"53",
          6156 => x"8e",
          6157 => x"56",
          6158 => x"09",
          6159 => x"38",
          6160 => x"b5",
          6161 => x"81",
          6162 => x"fd",
          6163 => x"b5",
          6164 => x"82",
          6165 => x"80",
          6166 => x"38",
          6167 => x"09",
          6168 => x"38",
          6169 => x"82",
          6170 => x"8b",
          6171 => x"fd",
          6172 => x"9a",
          6173 => x"eb",
          6174 => x"b5",
          6175 => x"ff",
          6176 => x"70",
          6177 => x"53",
          6178 => x"09",
          6179 => x"38",
          6180 => x"eb",
          6181 => x"b5",
          6182 => x"2b",
          6183 => x"72",
          6184 => x"0c",
          6185 => x"04",
          6186 => x"77",
          6187 => x"ff",
          6188 => x"9a",
          6189 => x"55",
          6190 => x"76",
          6191 => x"53",
          6192 => x"09",
          6193 => x"38",
          6194 => x"52",
          6195 => x"eb",
          6196 => x"3d",
          6197 => x"3d",
          6198 => x"5b",
          6199 => x"08",
          6200 => x"15",
          6201 => x"81",
          6202 => x"15",
          6203 => x"51",
          6204 => x"82",
          6205 => x"58",
          6206 => x"08",
          6207 => x"9c",
          6208 => x"33",
          6209 => x"86",
          6210 => x"80",
          6211 => x"13",
          6212 => x"06",
          6213 => x"06",
          6214 => x"72",
          6215 => x"82",
          6216 => x"53",
          6217 => x"2e",
          6218 => x"53",
          6219 => x"a9",
          6220 => x"74",
          6221 => x"72",
          6222 => x"38",
          6223 => x"99",
          6224 => x"a8",
          6225 => x"06",
          6226 => x"88",
          6227 => x"06",
          6228 => x"54",
          6229 => x"a0",
          6230 => x"74",
          6231 => x"3f",
          6232 => x"08",
          6233 => x"a8",
          6234 => x"98",
          6235 => x"fa",
          6236 => x"80",
          6237 => x"0c",
          6238 => x"a8",
          6239 => x"0d",
          6240 => x"0d",
          6241 => x"57",
          6242 => x"73",
          6243 => x"3f",
          6244 => x"08",
          6245 => x"a8",
          6246 => x"98",
          6247 => x"75",
          6248 => x"3f",
          6249 => x"08",
          6250 => x"a8",
          6251 => x"a0",
          6252 => x"a8",
          6253 => x"14",
          6254 => x"db",
          6255 => x"a0",
          6256 => x"14",
          6257 => x"ac",
          6258 => x"83",
          6259 => x"82",
          6260 => x"87",
          6261 => x"fd",
          6262 => x"70",
          6263 => x"08",
          6264 => x"55",
          6265 => x"3f",
          6266 => x"08",
          6267 => x"13",
          6268 => x"73",
          6269 => x"83",
          6270 => x"3d",
          6271 => x"3d",
          6272 => x"57",
          6273 => x"89",
          6274 => x"17",
          6275 => x"81",
          6276 => x"70",
          6277 => x"55",
          6278 => x"08",
          6279 => x"81",
          6280 => x"52",
          6281 => x"a8",
          6282 => x"2e",
          6283 => x"84",
          6284 => x"52",
          6285 => x"09",
          6286 => x"38",
          6287 => x"81",
          6288 => x"81",
          6289 => x"73",
          6290 => x"55",
          6291 => x"55",
          6292 => x"c5",
          6293 => x"88",
          6294 => x"0b",
          6295 => x"9c",
          6296 => x"8b",
          6297 => x"17",
          6298 => x"08",
          6299 => x"52",
          6300 => x"82",
          6301 => x"76",
          6302 => x"51",
          6303 => x"82",
          6304 => x"86",
          6305 => x"12",
          6306 => x"3f",
          6307 => x"08",
          6308 => x"88",
          6309 => x"f3",
          6310 => x"70",
          6311 => x"80",
          6312 => x"51",
          6313 => x"af",
          6314 => x"81",
          6315 => x"dc",
          6316 => x"74",
          6317 => x"38",
          6318 => x"88",
          6319 => x"39",
          6320 => x"80",
          6321 => x"56",
          6322 => x"af",
          6323 => x"06",
          6324 => x"56",
          6325 => x"32",
          6326 => x"80",
          6327 => x"51",
          6328 => x"dc",
          6329 => x"1c",
          6330 => x"33",
          6331 => x"9f",
          6332 => x"ff",
          6333 => x"1c",
          6334 => x"7a",
          6335 => x"3f",
          6336 => x"08",
          6337 => x"39",
          6338 => x"a0",
          6339 => x"5e",
          6340 => x"52",
          6341 => x"ff",
          6342 => x"59",
          6343 => x"33",
          6344 => x"ae",
          6345 => x"06",
          6346 => x"78",
          6347 => x"81",
          6348 => x"32",
          6349 => x"9f",
          6350 => x"26",
          6351 => x"53",
          6352 => x"73",
          6353 => x"17",
          6354 => x"34",
          6355 => x"db",
          6356 => x"32",
          6357 => x"9f",
          6358 => x"54",
          6359 => x"2e",
          6360 => x"80",
          6361 => x"75",
          6362 => x"bd",
          6363 => x"7e",
          6364 => x"a0",
          6365 => x"bd",
          6366 => x"82",
          6367 => x"18",
          6368 => x"1a",
          6369 => x"a0",
          6370 => x"fc",
          6371 => x"32",
          6372 => x"80",
          6373 => x"30",
          6374 => x"71",
          6375 => x"51",
          6376 => x"55",
          6377 => x"ac",
          6378 => x"81",
          6379 => x"78",
          6380 => x"51",
          6381 => x"af",
          6382 => x"06",
          6383 => x"55",
          6384 => x"32",
          6385 => x"80",
          6386 => x"51",
          6387 => x"db",
          6388 => x"39",
          6389 => x"09",
          6390 => x"38",
          6391 => x"7c",
          6392 => x"54",
          6393 => x"a2",
          6394 => x"32",
          6395 => x"ae",
          6396 => x"72",
          6397 => x"9f",
          6398 => x"51",
          6399 => x"74",
          6400 => x"88",
          6401 => x"fe",
          6402 => x"98",
          6403 => x"80",
          6404 => x"75",
          6405 => x"82",
          6406 => x"33",
          6407 => x"51",
          6408 => x"82",
          6409 => x"80",
          6410 => x"78",
          6411 => x"81",
          6412 => x"5a",
          6413 => x"d2",
          6414 => x"a8",
          6415 => x"80",
          6416 => x"1c",
          6417 => x"27",
          6418 => x"79",
          6419 => x"74",
          6420 => x"7a",
          6421 => x"74",
          6422 => x"39",
          6423 => x"ae",
          6424 => x"fe",
          6425 => x"a8",
          6426 => x"ff",
          6427 => x"73",
          6428 => x"38",
          6429 => x"81",
          6430 => x"54",
          6431 => x"75",
          6432 => x"17",
          6433 => x"39",
          6434 => x"0c",
          6435 => x"99",
          6436 => x"54",
          6437 => x"2e",
          6438 => x"84",
          6439 => x"34",
          6440 => x"76",
          6441 => x"8b",
          6442 => x"81",
          6443 => x"56",
          6444 => x"80",
          6445 => x"1b",
          6446 => x"08",
          6447 => x"51",
          6448 => x"82",
          6449 => x"56",
          6450 => x"08",
          6451 => x"98",
          6452 => x"76",
          6453 => x"3f",
          6454 => x"08",
          6455 => x"a8",
          6456 => x"38",
          6457 => x"70",
          6458 => x"73",
          6459 => x"be",
          6460 => x"33",
          6461 => x"73",
          6462 => x"8b",
          6463 => x"83",
          6464 => x"06",
          6465 => x"73",
          6466 => x"53",
          6467 => x"51",
          6468 => x"82",
          6469 => x"80",
          6470 => x"75",
          6471 => x"f3",
          6472 => x"9f",
          6473 => x"1c",
          6474 => x"74",
          6475 => x"38",
          6476 => x"09",
          6477 => x"e7",
          6478 => x"2a",
          6479 => x"77",
          6480 => x"51",
          6481 => x"2e",
          6482 => x"81",
          6483 => x"80",
          6484 => x"38",
          6485 => x"ab",
          6486 => x"55",
          6487 => x"75",
          6488 => x"73",
          6489 => x"55",
          6490 => x"82",
          6491 => x"06",
          6492 => x"ab",
          6493 => x"33",
          6494 => x"70",
          6495 => x"55",
          6496 => x"2e",
          6497 => x"1b",
          6498 => x"06",
          6499 => x"52",
          6500 => x"db",
          6501 => x"a8",
          6502 => x"0c",
          6503 => x"74",
          6504 => x"0c",
          6505 => x"04",
          6506 => x"7c",
          6507 => x"08",
          6508 => x"55",
          6509 => x"59",
          6510 => x"81",
          6511 => x"70",
          6512 => x"33",
          6513 => x"52",
          6514 => x"2e",
          6515 => x"ee",
          6516 => x"2e",
          6517 => x"81",
          6518 => x"33",
          6519 => x"81",
          6520 => x"52",
          6521 => x"26",
          6522 => x"14",
          6523 => x"06",
          6524 => x"52",
          6525 => x"80",
          6526 => x"0b",
          6527 => x"59",
          6528 => x"7a",
          6529 => x"70",
          6530 => x"33",
          6531 => x"05",
          6532 => x"9f",
          6533 => x"53",
          6534 => x"89",
          6535 => x"70",
          6536 => x"54",
          6537 => x"12",
          6538 => x"26",
          6539 => x"12",
          6540 => x"06",
          6541 => x"30",
          6542 => x"51",
          6543 => x"2e",
          6544 => x"85",
          6545 => x"be",
          6546 => x"74",
          6547 => x"30",
          6548 => x"9f",
          6549 => x"2a",
          6550 => x"54",
          6551 => x"2e",
          6552 => x"15",
          6553 => x"55",
          6554 => x"ff",
          6555 => x"39",
          6556 => x"86",
          6557 => x"7c",
          6558 => x"51",
          6559 => x"cc",
          6560 => x"70",
          6561 => x"0c",
          6562 => x"04",
          6563 => x"78",
          6564 => x"83",
          6565 => x"0b",
          6566 => x"79",
          6567 => x"e2",
          6568 => x"55",
          6569 => x"08",
          6570 => x"84",
          6571 => x"df",
          6572 => x"b5",
          6573 => x"ff",
          6574 => x"83",
          6575 => x"d4",
          6576 => x"81",
          6577 => x"38",
          6578 => x"17",
          6579 => x"74",
          6580 => x"09",
          6581 => x"38",
          6582 => x"81",
          6583 => x"30",
          6584 => x"79",
          6585 => x"54",
          6586 => x"74",
          6587 => x"09",
          6588 => x"38",
          6589 => x"ae",
          6590 => x"ea",
          6591 => x"b1",
          6592 => x"a8",
          6593 => x"b5",
          6594 => x"2e",
          6595 => x"53",
          6596 => x"52",
          6597 => x"51",
          6598 => x"82",
          6599 => x"55",
          6600 => x"08",
          6601 => x"38",
          6602 => x"82",
          6603 => x"88",
          6604 => x"f2",
          6605 => x"02",
          6606 => x"cb",
          6607 => x"55",
          6608 => x"60",
          6609 => x"3f",
          6610 => x"08",
          6611 => x"80",
          6612 => x"a8",
          6613 => x"fc",
          6614 => x"a8",
          6615 => x"82",
          6616 => x"70",
          6617 => x"8c",
          6618 => x"2e",
          6619 => x"73",
          6620 => x"81",
          6621 => x"33",
          6622 => x"80",
          6623 => x"81",
          6624 => x"d7",
          6625 => x"b5",
          6626 => x"ff",
          6627 => x"06",
          6628 => x"98",
          6629 => x"2e",
          6630 => x"74",
          6631 => x"81",
          6632 => x"8a",
          6633 => x"ac",
          6634 => x"39",
          6635 => x"77",
          6636 => x"81",
          6637 => x"33",
          6638 => x"3f",
          6639 => x"08",
          6640 => x"70",
          6641 => x"55",
          6642 => x"86",
          6643 => x"80",
          6644 => x"74",
          6645 => x"81",
          6646 => x"8a",
          6647 => x"f4",
          6648 => x"53",
          6649 => x"fd",
          6650 => x"b5",
          6651 => x"ff",
          6652 => x"82",
          6653 => x"06",
          6654 => x"8c",
          6655 => x"58",
          6656 => x"f6",
          6657 => x"58",
          6658 => x"2e",
          6659 => x"fa",
          6660 => x"e8",
          6661 => x"a8",
          6662 => x"78",
          6663 => x"5a",
          6664 => x"90",
          6665 => x"75",
          6666 => x"38",
          6667 => x"3d",
          6668 => x"70",
          6669 => x"08",
          6670 => x"7a",
          6671 => x"38",
          6672 => x"51",
          6673 => x"82",
          6674 => x"81",
          6675 => x"81",
          6676 => x"38",
          6677 => x"83",
          6678 => x"38",
          6679 => x"84",
          6680 => x"38",
          6681 => x"81",
          6682 => x"38",
          6683 => x"db",
          6684 => x"b5",
          6685 => x"ff",
          6686 => x"72",
          6687 => x"09",
          6688 => x"d0",
          6689 => x"14",
          6690 => x"3f",
          6691 => x"08",
          6692 => x"06",
          6693 => x"38",
          6694 => x"51",
          6695 => x"82",
          6696 => x"58",
          6697 => x"0c",
          6698 => x"33",
          6699 => x"80",
          6700 => x"ff",
          6701 => x"ff",
          6702 => x"55",
          6703 => x"81",
          6704 => x"38",
          6705 => x"06",
          6706 => x"80",
          6707 => x"52",
          6708 => x"8a",
          6709 => x"80",
          6710 => x"ff",
          6711 => x"53",
          6712 => x"86",
          6713 => x"83",
          6714 => x"c5",
          6715 => x"f5",
          6716 => x"a8",
          6717 => x"b5",
          6718 => x"15",
          6719 => x"06",
          6720 => x"76",
          6721 => x"80",
          6722 => x"da",
          6723 => x"b5",
          6724 => x"ff",
          6725 => x"74",
          6726 => x"d4",
          6727 => x"dc",
          6728 => x"a8",
          6729 => x"c2",
          6730 => x"b9",
          6731 => x"a8",
          6732 => x"ff",
          6733 => x"56",
          6734 => x"83",
          6735 => x"14",
          6736 => x"71",
          6737 => x"5a",
          6738 => x"26",
          6739 => x"8a",
          6740 => x"74",
          6741 => x"fe",
          6742 => x"82",
          6743 => x"55",
          6744 => x"08",
          6745 => x"ec",
          6746 => x"a8",
          6747 => x"ff",
          6748 => x"83",
          6749 => x"74",
          6750 => x"26",
          6751 => x"57",
          6752 => x"26",
          6753 => x"57",
          6754 => x"56",
          6755 => x"82",
          6756 => x"15",
          6757 => x"0c",
          6758 => x"0c",
          6759 => x"a4",
          6760 => x"1d",
          6761 => x"54",
          6762 => x"2e",
          6763 => x"af",
          6764 => x"14",
          6765 => x"3f",
          6766 => x"08",
          6767 => x"06",
          6768 => x"72",
          6769 => x"79",
          6770 => x"80",
          6771 => x"d9",
          6772 => x"b5",
          6773 => x"15",
          6774 => x"2b",
          6775 => x"8d",
          6776 => x"2e",
          6777 => x"77",
          6778 => x"0c",
          6779 => x"76",
          6780 => x"38",
          6781 => x"70",
          6782 => x"81",
          6783 => x"53",
          6784 => x"89",
          6785 => x"56",
          6786 => x"08",
          6787 => x"38",
          6788 => x"15",
          6789 => x"8c",
          6790 => x"80",
          6791 => x"34",
          6792 => x"09",
          6793 => x"92",
          6794 => x"14",
          6795 => x"3f",
          6796 => x"08",
          6797 => x"06",
          6798 => x"2e",
          6799 => x"80",
          6800 => x"1b",
          6801 => x"db",
          6802 => x"b5",
          6803 => x"ea",
          6804 => x"a8",
          6805 => x"34",
          6806 => x"51",
          6807 => x"82",
          6808 => x"83",
          6809 => x"53",
          6810 => x"d5",
          6811 => x"06",
          6812 => x"b4",
          6813 => x"84",
          6814 => x"a8",
          6815 => x"85",
          6816 => x"09",
          6817 => x"38",
          6818 => x"51",
          6819 => x"82",
          6820 => x"86",
          6821 => x"f2",
          6822 => x"06",
          6823 => x"9c",
          6824 => x"d8",
          6825 => x"a8",
          6826 => x"0c",
          6827 => x"51",
          6828 => x"82",
          6829 => x"8c",
          6830 => x"74",
          6831 => x"f0",
          6832 => x"53",
          6833 => x"f0",
          6834 => x"15",
          6835 => x"94",
          6836 => x"56",
          6837 => x"a8",
          6838 => x"0d",
          6839 => x"0d",
          6840 => x"55",
          6841 => x"b9",
          6842 => x"53",
          6843 => x"b1",
          6844 => x"52",
          6845 => x"a9",
          6846 => x"22",
          6847 => x"57",
          6848 => x"2e",
          6849 => x"99",
          6850 => x"33",
          6851 => x"3f",
          6852 => x"08",
          6853 => x"71",
          6854 => x"74",
          6855 => x"83",
          6856 => x"78",
          6857 => x"52",
          6858 => x"a8",
          6859 => x"0d",
          6860 => x"0d",
          6861 => x"33",
          6862 => x"3d",
          6863 => x"56",
          6864 => x"8b",
          6865 => x"82",
          6866 => x"24",
          6867 => x"b5",
          6868 => x"29",
          6869 => x"05",
          6870 => x"55",
          6871 => x"84",
          6872 => x"34",
          6873 => x"80",
          6874 => x"80",
          6875 => x"75",
          6876 => x"75",
          6877 => x"38",
          6878 => x"3d",
          6879 => x"05",
          6880 => x"3f",
          6881 => x"08",
          6882 => x"b5",
          6883 => x"3d",
          6884 => x"3d",
          6885 => x"84",
          6886 => x"05",
          6887 => x"89",
          6888 => x"2e",
          6889 => x"77",
          6890 => x"54",
          6891 => x"05",
          6892 => x"84",
          6893 => x"f6",
          6894 => x"b5",
          6895 => x"82",
          6896 => x"84",
          6897 => x"5c",
          6898 => x"3d",
          6899 => x"ed",
          6900 => x"b5",
          6901 => x"82",
          6902 => x"92",
          6903 => x"d7",
          6904 => x"98",
          6905 => x"73",
          6906 => x"38",
          6907 => x"9c",
          6908 => x"80",
          6909 => x"38",
          6910 => x"95",
          6911 => x"2e",
          6912 => x"aa",
          6913 => x"ea",
          6914 => x"b5",
          6915 => x"9e",
          6916 => x"05",
          6917 => x"54",
          6918 => x"38",
          6919 => x"70",
          6920 => x"54",
          6921 => x"8e",
          6922 => x"83",
          6923 => x"88",
          6924 => x"83",
          6925 => x"83",
          6926 => x"06",
          6927 => x"80",
          6928 => x"38",
          6929 => x"51",
          6930 => x"82",
          6931 => x"56",
          6932 => x"0a",
          6933 => x"05",
          6934 => x"3f",
          6935 => x"0b",
          6936 => x"80",
          6937 => x"7a",
          6938 => x"3f",
          6939 => x"9c",
          6940 => x"d1",
          6941 => x"81",
          6942 => x"34",
          6943 => x"80",
          6944 => x"b0",
          6945 => x"54",
          6946 => x"52",
          6947 => x"05",
          6948 => x"3f",
          6949 => x"08",
          6950 => x"a8",
          6951 => x"38",
          6952 => x"82",
          6953 => x"b2",
          6954 => x"84",
          6955 => x"06",
          6956 => x"73",
          6957 => x"38",
          6958 => x"ad",
          6959 => x"2a",
          6960 => x"51",
          6961 => x"2e",
          6962 => x"81",
          6963 => x"80",
          6964 => x"87",
          6965 => x"39",
          6966 => x"51",
          6967 => x"82",
          6968 => x"7b",
          6969 => x"12",
          6970 => x"82",
          6971 => x"81",
          6972 => x"83",
          6973 => x"06",
          6974 => x"80",
          6975 => x"77",
          6976 => x"58",
          6977 => x"08",
          6978 => x"63",
          6979 => x"63",
          6980 => x"57",
          6981 => x"82",
          6982 => x"82",
          6983 => x"88",
          6984 => x"9c",
          6985 => x"d2",
          6986 => x"b5",
          6987 => x"b5",
          6988 => x"1b",
          6989 => x"0c",
          6990 => x"22",
          6991 => x"77",
          6992 => x"80",
          6993 => x"34",
          6994 => x"1a",
          6995 => x"94",
          6996 => x"85",
          6997 => x"06",
          6998 => x"80",
          6999 => x"38",
          7000 => x"08",
          7001 => x"84",
          7002 => x"a8",
          7003 => x"0c",
          7004 => x"70",
          7005 => x"52",
          7006 => x"39",
          7007 => x"51",
          7008 => x"82",
          7009 => x"57",
          7010 => x"08",
          7011 => x"38",
          7012 => x"b5",
          7013 => x"2e",
          7014 => x"83",
          7015 => x"75",
          7016 => x"74",
          7017 => x"07",
          7018 => x"54",
          7019 => x"8a",
          7020 => x"75",
          7021 => x"73",
          7022 => x"98",
          7023 => x"a9",
          7024 => x"ff",
          7025 => x"80",
          7026 => x"76",
          7027 => x"d6",
          7028 => x"b5",
          7029 => x"38",
          7030 => x"39",
          7031 => x"82",
          7032 => x"05",
          7033 => x"84",
          7034 => x"0c",
          7035 => x"82",
          7036 => x"97",
          7037 => x"f2",
          7038 => x"63",
          7039 => x"40",
          7040 => x"7e",
          7041 => x"fc",
          7042 => x"51",
          7043 => x"82",
          7044 => x"55",
          7045 => x"08",
          7046 => x"19",
          7047 => x"80",
          7048 => x"74",
          7049 => x"39",
          7050 => x"81",
          7051 => x"56",
          7052 => x"82",
          7053 => x"39",
          7054 => x"1a",
          7055 => x"82",
          7056 => x"0b",
          7057 => x"81",
          7058 => x"39",
          7059 => x"94",
          7060 => x"55",
          7061 => x"83",
          7062 => x"7b",
          7063 => x"89",
          7064 => x"08",
          7065 => x"06",
          7066 => x"81",
          7067 => x"8a",
          7068 => x"05",
          7069 => x"06",
          7070 => x"a8",
          7071 => x"38",
          7072 => x"55",
          7073 => x"19",
          7074 => x"51",
          7075 => x"82",
          7076 => x"55",
          7077 => x"ff",
          7078 => x"ff",
          7079 => x"38",
          7080 => x"0c",
          7081 => x"52",
          7082 => x"cb",
          7083 => x"a8",
          7084 => x"ff",
          7085 => x"b5",
          7086 => x"7c",
          7087 => x"57",
          7088 => x"80",
          7089 => x"1a",
          7090 => x"22",
          7091 => x"75",
          7092 => x"38",
          7093 => x"58",
          7094 => x"53",
          7095 => x"1b",
          7096 => x"88",
          7097 => x"a8",
          7098 => x"38",
          7099 => x"33",
          7100 => x"80",
          7101 => x"b0",
          7102 => x"31",
          7103 => x"27",
          7104 => x"80",
          7105 => x"52",
          7106 => x"77",
          7107 => x"7d",
          7108 => x"e0",
          7109 => x"2b",
          7110 => x"76",
          7111 => x"94",
          7112 => x"ff",
          7113 => x"71",
          7114 => x"7b",
          7115 => x"38",
          7116 => x"19",
          7117 => x"51",
          7118 => x"82",
          7119 => x"fe",
          7120 => x"53",
          7121 => x"83",
          7122 => x"b4",
          7123 => x"51",
          7124 => x"7b",
          7125 => x"08",
          7126 => x"76",
          7127 => x"08",
          7128 => x"0c",
          7129 => x"f3",
          7130 => x"75",
          7131 => x"0c",
          7132 => x"04",
          7133 => x"60",
          7134 => x"40",
          7135 => x"80",
          7136 => x"3d",
          7137 => x"77",
          7138 => x"3f",
          7139 => x"08",
          7140 => x"a8",
          7141 => x"91",
          7142 => x"74",
          7143 => x"38",
          7144 => x"b8",
          7145 => x"33",
          7146 => x"70",
          7147 => x"56",
          7148 => x"74",
          7149 => x"a4",
          7150 => x"82",
          7151 => x"34",
          7152 => x"98",
          7153 => x"91",
          7154 => x"56",
          7155 => x"94",
          7156 => x"11",
          7157 => x"76",
          7158 => x"75",
          7159 => x"80",
          7160 => x"38",
          7161 => x"70",
          7162 => x"56",
          7163 => x"fd",
          7164 => x"11",
          7165 => x"77",
          7166 => x"5c",
          7167 => x"38",
          7168 => x"88",
          7169 => x"74",
          7170 => x"52",
          7171 => x"18",
          7172 => x"51",
          7173 => x"82",
          7174 => x"55",
          7175 => x"08",
          7176 => x"ab",
          7177 => x"2e",
          7178 => x"74",
          7179 => x"95",
          7180 => x"19",
          7181 => x"08",
          7182 => x"88",
          7183 => x"55",
          7184 => x"9c",
          7185 => x"09",
          7186 => x"38",
          7187 => x"c1",
          7188 => x"a8",
          7189 => x"38",
          7190 => x"52",
          7191 => x"97",
          7192 => x"a8",
          7193 => x"fe",
          7194 => x"b5",
          7195 => x"7c",
          7196 => x"57",
          7197 => x"80",
          7198 => x"1b",
          7199 => x"22",
          7200 => x"75",
          7201 => x"38",
          7202 => x"59",
          7203 => x"53",
          7204 => x"1a",
          7205 => x"be",
          7206 => x"a8",
          7207 => x"38",
          7208 => x"08",
          7209 => x"56",
          7210 => x"9b",
          7211 => x"53",
          7212 => x"77",
          7213 => x"7d",
          7214 => x"16",
          7215 => x"3f",
          7216 => x"0b",
          7217 => x"78",
          7218 => x"80",
          7219 => x"18",
          7220 => x"08",
          7221 => x"7e",
          7222 => x"3f",
          7223 => x"08",
          7224 => x"7e",
          7225 => x"0c",
          7226 => x"19",
          7227 => x"08",
          7228 => x"84",
          7229 => x"57",
          7230 => x"27",
          7231 => x"56",
          7232 => x"52",
          7233 => x"f9",
          7234 => x"a8",
          7235 => x"38",
          7236 => x"52",
          7237 => x"83",
          7238 => x"b4",
          7239 => x"d4",
          7240 => x"81",
          7241 => x"34",
          7242 => x"7e",
          7243 => x"0c",
          7244 => x"1a",
          7245 => x"94",
          7246 => x"1b",
          7247 => x"5e",
          7248 => x"27",
          7249 => x"55",
          7250 => x"0c",
          7251 => x"90",
          7252 => x"c0",
          7253 => x"90",
          7254 => x"56",
          7255 => x"a8",
          7256 => x"0d",
          7257 => x"0d",
          7258 => x"fc",
          7259 => x"52",
          7260 => x"3f",
          7261 => x"08",
          7262 => x"a8",
          7263 => x"38",
          7264 => x"70",
          7265 => x"81",
          7266 => x"55",
          7267 => x"80",
          7268 => x"16",
          7269 => x"51",
          7270 => x"82",
          7271 => x"57",
          7272 => x"08",
          7273 => x"a4",
          7274 => x"11",
          7275 => x"55",
          7276 => x"16",
          7277 => x"08",
          7278 => x"75",
          7279 => x"e8",
          7280 => x"08",
          7281 => x"51",
          7282 => x"82",
          7283 => x"52",
          7284 => x"c9",
          7285 => x"52",
          7286 => x"c9",
          7287 => x"54",
          7288 => x"15",
          7289 => x"cc",
          7290 => x"b5",
          7291 => x"17",
          7292 => x"06",
          7293 => x"90",
          7294 => x"82",
          7295 => x"8a",
          7296 => x"fc",
          7297 => x"70",
          7298 => x"d9",
          7299 => x"a8",
          7300 => x"b5",
          7301 => x"38",
          7302 => x"05",
          7303 => x"f1",
          7304 => x"b5",
          7305 => x"82",
          7306 => x"87",
          7307 => x"a8",
          7308 => x"72",
          7309 => x"0c",
          7310 => x"04",
          7311 => x"84",
          7312 => x"e4",
          7313 => x"80",
          7314 => x"a8",
          7315 => x"38",
          7316 => x"08",
          7317 => x"34",
          7318 => x"82",
          7319 => x"83",
          7320 => x"ef",
          7321 => x"53",
          7322 => x"05",
          7323 => x"51",
          7324 => x"82",
          7325 => x"55",
          7326 => x"08",
          7327 => x"76",
          7328 => x"93",
          7329 => x"51",
          7330 => x"82",
          7331 => x"55",
          7332 => x"08",
          7333 => x"80",
          7334 => x"70",
          7335 => x"56",
          7336 => x"89",
          7337 => x"94",
          7338 => x"b2",
          7339 => x"05",
          7340 => x"2a",
          7341 => x"51",
          7342 => x"80",
          7343 => x"76",
          7344 => x"52",
          7345 => x"3f",
          7346 => x"08",
          7347 => x"8e",
          7348 => x"a8",
          7349 => x"09",
          7350 => x"38",
          7351 => x"82",
          7352 => x"93",
          7353 => x"e4",
          7354 => x"6f",
          7355 => x"7a",
          7356 => x"9e",
          7357 => x"05",
          7358 => x"51",
          7359 => x"82",
          7360 => x"57",
          7361 => x"08",
          7362 => x"7b",
          7363 => x"94",
          7364 => x"55",
          7365 => x"73",
          7366 => x"ed",
          7367 => x"93",
          7368 => x"55",
          7369 => x"82",
          7370 => x"57",
          7371 => x"08",
          7372 => x"68",
          7373 => x"c9",
          7374 => x"b5",
          7375 => x"82",
          7376 => x"82",
          7377 => x"52",
          7378 => x"a3",
          7379 => x"a8",
          7380 => x"52",
          7381 => x"b8",
          7382 => x"a8",
          7383 => x"b5",
          7384 => x"a2",
          7385 => x"74",
          7386 => x"3f",
          7387 => x"08",
          7388 => x"a8",
          7389 => x"69",
          7390 => x"d9",
          7391 => x"82",
          7392 => x"2e",
          7393 => x"52",
          7394 => x"cf",
          7395 => x"a8",
          7396 => x"b5",
          7397 => x"2e",
          7398 => x"84",
          7399 => x"06",
          7400 => x"57",
          7401 => x"76",
          7402 => x"9e",
          7403 => x"05",
          7404 => x"dc",
          7405 => x"90",
          7406 => x"81",
          7407 => x"56",
          7408 => x"80",
          7409 => x"02",
          7410 => x"81",
          7411 => x"70",
          7412 => x"56",
          7413 => x"81",
          7414 => x"78",
          7415 => x"38",
          7416 => x"99",
          7417 => x"81",
          7418 => x"18",
          7419 => x"18",
          7420 => x"58",
          7421 => x"33",
          7422 => x"ee",
          7423 => x"6f",
          7424 => x"af",
          7425 => x"8d",
          7426 => x"2e",
          7427 => x"8a",
          7428 => x"6f",
          7429 => x"af",
          7430 => x"0b",
          7431 => x"33",
          7432 => x"82",
          7433 => x"70",
          7434 => x"52",
          7435 => x"56",
          7436 => x"8d",
          7437 => x"70",
          7438 => x"51",
          7439 => x"f5",
          7440 => x"54",
          7441 => x"a7",
          7442 => x"74",
          7443 => x"38",
          7444 => x"73",
          7445 => x"81",
          7446 => x"81",
          7447 => x"39",
          7448 => x"81",
          7449 => x"74",
          7450 => x"81",
          7451 => x"91",
          7452 => x"6e",
          7453 => x"59",
          7454 => x"7a",
          7455 => x"5c",
          7456 => x"26",
          7457 => x"7a",
          7458 => x"b5",
          7459 => x"3d",
          7460 => x"3d",
          7461 => x"8d",
          7462 => x"54",
          7463 => x"55",
          7464 => x"82",
          7465 => x"53",
          7466 => x"08",
          7467 => x"91",
          7468 => x"72",
          7469 => x"8c",
          7470 => x"73",
          7471 => x"38",
          7472 => x"70",
          7473 => x"81",
          7474 => x"57",
          7475 => x"73",
          7476 => x"08",
          7477 => x"94",
          7478 => x"75",
          7479 => x"97",
          7480 => x"11",
          7481 => x"2b",
          7482 => x"73",
          7483 => x"38",
          7484 => x"16",
          7485 => x"ac",
          7486 => x"a8",
          7487 => x"78",
          7488 => x"55",
          7489 => x"9c",
          7490 => x"a8",
          7491 => x"96",
          7492 => x"70",
          7493 => x"94",
          7494 => x"71",
          7495 => x"08",
          7496 => x"53",
          7497 => x"15",
          7498 => x"a6",
          7499 => x"74",
          7500 => x"3f",
          7501 => x"08",
          7502 => x"a8",
          7503 => x"81",
          7504 => x"b5",
          7505 => x"2e",
          7506 => x"82",
          7507 => x"88",
          7508 => x"98",
          7509 => x"80",
          7510 => x"38",
          7511 => x"80",
          7512 => x"77",
          7513 => x"08",
          7514 => x"0c",
          7515 => x"70",
          7516 => x"81",
          7517 => x"5a",
          7518 => x"2e",
          7519 => x"52",
          7520 => x"f9",
          7521 => x"a8",
          7522 => x"b5",
          7523 => x"38",
          7524 => x"08",
          7525 => x"73",
          7526 => x"c7",
          7527 => x"b5",
          7528 => x"73",
          7529 => x"38",
          7530 => x"af",
          7531 => x"73",
          7532 => x"27",
          7533 => x"98",
          7534 => x"a0",
          7535 => x"08",
          7536 => x"0c",
          7537 => x"06",
          7538 => x"2e",
          7539 => x"52",
          7540 => x"a3",
          7541 => x"a8",
          7542 => x"82",
          7543 => x"34",
          7544 => x"c4",
          7545 => x"91",
          7546 => x"53",
          7547 => x"89",
          7548 => x"a8",
          7549 => x"94",
          7550 => x"8c",
          7551 => x"27",
          7552 => x"8c",
          7553 => x"15",
          7554 => x"07",
          7555 => x"16",
          7556 => x"ff",
          7557 => x"80",
          7558 => x"77",
          7559 => x"2e",
          7560 => x"9c",
          7561 => x"53",
          7562 => x"a8",
          7563 => x"0d",
          7564 => x"0d",
          7565 => x"54",
          7566 => x"81",
          7567 => x"53",
          7568 => x"05",
          7569 => x"84",
          7570 => x"e7",
          7571 => x"a8",
          7572 => x"b5",
          7573 => x"ea",
          7574 => x"0c",
          7575 => x"51",
          7576 => x"82",
          7577 => x"55",
          7578 => x"08",
          7579 => x"ab",
          7580 => x"98",
          7581 => x"80",
          7582 => x"38",
          7583 => x"70",
          7584 => x"81",
          7585 => x"57",
          7586 => x"ad",
          7587 => x"08",
          7588 => x"d3",
          7589 => x"b5",
          7590 => x"17",
          7591 => x"86",
          7592 => x"17",
          7593 => x"75",
          7594 => x"3f",
          7595 => x"08",
          7596 => x"2e",
          7597 => x"85",
          7598 => x"86",
          7599 => x"2e",
          7600 => x"76",
          7601 => x"73",
          7602 => x"0c",
          7603 => x"04",
          7604 => x"76",
          7605 => x"05",
          7606 => x"53",
          7607 => x"82",
          7608 => x"87",
          7609 => x"a8",
          7610 => x"86",
          7611 => x"fb",
          7612 => x"79",
          7613 => x"05",
          7614 => x"56",
          7615 => x"3f",
          7616 => x"08",
          7617 => x"a8",
          7618 => x"38",
          7619 => x"82",
          7620 => x"52",
          7621 => x"f8",
          7622 => x"a8",
          7623 => x"ca",
          7624 => x"a8",
          7625 => x"51",
          7626 => x"82",
          7627 => x"53",
          7628 => x"08",
          7629 => x"81",
          7630 => x"80",
          7631 => x"82",
          7632 => x"a6",
          7633 => x"73",
          7634 => x"3f",
          7635 => x"51",
          7636 => x"82",
          7637 => x"84",
          7638 => x"70",
          7639 => x"2c",
          7640 => x"a8",
          7641 => x"51",
          7642 => x"82",
          7643 => x"87",
          7644 => x"ee",
          7645 => x"57",
          7646 => x"3d",
          7647 => x"3d",
          7648 => x"af",
          7649 => x"a8",
          7650 => x"b5",
          7651 => x"38",
          7652 => x"51",
          7653 => x"82",
          7654 => x"55",
          7655 => x"08",
          7656 => x"80",
          7657 => x"70",
          7658 => x"58",
          7659 => x"85",
          7660 => x"8d",
          7661 => x"2e",
          7662 => x"52",
          7663 => x"be",
          7664 => x"b5",
          7665 => x"3d",
          7666 => x"3d",
          7667 => x"55",
          7668 => x"92",
          7669 => x"52",
          7670 => x"de",
          7671 => x"b5",
          7672 => x"82",
          7673 => x"82",
          7674 => x"74",
          7675 => x"98",
          7676 => x"11",
          7677 => x"59",
          7678 => x"75",
          7679 => x"38",
          7680 => x"81",
          7681 => x"5b",
          7682 => x"82",
          7683 => x"39",
          7684 => x"08",
          7685 => x"59",
          7686 => x"09",
          7687 => x"38",
          7688 => x"57",
          7689 => x"3d",
          7690 => x"c1",
          7691 => x"b5",
          7692 => x"2e",
          7693 => x"b5",
          7694 => x"2e",
          7695 => x"b5",
          7696 => x"70",
          7697 => x"08",
          7698 => x"7a",
          7699 => x"7f",
          7700 => x"54",
          7701 => x"77",
          7702 => x"80",
          7703 => x"15",
          7704 => x"a8",
          7705 => x"75",
          7706 => x"52",
          7707 => x"52",
          7708 => x"8d",
          7709 => x"a8",
          7710 => x"b5",
          7711 => x"d6",
          7712 => x"33",
          7713 => x"1a",
          7714 => x"54",
          7715 => x"09",
          7716 => x"38",
          7717 => x"ff",
          7718 => x"82",
          7719 => x"83",
          7720 => x"70",
          7721 => x"25",
          7722 => x"59",
          7723 => x"9b",
          7724 => x"51",
          7725 => x"3f",
          7726 => x"08",
          7727 => x"70",
          7728 => x"25",
          7729 => x"59",
          7730 => x"75",
          7731 => x"7a",
          7732 => x"ff",
          7733 => x"7c",
          7734 => x"90",
          7735 => x"11",
          7736 => x"56",
          7737 => x"15",
          7738 => x"b5",
          7739 => x"3d",
          7740 => x"3d",
          7741 => x"3d",
          7742 => x"70",
          7743 => x"dd",
          7744 => x"a8",
          7745 => x"b5",
          7746 => x"a8",
          7747 => x"33",
          7748 => x"a0",
          7749 => x"33",
          7750 => x"70",
          7751 => x"55",
          7752 => x"73",
          7753 => x"8e",
          7754 => x"08",
          7755 => x"18",
          7756 => x"80",
          7757 => x"38",
          7758 => x"08",
          7759 => x"08",
          7760 => x"c4",
          7761 => x"b5",
          7762 => x"88",
          7763 => x"80",
          7764 => x"17",
          7765 => x"51",
          7766 => x"3f",
          7767 => x"08",
          7768 => x"81",
          7769 => x"81",
          7770 => x"a8",
          7771 => x"09",
          7772 => x"38",
          7773 => x"39",
          7774 => x"77",
          7775 => x"a8",
          7776 => x"08",
          7777 => x"98",
          7778 => x"82",
          7779 => x"52",
          7780 => x"bd",
          7781 => x"a8",
          7782 => x"17",
          7783 => x"0c",
          7784 => x"80",
          7785 => x"73",
          7786 => x"75",
          7787 => x"38",
          7788 => x"34",
          7789 => x"82",
          7790 => x"89",
          7791 => x"e2",
          7792 => x"53",
          7793 => x"a4",
          7794 => x"3d",
          7795 => x"3f",
          7796 => x"08",
          7797 => x"a8",
          7798 => x"38",
          7799 => x"3d",
          7800 => x"3d",
          7801 => x"d1",
          7802 => x"b5",
          7803 => x"82",
          7804 => x"81",
          7805 => x"80",
          7806 => x"70",
          7807 => x"81",
          7808 => x"56",
          7809 => x"81",
          7810 => x"98",
          7811 => x"74",
          7812 => x"38",
          7813 => x"05",
          7814 => x"06",
          7815 => x"55",
          7816 => x"38",
          7817 => x"51",
          7818 => x"82",
          7819 => x"74",
          7820 => x"81",
          7821 => x"56",
          7822 => x"80",
          7823 => x"54",
          7824 => x"08",
          7825 => x"2e",
          7826 => x"73",
          7827 => x"a8",
          7828 => x"52",
          7829 => x"52",
          7830 => x"3f",
          7831 => x"08",
          7832 => x"a8",
          7833 => x"38",
          7834 => x"08",
          7835 => x"cc",
          7836 => x"b5",
          7837 => x"82",
          7838 => x"86",
          7839 => x"80",
          7840 => x"b5",
          7841 => x"2e",
          7842 => x"b5",
          7843 => x"c0",
          7844 => x"ce",
          7845 => x"b5",
          7846 => x"b5",
          7847 => x"70",
          7848 => x"08",
          7849 => x"51",
          7850 => x"80",
          7851 => x"73",
          7852 => x"38",
          7853 => x"52",
          7854 => x"95",
          7855 => x"a8",
          7856 => x"8c",
          7857 => x"ff",
          7858 => x"82",
          7859 => x"55",
          7860 => x"a8",
          7861 => x"0d",
          7862 => x"0d",
          7863 => x"3d",
          7864 => x"9a",
          7865 => x"cb",
          7866 => x"a8",
          7867 => x"b5",
          7868 => x"b0",
          7869 => x"69",
          7870 => x"70",
          7871 => x"97",
          7872 => x"a8",
          7873 => x"b5",
          7874 => x"38",
          7875 => x"94",
          7876 => x"a8",
          7877 => x"09",
          7878 => x"88",
          7879 => x"df",
          7880 => x"85",
          7881 => x"51",
          7882 => x"74",
          7883 => x"78",
          7884 => x"8a",
          7885 => x"57",
          7886 => x"82",
          7887 => x"75",
          7888 => x"b5",
          7889 => x"38",
          7890 => x"b5",
          7891 => x"2e",
          7892 => x"83",
          7893 => x"82",
          7894 => x"ff",
          7895 => x"06",
          7896 => x"54",
          7897 => x"73",
          7898 => x"82",
          7899 => x"52",
          7900 => x"a4",
          7901 => x"a8",
          7902 => x"b5",
          7903 => x"9a",
          7904 => x"a0",
          7905 => x"51",
          7906 => x"3f",
          7907 => x"0b",
          7908 => x"78",
          7909 => x"bf",
          7910 => x"88",
          7911 => x"80",
          7912 => x"ff",
          7913 => x"75",
          7914 => x"11",
          7915 => x"f8",
          7916 => x"78",
          7917 => x"80",
          7918 => x"ff",
          7919 => x"78",
          7920 => x"80",
          7921 => x"7f",
          7922 => x"d4",
          7923 => x"c9",
          7924 => x"54",
          7925 => x"15",
          7926 => x"cb",
          7927 => x"b5",
          7928 => x"82",
          7929 => x"b2",
          7930 => x"b2",
          7931 => x"96",
          7932 => x"b5",
          7933 => x"53",
          7934 => x"51",
          7935 => x"64",
          7936 => x"8b",
          7937 => x"54",
          7938 => x"15",
          7939 => x"ff",
          7940 => x"82",
          7941 => x"54",
          7942 => x"53",
          7943 => x"51",
          7944 => x"3f",
          7945 => x"a8",
          7946 => x"0d",
          7947 => x"0d",
          7948 => x"05",
          7949 => x"3f",
          7950 => x"3d",
          7951 => x"52",
          7952 => x"d5",
          7953 => x"b5",
          7954 => x"82",
          7955 => x"82",
          7956 => x"4d",
          7957 => x"52",
          7958 => x"52",
          7959 => x"3f",
          7960 => x"08",
          7961 => x"a8",
          7962 => x"38",
          7963 => x"05",
          7964 => x"06",
          7965 => x"73",
          7966 => x"a0",
          7967 => x"08",
          7968 => x"ff",
          7969 => x"ff",
          7970 => x"ac",
          7971 => x"92",
          7972 => x"54",
          7973 => x"3f",
          7974 => x"52",
          7975 => x"f7",
          7976 => x"a8",
          7977 => x"b5",
          7978 => x"38",
          7979 => x"09",
          7980 => x"38",
          7981 => x"08",
          7982 => x"88",
          7983 => x"39",
          7984 => x"08",
          7985 => x"81",
          7986 => x"38",
          7987 => x"b1",
          7988 => x"a8",
          7989 => x"b5",
          7990 => x"c8",
          7991 => x"93",
          7992 => x"ff",
          7993 => x"8d",
          7994 => x"b4",
          7995 => x"af",
          7996 => x"17",
          7997 => x"33",
          7998 => x"70",
          7999 => x"55",
          8000 => x"38",
          8001 => x"54",
          8002 => x"34",
          8003 => x"0b",
          8004 => x"8b",
          8005 => x"84",
          8006 => x"06",
          8007 => x"73",
          8008 => x"e5",
          8009 => x"2e",
          8010 => x"75",
          8011 => x"c6",
          8012 => x"b5",
          8013 => x"78",
          8014 => x"bb",
          8015 => x"82",
          8016 => x"80",
          8017 => x"38",
          8018 => x"08",
          8019 => x"ff",
          8020 => x"82",
          8021 => x"79",
          8022 => x"58",
          8023 => x"b5",
          8024 => x"c0",
          8025 => x"33",
          8026 => x"2e",
          8027 => x"99",
          8028 => x"75",
          8029 => x"c6",
          8030 => x"54",
          8031 => x"15",
          8032 => x"82",
          8033 => x"9c",
          8034 => x"c8",
          8035 => x"b5",
          8036 => x"82",
          8037 => x"8c",
          8038 => x"ff",
          8039 => x"82",
          8040 => x"55",
          8041 => x"a8",
          8042 => x"0d",
          8043 => x"0d",
          8044 => x"05",
          8045 => x"05",
          8046 => x"33",
          8047 => x"53",
          8048 => x"05",
          8049 => x"51",
          8050 => x"82",
          8051 => x"55",
          8052 => x"08",
          8053 => x"78",
          8054 => x"95",
          8055 => x"51",
          8056 => x"82",
          8057 => x"55",
          8058 => x"08",
          8059 => x"80",
          8060 => x"81",
          8061 => x"86",
          8062 => x"38",
          8063 => x"61",
          8064 => x"12",
          8065 => x"7a",
          8066 => x"51",
          8067 => x"74",
          8068 => x"78",
          8069 => x"83",
          8070 => x"51",
          8071 => x"3f",
          8072 => x"08",
          8073 => x"b5",
          8074 => x"3d",
          8075 => x"3d",
          8076 => x"82",
          8077 => x"d0",
          8078 => x"3d",
          8079 => x"3f",
          8080 => x"08",
          8081 => x"a8",
          8082 => x"38",
          8083 => x"52",
          8084 => x"05",
          8085 => x"3f",
          8086 => x"08",
          8087 => x"a8",
          8088 => x"02",
          8089 => x"33",
          8090 => x"54",
          8091 => x"a6",
          8092 => x"22",
          8093 => x"71",
          8094 => x"53",
          8095 => x"51",
          8096 => x"3f",
          8097 => x"0b",
          8098 => x"76",
          8099 => x"b8",
          8100 => x"a8",
          8101 => x"82",
          8102 => x"93",
          8103 => x"ea",
          8104 => x"6b",
          8105 => x"53",
          8106 => x"05",
          8107 => x"51",
          8108 => x"82",
          8109 => x"82",
          8110 => x"30",
          8111 => x"a8",
          8112 => x"25",
          8113 => x"79",
          8114 => x"85",
          8115 => x"75",
          8116 => x"73",
          8117 => x"f9",
          8118 => x"80",
          8119 => x"8d",
          8120 => x"54",
          8121 => x"3f",
          8122 => x"08",
          8123 => x"a8",
          8124 => x"38",
          8125 => x"51",
          8126 => x"82",
          8127 => x"57",
          8128 => x"08",
          8129 => x"b5",
          8130 => x"b5",
          8131 => x"5b",
          8132 => x"18",
          8133 => x"18",
          8134 => x"74",
          8135 => x"81",
          8136 => x"78",
          8137 => x"8b",
          8138 => x"54",
          8139 => x"75",
          8140 => x"38",
          8141 => x"1b",
          8142 => x"55",
          8143 => x"2e",
          8144 => x"39",
          8145 => x"09",
          8146 => x"38",
          8147 => x"80",
          8148 => x"70",
          8149 => x"25",
          8150 => x"80",
          8151 => x"38",
          8152 => x"bc",
          8153 => x"11",
          8154 => x"ff",
          8155 => x"82",
          8156 => x"57",
          8157 => x"08",
          8158 => x"70",
          8159 => x"80",
          8160 => x"83",
          8161 => x"80",
          8162 => x"84",
          8163 => x"a7",
          8164 => x"b4",
          8165 => x"ad",
          8166 => x"b5",
          8167 => x"0c",
          8168 => x"a8",
          8169 => x"0d",
          8170 => x"0d",
          8171 => x"3d",
          8172 => x"52",
          8173 => x"ce",
          8174 => x"b5",
          8175 => x"b5",
          8176 => x"54",
          8177 => x"08",
          8178 => x"8b",
          8179 => x"8b",
          8180 => x"59",
          8181 => x"3f",
          8182 => x"33",
          8183 => x"06",
          8184 => x"57",
          8185 => x"81",
          8186 => x"58",
          8187 => x"06",
          8188 => x"4e",
          8189 => x"ff",
          8190 => x"82",
          8191 => x"80",
          8192 => x"6c",
          8193 => x"53",
          8194 => x"ae",
          8195 => x"b5",
          8196 => x"2e",
          8197 => x"88",
          8198 => x"6d",
          8199 => x"55",
          8200 => x"b5",
          8201 => x"ff",
          8202 => x"83",
          8203 => x"51",
          8204 => x"26",
          8205 => x"15",
          8206 => x"ff",
          8207 => x"80",
          8208 => x"87",
          8209 => x"f0",
          8210 => x"74",
          8211 => x"38",
          8212 => x"af",
          8213 => x"ae",
          8214 => x"b5",
          8215 => x"38",
          8216 => x"27",
          8217 => x"89",
          8218 => x"8b",
          8219 => x"27",
          8220 => x"55",
          8221 => x"81",
          8222 => x"8f",
          8223 => x"2a",
          8224 => x"70",
          8225 => x"34",
          8226 => x"74",
          8227 => x"05",
          8228 => x"17",
          8229 => x"70",
          8230 => x"52",
          8231 => x"73",
          8232 => x"c8",
          8233 => x"33",
          8234 => x"73",
          8235 => x"81",
          8236 => x"80",
          8237 => x"02",
          8238 => x"76",
          8239 => x"51",
          8240 => x"2e",
          8241 => x"87",
          8242 => x"57",
          8243 => x"79",
          8244 => x"80",
          8245 => x"70",
          8246 => x"ba",
          8247 => x"b5",
          8248 => x"82",
          8249 => x"80",
          8250 => x"52",
          8251 => x"bf",
          8252 => x"b5",
          8253 => x"82",
          8254 => x"8d",
          8255 => x"c4",
          8256 => x"e5",
          8257 => x"c6",
          8258 => x"a8",
          8259 => x"09",
          8260 => x"cc",
          8261 => x"76",
          8262 => x"c4",
          8263 => x"74",
          8264 => x"b0",
          8265 => x"a8",
          8266 => x"b5",
          8267 => x"38",
          8268 => x"b5",
          8269 => x"67",
          8270 => x"db",
          8271 => x"88",
          8272 => x"34",
          8273 => x"52",
          8274 => x"ab",
          8275 => x"54",
          8276 => x"15",
          8277 => x"ff",
          8278 => x"82",
          8279 => x"54",
          8280 => x"82",
          8281 => x"9c",
          8282 => x"f2",
          8283 => x"62",
          8284 => x"80",
          8285 => x"93",
          8286 => x"55",
          8287 => x"5e",
          8288 => x"3f",
          8289 => x"08",
          8290 => x"a8",
          8291 => x"38",
          8292 => x"58",
          8293 => x"38",
          8294 => x"97",
          8295 => x"08",
          8296 => x"38",
          8297 => x"70",
          8298 => x"81",
          8299 => x"55",
          8300 => x"87",
          8301 => x"39",
          8302 => x"90",
          8303 => x"82",
          8304 => x"8a",
          8305 => x"89",
          8306 => x"7f",
          8307 => x"56",
          8308 => x"3f",
          8309 => x"06",
          8310 => x"72",
          8311 => x"82",
          8312 => x"05",
          8313 => x"7c",
          8314 => x"55",
          8315 => x"27",
          8316 => x"16",
          8317 => x"83",
          8318 => x"76",
          8319 => x"80",
          8320 => x"79",
          8321 => x"99",
          8322 => x"7f",
          8323 => x"14",
          8324 => x"83",
          8325 => x"82",
          8326 => x"81",
          8327 => x"38",
          8328 => x"08",
          8329 => x"95",
          8330 => x"a8",
          8331 => x"81",
          8332 => x"7b",
          8333 => x"06",
          8334 => x"39",
          8335 => x"56",
          8336 => x"09",
          8337 => x"b9",
          8338 => x"80",
          8339 => x"80",
          8340 => x"78",
          8341 => x"7a",
          8342 => x"38",
          8343 => x"73",
          8344 => x"81",
          8345 => x"ff",
          8346 => x"74",
          8347 => x"ff",
          8348 => x"82",
          8349 => x"58",
          8350 => x"08",
          8351 => x"74",
          8352 => x"16",
          8353 => x"73",
          8354 => x"39",
          8355 => x"7e",
          8356 => x"0c",
          8357 => x"2e",
          8358 => x"88",
          8359 => x"8c",
          8360 => x"1a",
          8361 => x"07",
          8362 => x"1b",
          8363 => x"08",
          8364 => x"16",
          8365 => x"75",
          8366 => x"38",
          8367 => x"90",
          8368 => x"15",
          8369 => x"54",
          8370 => x"34",
          8371 => x"82",
          8372 => x"90",
          8373 => x"e9",
          8374 => x"6d",
          8375 => x"80",
          8376 => x"9d",
          8377 => x"5c",
          8378 => x"3f",
          8379 => x"0b",
          8380 => x"08",
          8381 => x"38",
          8382 => x"08",
          8383 => x"cc",
          8384 => x"08",
          8385 => x"80",
          8386 => x"80",
          8387 => x"b5",
          8388 => x"ff",
          8389 => x"52",
          8390 => x"a0",
          8391 => x"b5",
          8392 => x"ff",
          8393 => x"06",
          8394 => x"56",
          8395 => x"38",
          8396 => x"70",
          8397 => x"55",
          8398 => x"8b",
          8399 => x"3d",
          8400 => x"83",
          8401 => x"ff",
          8402 => x"82",
          8403 => x"99",
          8404 => x"74",
          8405 => x"38",
          8406 => x"80",
          8407 => x"ff",
          8408 => x"55",
          8409 => x"83",
          8410 => x"78",
          8411 => x"38",
          8412 => x"26",
          8413 => x"81",
          8414 => x"8b",
          8415 => x"79",
          8416 => x"80",
          8417 => x"93",
          8418 => x"39",
          8419 => x"6e",
          8420 => x"89",
          8421 => x"48",
          8422 => x"83",
          8423 => x"61",
          8424 => x"25",
          8425 => x"55",
          8426 => x"8a",
          8427 => x"3d",
          8428 => x"81",
          8429 => x"ff",
          8430 => x"81",
          8431 => x"a8",
          8432 => x"38",
          8433 => x"70",
          8434 => x"b5",
          8435 => x"56",
          8436 => x"38",
          8437 => x"55",
          8438 => x"75",
          8439 => x"38",
          8440 => x"70",
          8441 => x"ff",
          8442 => x"83",
          8443 => x"78",
          8444 => x"89",
          8445 => x"81",
          8446 => x"06",
          8447 => x"80",
          8448 => x"77",
          8449 => x"74",
          8450 => x"8d",
          8451 => x"06",
          8452 => x"2e",
          8453 => x"77",
          8454 => x"93",
          8455 => x"74",
          8456 => x"cb",
          8457 => x"7d",
          8458 => x"81",
          8459 => x"38",
          8460 => x"66",
          8461 => x"81",
          8462 => x"94",
          8463 => x"74",
          8464 => x"38",
          8465 => x"98",
          8466 => x"94",
          8467 => x"82",
          8468 => x"57",
          8469 => x"80",
          8470 => x"76",
          8471 => x"38",
          8472 => x"51",
          8473 => x"3f",
          8474 => x"08",
          8475 => x"87",
          8476 => x"2a",
          8477 => x"5c",
          8478 => x"b5",
          8479 => x"80",
          8480 => x"44",
          8481 => x"0a",
          8482 => x"ec",
          8483 => x"39",
          8484 => x"66",
          8485 => x"81",
          8486 => x"84",
          8487 => x"74",
          8488 => x"38",
          8489 => x"98",
          8490 => x"84",
          8491 => x"82",
          8492 => x"57",
          8493 => x"80",
          8494 => x"76",
          8495 => x"38",
          8496 => x"51",
          8497 => x"3f",
          8498 => x"08",
          8499 => x"57",
          8500 => x"08",
          8501 => x"96",
          8502 => x"82",
          8503 => x"10",
          8504 => x"08",
          8505 => x"72",
          8506 => x"59",
          8507 => x"ff",
          8508 => x"5d",
          8509 => x"44",
          8510 => x"11",
          8511 => x"70",
          8512 => x"71",
          8513 => x"06",
          8514 => x"52",
          8515 => x"40",
          8516 => x"09",
          8517 => x"38",
          8518 => x"18",
          8519 => x"39",
          8520 => x"79",
          8521 => x"70",
          8522 => x"58",
          8523 => x"76",
          8524 => x"38",
          8525 => x"7d",
          8526 => x"70",
          8527 => x"55",
          8528 => x"3f",
          8529 => x"08",
          8530 => x"2e",
          8531 => x"9b",
          8532 => x"a8",
          8533 => x"f5",
          8534 => x"38",
          8535 => x"38",
          8536 => x"59",
          8537 => x"38",
          8538 => x"7d",
          8539 => x"81",
          8540 => x"38",
          8541 => x"0b",
          8542 => x"08",
          8543 => x"78",
          8544 => x"1a",
          8545 => x"c0",
          8546 => x"74",
          8547 => x"39",
          8548 => x"55",
          8549 => x"8f",
          8550 => x"fd",
          8551 => x"b5",
          8552 => x"f5",
          8553 => x"78",
          8554 => x"79",
          8555 => x"80",
          8556 => x"f1",
          8557 => x"39",
          8558 => x"81",
          8559 => x"06",
          8560 => x"55",
          8561 => x"27",
          8562 => x"81",
          8563 => x"56",
          8564 => x"38",
          8565 => x"80",
          8566 => x"ff",
          8567 => x"8b",
          8568 => x"ac",
          8569 => x"ff",
          8570 => x"84",
          8571 => x"1b",
          8572 => x"b3",
          8573 => x"1c",
          8574 => x"ff",
          8575 => x"8e",
          8576 => x"a1",
          8577 => x"0b",
          8578 => x"7d",
          8579 => x"30",
          8580 => x"84",
          8581 => x"51",
          8582 => x"51",
          8583 => x"3f",
          8584 => x"83",
          8585 => x"90",
          8586 => x"ff",
          8587 => x"93",
          8588 => x"a0",
          8589 => x"39",
          8590 => x"1b",
          8591 => x"85",
          8592 => x"95",
          8593 => x"52",
          8594 => x"ff",
          8595 => x"81",
          8596 => x"1b",
          8597 => x"cf",
          8598 => x"9c",
          8599 => x"a0",
          8600 => x"83",
          8601 => x"06",
          8602 => x"82",
          8603 => x"52",
          8604 => x"51",
          8605 => x"3f",
          8606 => x"1b",
          8607 => x"c5",
          8608 => x"ac",
          8609 => x"a0",
          8610 => x"52",
          8611 => x"ff",
          8612 => x"86",
          8613 => x"51",
          8614 => x"3f",
          8615 => x"80",
          8616 => x"a9",
          8617 => x"1c",
          8618 => x"82",
          8619 => x"80",
          8620 => x"ae",
          8621 => x"b2",
          8622 => x"1b",
          8623 => x"85",
          8624 => x"ff",
          8625 => x"96",
          8626 => x"9f",
          8627 => x"80",
          8628 => x"34",
          8629 => x"1c",
          8630 => x"82",
          8631 => x"ab",
          8632 => x"a0",
          8633 => x"d4",
          8634 => x"fe",
          8635 => x"59",
          8636 => x"3f",
          8637 => x"53",
          8638 => x"51",
          8639 => x"3f",
          8640 => x"b5",
          8641 => x"e7",
          8642 => x"2e",
          8643 => x"80",
          8644 => x"54",
          8645 => x"53",
          8646 => x"51",
          8647 => x"3f",
          8648 => x"80",
          8649 => x"ff",
          8650 => x"84",
          8651 => x"d2",
          8652 => x"ff",
          8653 => x"86",
          8654 => x"f2",
          8655 => x"1b",
          8656 => x"81",
          8657 => x"52",
          8658 => x"51",
          8659 => x"3f",
          8660 => x"ec",
          8661 => x"9e",
          8662 => x"d4",
          8663 => x"51",
          8664 => x"3f",
          8665 => x"87",
          8666 => x"52",
          8667 => x"9a",
          8668 => x"54",
          8669 => x"7a",
          8670 => x"ff",
          8671 => x"65",
          8672 => x"7a",
          8673 => x"8f",
          8674 => x"80",
          8675 => x"2e",
          8676 => x"9a",
          8677 => x"7a",
          8678 => x"a9",
          8679 => x"84",
          8680 => x"9e",
          8681 => x"0a",
          8682 => x"51",
          8683 => x"ff",
          8684 => x"7d",
          8685 => x"38",
          8686 => x"52",
          8687 => x"9e",
          8688 => x"55",
          8689 => x"62",
          8690 => x"74",
          8691 => x"75",
          8692 => x"7e",
          8693 => x"fe",
          8694 => x"a8",
          8695 => x"38",
          8696 => x"82",
          8697 => x"52",
          8698 => x"9e",
          8699 => x"16",
          8700 => x"56",
          8701 => x"38",
          8702 => x"77",
          8703 => x"8d",
          8704 => x"7d",
          8705 => x"38",
          8706 => x"57",
          8707 => x"83",
          8708 => x"76",
          8709 => x"7a",
          8710 => x"ff",
          8711 => x"82",
          8712 => x"81",
          8713 => x"16",
          8714 => x"56",
          8715 => x"38",
          8716 => x"83",
          8717 => x"86",
          8718 => x"ff",
          8719 => x"38",
          8720 => x"82",
          8721 => x"81",
          8722 => x"06",
          8723 => x"fe",
          8724 => x"53",
          8725 => x"51",
          8726 => x"3f",
          8727 => x"52",
          8728 => x"9c",
          8729 => x"be",
          8730 => x"75",
          8731 => x"81",
          8732 => x"0b",
          8733 => x"77",
          8734 => x"75",
          8735 => x"60",
          8736 => x"80",
          8737 => x"75",
          8738 => x"98",
          8739 => x"85",
          8740 => x"b5",
          8741 => x"2a",
          8742 => x"75",
          8743 => x"82",
          8744 => x"87",
          8745 => x"52",
          8746 => x"51",
          8747 => x"3f",
          8748 => x"ca",
          8749 => x"9c",
          8750 => x"54",
          8751 => x"52",
          8752 => x"98",
          8753 => x"56",
          8754 => x"08",
          8755 => x"53",
          8756 => x"51",
          8757 => x"3f",
          8758 => x"b5",
          8759 => x"38",
          8760 => x"56",
          8761 => x"56",
          8762 => x"b5",
          8763 => x"75",
          8764 => x"0c",
          8765 => x"04",
          8766 => x"7d",
          8767 => x"80",
          8768 => x"05",
          8769 => x"76",
          8770 => x"38",
          8771 => x"11",
          8772 => x"53",
          8773 => x"79",
          8774 => x"3f",
          8775 => x"09",
          8776 => x"38",
          8777 => x"55",
          8778 => x"db",
          8779 => x"70",
          8780 => x"34",
          8781 => x"74",
          8782 => x"81",
          8783 => x"80",
          8784 => x"55",
          8785 => x"76",
          8786 => x"b5",
          8787 => x"3d",
          8788 => x"3d",
          8789 => x"84",
          8790 => x"33",
          8791 => x"8a",
          8792 => x"06",
          8793 => x"52",
          8794 => x"3f",
          8795 => x"56",
          8796 => x"be",
          8797 => x"08",
          8798 => x"05",
          8799 => x"75",
          8800 => x"56",
          8801 => x"a1",
          8802 => x"fc",
          8803 => x"53",
          8804 => x"76",
          8805 => x"dc",
          8806 => x"32",
          8807 => x"72",
          8808 => x"70",
          8809 => x"56",
          8810 => x"18",
          8811 => x"88",
          8812 => x"3d",
          8813 => x"3d",
          8814 => x"11",
          8815 => x"80",
          8816 => x"38",
          8817 => x"05",
          8818 => x"8c",
          8819 => x"08",
          8820 => x"3f",
          8821 => x"08",
          8822 => x"16",
          8823 => x"09",
          8824 => x"38",
          8825 => x"55",
          8826 => x"55",
          8827 => x"a8",
          8828 => x"0d",
          8829 => x"0d",
          8830 => x"cc",
          8831 => x"73",
          8832 => x"93",
          8833 => x"0c",
          8834 => x"04",
          8835 => x"02",
          8836 => x"33",
          8837 => x"3d",
          8838 => x"54",
          8839 => x"52",
          8840 => x"ae",
          8841 => x"ff",
          8842 => x"3d",
          8843 => x"00",
          8844 => x"ff",
          8845 => x"ff",
          8846 => x"00",
          8847 => x"ff",
          8848 => x"2b",
          8849 => x"2b",
          8850 => x"2b",
          8851 => x"2b",
          8852 => x"2b",
          8853 => x"2b",
          8854 => x"2b",
          8855 => x"2b",
          8856 => x"2b",
          8857 => x"2b",
          8858 => x"2b",
          8859 => x"2b",
          8860 => x"2b",
          8861 => x"2b",
          8862 => x"2b",
          8863 => x"2b",
          8864 => x"2b",
          8865 => x"2b",
          8866 => x"2b",
          8867 => x"2b",
          8868 => x"41",
          8869 => x"41",
          8870 => x"41",
          8871 => x"41",
          8872 => x"41",
          8873 => x"47",
          8874 => x"48",
          8875 => x"49",
          8876 => x"4b",
          8877 => x"47",
          8878 => x"45",
          8879 => x"49",
          8880 => x"4b",
          8881 => x"4a",
          8882 => x"4a",
          8883 => x"4a",
          8884 => x"48",
          8885 => x"45",
          8886 => x"49",
          8887 => x"49",
          8888 => x"49",
          8889 => x"45",
          8890 => x"45",
          8891 => x"4a",
          8892 => x"4a",
          8893 => x"4b",
          8894 => x"4b",
          8895 => x"0e",
          8896 => x"17",
          8897 => x"17",
          8898 => x"0e",
          8899 => x"17",
          8900 => x"17",
          8901 => x"17",
          8902 => x"17",
          8903 => x"17",
          8904 => x"17",
          8905 => x"17",
          8906 => x"0e",
          8907 => x"17",
          8908 => x"0e",
          8909 => x"0e",
          8910 => x"17",
          8911 => x"17",
          8912 => x"17",
          8913 => x"17",
          8914 => x"17",
          8915 => x"17",
          8916 => x"17",
          8917 => x"17",
          8918 => x"17",
          8919 => x"17",
          8920 => x"17",
          8921 => x"17",
          8922 => x"17",
          8923 => x"17",
          8924 => x"17",
          8925 => x"17",
          8926 => x"17",
          8927 => x"17",
          8928 => x"17",
          8929 => x"17",
          8930 => x"17",
          8931 => x"17",
          8932 => x"17",
          8933 => x"17",
          8934 => x"17",
          8935 => x"17",
          8936 => x"17",
          8937 => x"17",
          8938 => x"17",
          8939 => x"17",
          8940 => x"17",
          8941 => x"17",
          8942 => x"17",
          8943 => x"17",
          8944 => x"17",
          8945 => x"17",
          8946 => x"0f",
          8947 => x"17",
          8948 => x"17",
          8949 => x"17",
          8950 => x"17",
          8951 => x"11",
          8952 => x"17",
          8953 => x"17",
          8954 => x"17",
          8955 => x"17",
          8956 => x"17",
          8957 => x"17",
          8958 => x"17",
          8959 => x"17",
          8960 => x"17",
          8961 => x"17",
          8962 => x"0e",
          8963 => x"10",
          8964 => x"0e",
          8965 => x"0e",
          8966 => x"0e",
          8967 => x"17",
          8968 => x"10",
          8969 => x"17",
          8970 => x"17",
          8971 => x"0e",
          8972 => x"17",
          8973 => x"17",
          8974 => x"10",
          8975 => x"10",
          8976 => x"17",
          8977 => x"17",
          8978 => x"0f",
          8979 => x"17",
          8980 => x"11",
          8981 => x"17",
          8982 => x"17",
          8983 => x"11",
          8984 => x"6e",
          8985 => x"00",
          8986 => x"6f",
          8987 => x"00",
          8988 => x"6e",
          8989 => x"00",
          8990 => x"6f",
          8991 => x"00",
          8992 => x"78",
          8993 => x"00",
          8994 => x"6c",
          8995 => x"00",
          8996 => x"6f",
          8997 => x"00",
          8998 => x"69",
          8999 => x"00",
          9000 => x"75",
          9001 => x"00",
          9002 => x"62",
          9003 => x"68",
          9004 => x"77",
          9005 => x"64",
          9006 => x"65",
          9007 => x"64",
          9008 => x"65",
          9009 => x"6c",
          9010 => x"00",
          9011 => x"70",
          9012 => x"73",
          9013 => x"74",
          9014 => x"73",
          9015 => x"00",
          9016 => x"66",
          9017 => x"00",
          9018 => x"73",
          9019 => x"00",
          9020 => x"61",
          9021 => x"00",
          9022 => x"61",
          9023 => x"00",
          9024 => x"6c",
          9025 => x"00",
          9026 => x"00",
          9027 => x"73",
          9028 => x"72",
          9029 => x"0a",
          9030 => x"74",
          9031 => x"61",
          9032 => x"72",
          9033 => x"2e",
          9034 => x"00",
          9035 => x"73",
          9036 => x"6f",
          9037 => x"65",
          9038 => x"2e",
          9039 => x"00",
          9040 => x"20",
          9041 => x"65",
          9042 => x"75",
          9043 => x"0a",
          9044 => x"20",
          9045 => x"68",
          9046 => x"75",
          9047 => x"0a",
          9048 => x"76",
          9049 => x"64",
          9050 => x"6c",
          9051 => x"6d",
          9052 => x"00",
          9053 => x"63",
          9054 => x"20",
          9055 => x"69",
          9056 => x"0a",
          9057 => x"6c",
          9058 => x"6c",
          9059 => x"64",
          9060 => x"78",
          9061 => x"73",
          9062 => x"00",
          9063 => x"6c",
          9064 => x"61",
          9065 => x"65",
          9066 => x"76",
          9067 => x"64",
          9068 => x"00",
          9069 => x"20",
          9070 => x"77",
          9071 => x"65",
          9072 => x"6f",
          9073 => x"74",
          9074 => x"0a",
          9075 => x"69",
          9076 => x"6e",
          9077 => x"65",
          9078 => x"73",
          9079 => x"76",
          9080 => x"64",
          9081 => x"00",
          9082 => x"73",
          9083 => x"6f",
          9084 => x"6e",
          9085 => x"65",
          9086 => x"00",
          9087 => x"20",
          9088 => x"70",
          9089 => x"62",
          9090 => x"66",
          9091 => x"73",
          9092 => x"65",
          9093 => x"6f",
          9094 => x"20",
          9095 => x"64",
          9096 => x"2e",
          9097 => x"00",
          9098 => x"72",
          9099 => x"20",
          9100 => x"72",
          9101 => x"2e",
          9102 => x"00",
          9103 => x"6d",
          9104 => x"74",
          9105 => x"70",
          9106 => x"74",
          9107 => x"20",
          9108 => x"63",
          9109 => x"65",
          9110 => x"00",
          9111 => x"6c",
          9112 => x"73",
          9113 => x"63",
          9114 => x"2e",
          9115 => x"00",
          9116 => x"73",
          9117 => x"69",
          9118 => x"6e",
          9119 => x"65",
          9120 => x"79",
          9121 => x"00",
          9122 => x"6f",
          9123 => x"6e",
          9124 => x"70",
          9125 => x"66",
          9126 => x"73",
          9127 => x"00",
          9128 => x"72",
          9129 => x"74",
          9130 => x"20",
          9131 => x"6f",
          9132 => x"63",
          9133 => x"00",
          9134 => x"63",
          9135 => x"73",
          9136 => x"00",
          9137 => x"6b",
          9138 => x"6e",
          9139 => x"72",
          9140 => x"0a",
          9141 => x"6c",
          9142 => x"79",
          9143 => x"20",
          9144 => x"61",
          9145 => x"6c",
          9146 => x"79",
          9147 => x"2f",
          9148 => x"2e",
          9149 => x"00",
          9150 => x"61",
          9151 => x"00",
          9152 => x"38",
          9153 => x"00",
          9154 => x"20",
          9155 => x"34",
          9156 => x"00",
          9157 => x"20",
          9158 => x"20",
          9159 => x"00",
          9160 => x"32",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"0a",
          9165 => x"53",
          9166 => x"2a",
          9167 => x"20",
          9168 => x"00",
          9169 => x"2f",
          9170 => x"32",
          9171 => x"00",
          9172 => x"2e",
          9173 => x"00",
          9174 => x"50",
          9175 => x"72",
          9176 => x"25",
          9177 => x"29",
          9178 => x"20",
          9179 => x"2a",
          9180 => x"00",
          9181 => x"55",
          9182 => x"74",
          9183 => x"75",
          9184 => x"48",
          9185 => x"6c",
          9186 => x"00",
          9187 => x"6d",
          9188 => x"69",
          9189 => x"72",
          9190 => x"74",
          9191 => x"00",
          9192 => x"32",
          9193 => x"74",
          9194 => x"75",
          9195 => x"00",
          9196 => x"43",
          9197 => x"52",
          9198 => x"6e",
          9199 => x"72",
          9200 => x"0a",
          9201 => x"43",
          9202 => x"57",
          9203 => x"6e",
          9204 => x"72",
          9205 => x"0a",
          9206 => x"52",
          9207 => x"52",
          9208 => x"6e",
          9209 => x"72",
          9210 => x"0a",
          9211 => x"52",
          9212 => x"54",
          9213 => x"6e",
          9214 => x"72",
          9215 => x"0a",
          9216 => x"52",
          9217 => x"52",
          9218 => x"6e",
          9219 => x"72",
          9220 => x"0a",
          9221 => x"52",
          9222 => x"54",
          9223 => x"6e",
          9224 => x"72",
          9225 => x"0a",
          9226 => x"74",
          9227 => x"67",
          9228 => x"20",
          9229 => x"65",
          9230 => x"2e",
          9231 => x"00",
          9232 => x"61",
          9233 => x"6e",
          9234 => x"69",
          9235 => x"2e",
          9236 => x"00",
          9237 => x"74",
          9238 => x"65",
          9239 => x"61",
          9240 => x"00",
          9241 => x"53",
          9242 => x"74",
          9243 => x"00",
          9244 => x"69",
          9245 => x"20",
          9246 => x"69",
          9247 => x"69",
          9248 => x"73",
          9249 => x"64",
          9250 => x"72",
          9251 => x"2c",
          9252 => x"65",
          9253 => x"20",
          9254 => x"74",
          9255 => x"6e",
          9256 => x"6c",
          9257 => x"00",
          9258 => x"00",
          9259 => x"65",
          9260 => x"6e",
          9261 => x"2e",
          9262 => x"00",
          9263 => x"70",
          9264 => x"67",
          9265 => x"00",
          9266 => x"6d",
          9267 => x"69",
          9268 => x"2e",
          9269 => x"00",
          9270 => x"38",
          9271 => x"25",
          9272 => x"29",
          9273 => x"30",
          9274 => x"28",
          9275 => x"78",
          9276 => x"00",
          9277 => x"6d",
          9278 => x"65",
          9279 => x"79",
          9280 => x"00",
          9281 => x"6f",
          9282 => x"65",
          9283 => x"0a",
          9284 => x"38",
          9285 => x"30",
          9286 => x"00",
          9287 => x"3f",
          9288 => x"00",
          9289 => x"38",
          9290 => x"30",
          9291 => x"00",
          9292 => x"38",
          9293 => x"30",
          9294 => x"00",
          9295 => x"65",
          9296 => x"69",
          9297 => x"63",
          9298 => x"20",
          9299 => x"30",
          9300 => x"2e",
          9301 => x"00",
          9302 => x"6c",
          9303 => x"67",
          9304 => x"64",
          9305 => x"20",
          9306 => x"78",
          9307 => x"2e",
          9308 => x"00",
          9309 => x"6c",
          9310 => x"65",
          9311 => x"6e",
          9312 => x"63",
          9313 => x"20",
          9314 => x"29",
          9315 => x"00",
          9316 => x"73",
          9317 => x"74",
          9318 => x"20",
          9319 => x"6c",
          9320 => x"74",
          9321 => x"2e",
          9322 => x"00",
          9323 => x"6c",
          9324 => x"65",
          9325 => x"74",
          9326 => x"2e",
          9327 => x"00",
          9328 => x"55",
          9329 => x"6e",
          9330 => x"3a",
          9331 => x"5c",
          9332 => x"25",
          9333 => x"00",
          9334 => x"3a",
          9335 => x"5c",
          9336 => x"00",
          9337 => x"3a",
          9338 => x"00",
          9339 => x"64",
          9340 => x"6d",
          9341 => x"64",
          9342 => x"00",
          9343 => x"4c",
          9344 => x"31",
          9345 => x"4f",
          9346 => x"52",
          9347 => x"46",
          9348 => x"4c",
          9349 => x"32",
          9350 => x"4f",
          9351 => x"52",
          9352 => x"46",
          9353 => x"6e",
          9354 => x"67",
          9355 => x"0a",
          9356 => x"61",
          9357 => x"6e",
          9358 => x"6e",
          9359 => x"72",
          9360 => x"73",
          9361 => x"0a",
          9362 => x"2f",
          9363 => x"25",
          9364 => x"64",
          9365 => x"3a",
          9366 => x"25",
          9367 => x"0a",
          9368 => x"43",
          9369 => x"6e",
          9370 => x"75",
          9371 => x"69",
          9372 => x"00",
          9373 => x"66",
          9374 => x"20",
          9375 => x"20",
          9376 => x"66",
          9377 => x"00",
          9378 => x"44",
          9379 => x"63",
          9380 => x"69",
          9381 => x"65",
          9382 => x"74",
          9383 => x"0a",
          9384 => x"20",
          9385 => x"20",
          9386 => x"41",
          9387 => x"28",
          9388 => x"58",
          9389 => x"38",
          9390 => x"0a",
          9391 => x"20",
          9392 => x"52",
          9393 => x"20",
          9394 => x"28",
          9395 => x"58",
          9396 => x"38",
          9397 => x"0a",
          9398 => x"20",
          9399 => x"53",
          9400 => x"52",
          9401 => x"28",
          9402 => x"58",
          9403 => x"38",
          9404 => x"0a",
          9405 => x"20",
          9406 => x"41",
          9407 => x"20",
          9408 => x"28",
          9409 => x"58",
          9410 => x"38",
          9411 => x"0a",
          9412 => x"20",
          9413 => x"4d",
          9414 => x"20",
          9415 => x"28",
          9416 => x"58",
          9417 => x"38",
          9418 => x"0a",
          9419 => x"20",
          9420 => x"20",
          9421 => x"44",
          9422 => x"28",
          9423 => x"69",
          9424 => x"20",
          9425 => x"32",
          9426 => x"0a",
          9427 => x"20",
          9428 => x"4d",
          9429 => x"20",
          9430 => x"28",
          9431 => x"65",
          9432 => x"20",
          9433 => x"32",
          9434 => x"0a",
          9435 => x"20",
          9436 => x"54",
          9437 => x"54",
          9438 => x"28",
          9439 => x"6e",
          9440 => x"73",
          9441 => x"32",
          9442 => x"0a",
          9443 => x"20",
          9444 => x"53",
          9445 => x"4e",
          9446 => x"55",
          9447 => x"00",
          9448 => x"20",
          9449 => x"20",
          9450 => x"0a",
          9451 => x"20",
          9452 => x"43",
          9453 => x"00",
          9454 => x"20",
          9455 => x"32",
          9456 => x"00",
          9457 => x"20",
          9458 => x"49",
          9459 => x"00",
          9460 => x"64",
          9461 => x"73",
          9462 => x"0a",
          9463 => x"20",
          9464 => x"55",
          9465 => x"73",
          9466 => x"56",
          9467 => x"6f",
          9468 => x"64",
          9469 => x"73",
          9470 => x"20",
          9471 => x"58",
          9472 => x"00",
          9473 => x"20",
          9474 => x"55",
          9475 => x"6d",
          9476 => x"20",
          9477 => x"72",
          9478 => x"64",
          9479 => x"73",
          9480 => x"20",
          9481 => x"58",
          9482 => x"00",
          9483 => x"20",
          9484 => x"61",
          9485 => x"53",
          9486 => x"74",
          9487 => x"64",
          9488 => x"73",
          9489 => x"20",
          9490 => x"20",
          9491 => x"58",
          9492 => x"00",
          9493 => x"73",
          9494 => x"00",
          9495 => x"20",
          9496 => x"55",
          9497 => x"20",
          9498 => x"20",
          9499 => x"20",
          9500 => x"20",
          9501 => x"20",
          9502 => x"20",
          9503 => x"58",
          9504 => x"00",
          9505 => x"20",
          9506 => x"73",
          9507 => x"20",
          9508 => x"63",
          9509 => x"72",
          9510 => x"20",
          9511 => x"20",
          9512 => x"20",
          9513 => x"25",
          9514 => x"4d",
          9515 => x"00",
          9516 => x"20",
          9517 => x"52",
          9518 => x"43",
          9519 => x"6b",
          9520 => x"65",
          9521 => x"20",
          9522 => x"20",
          9523 => x"20",
          9524 => x"25",
          9525 => x"4d",
          9526 => x"00",
          9527 => x"20",
          9528 => x"73",
          9529 => x"6e",
          9530 => x"44",
          9531 => x"20",
          9532 => x"63",
          9533 => x"72",
          9534 => x"20",
          9535 => x"25",
          9536 => x"4d",
          9537 => x"00",
          9538 => x"61",
          9539 => x"00",
          9540 => x"64",
          9541 => x"00",
          9542 => x"65",
          9543 => x"00",
          9544 => x"4f",
          9545 => x"4f",
          9546 => x"00",
          9547 => x"6b",
          9548 => x"6e",
          9549 => x"96",
          9550 => x"00",
          9551 => x"00",
          9552 => x"96",
          9553 => x"00",
          9554 => x"00",
          9555 => x"96",
          9556 => x"00",
          9557 => x"00",
          9558 => x"96",
          9559 => x"00",
          9560 => x"00",
          9561 => x"96",
          9562 => x"00",
          9563 => x"00",
          9564 => x"96",
          9565 => x"00",
          9566 => x"00",
          9567 => x"96",
          9568 => x"00",
          9569 => x"00",
          9570 => x"96",
          9571 => x"00",
          9572 => x"00",
          9573 => x"96",
          9574 => x"00",
          9575 => x"00",
          9576 => x"96",
          9577 => x"00",
          9578 => x"00",
          9579 => x"96",
          9580 => x"00",
          9581 => x"00",
          9582 => x"96",
          9583 => x"00",
          9584 => x"00",
          9585 => x"96",
          9586 => x"00",
          9587 => x"00",
          9588 => x"96",
          9589 => x"00",
          9590 => x"00",
          9591 => x"96",
          9592 => x"00",
          9593 => x"00",
          9594 => x"96",
          9595 => x"00",
          9596 => x"00",
          9597 => x"96",
          9598 => x"00",
          9599 => x"00",
          9600 => x"96",
          9601 => x"00",
          9602 => x"00",
          9603 => x"96",
          9604 => x"00",
          9605 => x"00",
          9606 => x"96",
          9607 => x"00",
          9608 => x"00",
          9609 => x"96",
          9610 => x"00",
          9611 => x"00",
          9612 => x"96",
          9613 => x"00",
          9614 => x"00",
          9615 => x"44",
          9616 => x"43",
          9617 => x"42",
          9618 => x"41",
          9619 => x"36",
          9620 => x"35",
          9621 => x"34",
          9622 => x"46",
          9623 => x"33",
          9624 => x"32",
          9625 => x"31",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"73",
          9638 => x"79",
          9639 => x"73",
          9640 => x"00",
          9641 => x"00",
          9642 => x"34",
          9643 => x"25",
          9644 => x"00",
          9645 => x"69",
          9646 => x"20",
          9647 => x"72",
          9648 => x"74",
          9649 => x"65",
          9650 => x"73",
          9651 => x"79",
          9652 => x"6c",
          9653 => x"6f",
          9654 => x"46",
          9655 => x"00",
          9656 => x"6e",
          9657 => x"20",
          9658 => x"6e",
          9659 => x"65",
          9660 => x"20",
          9661 => x"74",
          9662 => x"20",
          9663 => x"65",
          9664 => x"69",
          9665 => x"6c",
          9666 => x"2e",
          9667 => x"00",
          9668 => x"2b",
          9669 => x"3c",
          9670 => x"5b",
          9671 => x"00",
          9672 => x"54",
          9673 => x"54",
          9674 => x"00",
          9675 => x"90",
          9676 => x"4f",
          9677 => x"30",
          9678 => x"20",
          9679 => x"45",
          9680 => x"20",
          9681 => x"33",
          9682 => x"20",
          9683 => x"20",
          9684 => x"45",
          9685 => x"20",
          9686 => x"20",
          9687 => x"20",
          9688 => x"97",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"45",
          9693 => x"8f",
          9694 => x"45",
          9695 => x"8e",
          9696 => x"92",
          9697 => x"55",
          9698 => x"9a",
          9699 => x"9e",
          9700 => x"4f",
          9701 => x"a6",
          9702 => x"aa",
          9703 => x"ae",
          9704 => x"b2",
          9705 => x"b6",
          9706 => x"ba",
          9707 => x"be",
          9708 => x"c2",
          9709 => x"c6",
          9710 => x"ca",
          9711 => x"ce",
          9712 => x"d2",
          9713 => x"d6",
          9714 => x"da",
          9715 => x"de",
          9716 => x"e2",
          9717 => x"e6",
          9718 => x"ea",
          9719 => x"ee",
          9720 => x"f2",
          9721 => x"f6",
          9722 => x"fa",
          9723 => x"fe",
          9724 => x"2c",
          9725 => x"5d",
          9726 => x"2a",
          9727 => x"3f",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"02",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"8c",
          9739 => x"01",
          9740 => x"00",
          9741 => x"00",
          9742 => x"8c",
          9743 => x"01",
          9744 => x"00",
          9745 => x"00",
          9746 => x"8c",
          9747 => x"03",
          9748 => x"00",
          9749 => x"00",
          9750 => x"8c",
          9751 => x"03",
          9752 => x"00",
          9753 => x"00",
          9754 => x"8c",
          9755 => x"03",
          9756 => x"00",
          9757 => x"00",
          9758 => x"8c",
          9759 => x"04",
          9760 => x"00",
          9761 => x"00",
          9762 => x"8c",
          9763 => x"04",
          9764 => x"00",
          9765 => x"00",
          9766 => x"8c",
          9767 => x"04",
          9768 => x"00",
          9769 => x"00",
          9770 => x"8c",
          9771 => x"04",
          9772 => x"00",
          9773 => x"00",
          9774 => x"8c",
          9775 => x"04",
          9776 => x"00",
          9777 => x"00",
          9778 => x"8c",
          9779 => x"04",
          9780 => x"00",
          9781 => x"00",
          9782 => x"8c",
          9783 => x"04",
          9784 => x"00",
          9785 => x"00",
          9786 => x"8c",
          9787 => x"05",
          9788 => x"00",
          9789 => x"00",
          9790 => x"8c",
          9791 => x"05",
          9792 => x"00",
          9793 => x"00",
          9794 => x"8c",
          9795 => x"05",
          9796 => x"00",
          9797 => x"00",
          9798 => x"8c",
          9799 => x"05",
          9800 => x"00",
          9801 => x"00",
          9802 => x"8c",
          9803 => x"07",
          9804 => x"00",
          9805 => x"00",
          9806 => x"8c",
          9807 => x"07",
          9808 => x"00",
          9809 => x"00",
          9810 => x"8c",
          9811 => x"08",
          9812 => x"00",
          9813 => x"00",
          9814 => x"8c",
          9815 => x"08",
          9816 => x"00",
          9817 => x"00",
          9818 => x"8c",
          9819 => x"08",
          9820 => x"00",
          9821 => x"00",
          9822 => x"8c",
          9823 => x"08",
          9824 => x"00",
          9825 => x"00",
          9826 => x"8c",
          9827 => x"09",
          9828 => x"00",
          9829 => x"00",
          9830 => x"8c",
          9831 => x"09",
          9832 => x"00",
          9833 => x"00",
          9834 => x"8d",
          9835 => x"09",
          9836 => x"00",
          9837 => x"00",
          9838 => x"8d",
          9839 => x"09",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"00",
          9844 => x"7f",
          9845 => x"00",
          9846 => x"7f",
          9847 => x"00",
          9848 => x"7f",
          9849 => x"00",
          9850 => x"00",
          9851 => x"00",
          9852 => x"ff",
          9853 => x"00",
          9854 => x"00",
          9855 => x"78",
          9856 => x"00",
          9857 => x"e1",
          9858 => x"e1",
          9859 => x"e1",
          9860 => x"00",
          9861 => x"01",
          9862 => x"01",
          9863 => x"10",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"00",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"96",
          9890 => x"00",
          9891 => x"96",
          9892 => x"00",
          9893 => x"96",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"83",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"be",
           391 => x"b5",
           392 => x"d0",
           393 => x"b5",
           394 => x"83",
           395 => x"b4",
           396 => x"90",
           397 => x"b4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"82",
           404 => x"82",
           405 => x"bc",
           406 => x"b5",
           407 => x"d0",
           408 => x"b5",
           409 => x"b2",
           410 => x"b4",
           411 => x"90",
           412 => x"b4",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"82",
           419 => x"82",
           420 => x"96",
           421 => x"b5",
           422 => x"d0",
           423 => x"b5",
           424 => x"cb",
           425 => x"b4",
           426 => x"90",
           427 => x"b4",
           428 => x"f0",
           429 => x"b4",
           430 => x"90",
           431 => x"b4",
           432 => x"ce",
           433 => x"b4",
           434 => x"90",
           435 => x"b4",
           436 => x"8a",
           437 => x"b4",
           438 => x"90",
           439 => x"b4",
           440 => x"82",
           441 => x"b4",
           442 => x"90",
           443 => x"b4",
           444 => x"b5",
           445 => x"b4",
           446 => x"90",
           447 => x"b4",
           448 => x"91",
           449 => x"b4",
           450 => x"90",
           451 => x"b4",
           452 => x"82",
           453 => x"b4",
           454 => x"90",
           455 => x"b4",
           456 => x"f6",
           457 => x"b4",
           458 => x"90",
           459 => x"b4",
           460 => x"f3",
           461 => x"b4",
           462 => x"90",
           463 => x"b4",
           464 => x"91",
           465 => x"b4",
           466 => x"90",
           467 => x"b4",
           468 => x"f1",
           469 => x"b4",
           470 => x"90",
           471 => x"b4",
           472 => x"e4",
           473 => x"b4",
           474 => x"90",
           475 => x"b4",
           476 => x"b0",
           477 => x"b4",
           478 => x"90",
           479 => x"b4",
           480 => x"cf",
           481 => x"b4",
           482 => x"90",
           483 => x"b4",
           484 => x"ee",
           485 => x"b4",
           486 => x"90",
           487 => x"b4",
           488 => x"d8",
           489 => x"b4",
           490 => x"90",
           491 => x"b4",
           492 => x"be",
           493 => x"b4",
           494 => x"90",
           495 => x"b4",
           496 => x"ac",
           497 => x"b4",
           498 => x"90",
           499 => x"b4",
           500 => x"f2",
           501 => x"b4",
           502 => x"90",
           503 => x"b4",
           504 => x"ac",
           505 => x"b4",
           506 => x"90",
           507 => x"b4",
           508 => x"ad",
           509 => x"b4",
           510 => x"90",
           511 => x"b4",
           512 => x"e2",
           513 => x"b4",
           514 => x"90",
           515 => x"b4",
           516 => x"bb",
           517 => x"b4",
           518 => x"90",
           519 => x"b4",
           520 => x"e6",
           521 => x"b4",
           522 => x"90",
           523 => x"b4",
           524 => x"c9",
           525 => x"b4",
           526 => x"90",
           527 => x"b4",
           528 => x"9e",
           529 => x"b4",
           530 => x"90",
           531 => x"b4",
           532 => x"a8",
           533 => x"b4",
           534 => x"90",
           535 => x"b4",
           536 => x"ea",
           537 => x"b4",
           538 => x"90",
           539 => x"b4",
           540 => x"b0",
           541 => x"b4",
           542 => x"90",
           543 => x"b4",
           544 => x"d6",
           545 => x"b4",
           546 => x"90",
           547 => x"b4",
           548 => x"8b",
           549 => x"b4",
           550 => x"90",
           551 => x"b4",
           552 => x"f7",
           553 => x"b4",
           554 => x"90",
           555 => x"b4",
           556 => x"eb",
           557 => x"b4",
           558 => x"90",
           559 => x"b4",
           560 => x"d5",
           561 => x"b4",
           562 => x"90",
           563 => x"b4",
           564 => x"b9",
           565 => x"b4",
           566 => x"90",
           567 => x"b4",
           568 => x"b3",
           569 => x"b4",
           570 => x"90",
           571 => x"b4",
           572 => x"d7",
           573 => x"b4",
           574 => x"90",
           575 => x"b4",
           576 => x"bb",
           577 => x"b4",
           578 => x"90",
           579 => x"b4",
           580 => x"96",
           581 => x"b4",
           582 => x"90",
           583 => x"b4",
           584 => x"ff",
           585 => x"b4",
           586 => x"90",
           587 => x"b4",
           588 => x"a7",
           589 => x"b4",
           590 => x"90",
           591 => x"b4",
           592 => x"9f",
           593 => x"b4",
           594 => x"90",
           595 => x"b4",
           596 => x"e9",
           597 => x"b4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"a8",
           623 => x"84",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"b4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"b5",
           637 => x"05",
           638 => x"b5",
           639 => x"05",
           640 => x"cc",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"b4",
           652 => x"b5",
           653 => x"3d",
           654 => x"b4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"b5",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"b5",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"b5",
           675 => x"05",
           676 => x"b4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"b5",
           683 => x"05",
           684 => x"b2",
           685 => x"a8",
           686 => x"b5",
           687 => x"05",
           688 => x"b5",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"b5",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"b5",
           709 => x"05",
           710 => x"72",
           711 => x"b4",
           712 => x"08",
           713 => x"b4",
           714 => x"0c",
           715 => x"b4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"b4",
           722 => x"0d",
           723 => x"b5",
           724 => x"05",
           725 => x"b4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"b5",
           730 => x"05",
           731 => x"b4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"b4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"b4",
           756 => x"b5",
           757 => x"3d",
           758 => x"b4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"b5",
           769 => x"82",
           770 => x"f8",
           771 => x"b5",
           772 => x"05",
           773 => x"b5",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"b4",
           779 => x"0d",
           780 => x"b5",
           781 => x"05",
           782 => x"b4",
           783 => x"08",
           784 => x"8c",
           785 => x"b5",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"b4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"b4",
           804 => x"08",
           805 => x"b5",
           806 => x"05",
           807 => x"b4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"b4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"b5",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"b4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"b5",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"b5",
           863 => x"05",
           864 => x"b4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"b4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"b5",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"b4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"b5",
           889 => x"05",
           890 => x"b4",
           891 => x"33",
           892 => x"b5",
           893 => x"05",
           894 => x"b5",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"fc",
           901 => x"51",
           902 => x"72",
           903 => x"b4",
           904 => x"22",
           905 => x"51",
           906 => x"b5",
           907 => x"05",
           908 => x"b4",
           909 => x"22",
           910 => x"51",
           911 => x"b5",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"b5",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"b5",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"b4",
           930 => x"23",
           931 => x"b5",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"b4",
           938 => x"23",
           939 => x"bf",
           940 => x"b4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"b5",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"b4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"b4",
           969 => x"0c",
           970 => x"b5",
           971 => x"05",
           972 => x"b4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"b5",
           982 => x"05",
           983 => x"ad",
           984 => x"b5",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"b4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"b5",
           993 => x"05",
           994 => x"b4",
           995 => x"22",
           996 => x"b4",
           997 => x"22",
           998 => x"54",
           999 => x"b5",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"b4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"b5",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"b4",
          1020 => x"08",
          1021 => x"e3",
          1022 => x"a8",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"b4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"b4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"b4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"b5",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"b5",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"b4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"b5",
          1072 => x"05",
          1073 => x"b4",
          1074 => x"08",
          1075 => x"b4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"b5",
          1081 => x"05",
          1082 => x"39",
          1083 => x"b5",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"b4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"b4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"b5",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"b5",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"b5",
          1127 => x"b5",
          1128 => x"05",
          1129 => x"b4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"b5",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"b5",
          1147 => x"05",
          1148 => x"33",
          1149 => x"b4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"b4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"b4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"b4",
          1172 => x"08",
          1173 => x"cd",
          1174 => x"a8",
          1175 => x"b5",
          1176 => x"05",
          1177 => x"b5",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"b4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"b4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"b4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"b5",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"b5",
          1225 => x"05",
          1226 => x"b4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"b5",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"b4",
          1247 => x"33",
          1248 => x"b4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"b5",
          1252 => x"05",
          1253 => x"b4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"b5",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"b4",
          1269 => x"23",
          1270 => x"b5",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"b4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"90",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ec",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"b4",
          1313 => x"08",
          1314 => x"95",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"b4",
          1322 => x"08",
          1323 => x"95",
          1324 => x"b5",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"9c",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"d8",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"b5",
          1381 => x"05",
          1382 => x"54",
          1383 => x"b5",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"b5",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"b4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"b5",
          1397 => x"05",
          1398 => x"b5",
          1399 => x"05",
          1400 => x"f0",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"b5",
          1407 => x"05",
          1408 => x"51",
          1409 => x"b5",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"b4",
          1420 => x"08",
          1421 => x"b5",
          1422 => x"05",
          1423 => x"94",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"b5",
          1430 => x"05",
          1431 => x"51",
          1432 => x"b5",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"c8",
          1443 => x"b4",
          1444 => x"08",
          1445 => x"b5",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"b4",
          1452 => x"08",
          1453 => x"b4",
          1454 => x"08",
          1455 => x"b5",
          1456 => x"05",
          1457 => x"b4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"b4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"b5",
          1479 => x"05",
          1480 => x"b5",
          1481 => x"05",
          1482 => x"a8",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"b4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"b4",
          1496 => x"34",
          1497 => x"b5",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"b5",
          1506 => x"05",
          1507 => x"08",
          1508 => x"b4",
          1509 => x"0c",
          1510 => x"b5",
          1511 => x"05",
          1512 => x"a8",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"b4",
          1516 => x"b5",
          1517 => x"3d",
          1518 => x"82",
          1519 => x"f0",
          1520 => x"b5",
          1521 => x"05",
          1522 => x"73",
          1523 => x"b4",
          1524 => x"08",
          1525 => x"53",
          1526 => x"72",
          1527 => x"08",
          1528 => x"72",
          1529 => x"53",
          1530 => x"09",
          1531 => x"38",
          1532 => x"08",
          1533 => x"70",
          1534 => x"71",
          1535 => x"39",
          1536 => x"08",
          1537 => x"53",
          1538 => x"09",
          1539 => x"38",
          1540 => x"b5",
          1541 => x"05",
          1542 => x"b4",
          1543 => x"08",
          1544 => x"05",
          1545 => x"08",
          1546 => x"33",
          1547 => x"08",
          1548 => x"82",
          1549 => x"f8",
          1550 => x"72",
          1551 => x"81",
          1552 => x"38",
          1553 => x"08",
          1554 => x"70",
          1555 => x"71",
          1556 => x"51",
          1557 => x"82",
          1558 => x"f8",
          1559 => x"b5",
          1560 => x"05",
          1561 => x"b4",
          1562 => x"0c",
          1563 => x"08",
          1564 => x"80",
          1565 => x"38",
          1566 => x"08",
          1567 => x"80",
          1568 => x"38",
          1569 => x"90",
          1570 => x"b4",
          1571 => x"34",
          1572 => x"08",
          1573 => x"70",
          1574 => x"71",
          1575 => x"51",
          1576 => x"82",
          1577 => x"f8",
          1578 => x"a4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"b5",
          1582 => x"05",
          1583 => x"81",
          1584 => x"70",
          1585 => x"72",
          1586 => x"b4",
          1587 => x"34",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"72",
          1591 => x"38",
          1592 => x"b5",
          1593 => x"05",
          1594 => x"39",
          1595 => x"08",
          1596 => x"53",
          1597 => x"90",
          1598 => x"b4",
          1599 => x"33",
          1600 => x"26",
          1601 => x"39",
          1602 => x"b5",
          1603 => x"05",
          1604 => x"39",
          1605 => x"b5",
          1606 => x"05",
          1607 => x"82",
          1608 => x"f8",
          1609 => x"af",
          1610 => x"38",
          1611 => x"08",
          1612 => x"53",
          1613 => x"83",
          1614 => x"80",
          1615 => x"b4",
          1616 => x"0c",
          1617 => x"8a",
          1618 => x"b4",
          1619 => x"34",
          1620 => x"b5",
          1621 => x"05",
          1622 => x"b4",
          1623 => x"33",
          1624 => x"27",
          1625 => x"82",
          1626 => x"f8",
          1627 => x"80",
          1628 => x"94",
          1629 => x"b4",
          1630 => x"33",
          1631 => x"53",
          1632 => x"b4",
          1633 => x"34",
          1634 => x"08",
          1635 => x"d0",
          1636 => x"72",
          1637 => x"08",
          1638 => x"82",
          1639 => x"f8",
          1640 => x"90",
          1641 => x"38",
          1642 => x"08",
          1643 => x"f9",
          1644 => x"72",
          1645 => x"08",
          1646 => x"82",
          1647 => x"f8",
          1648 => x"72",
          1649 => x"38",
          1650 => x"b5",
          1651 => x"05",
          1652 => x"39",
          1653 => x"08",
          1654 => x"82",
          1655 => x"f4",
          1656 => x"54",
          1657 => x"8d",
          1658 => x"82",
          1659 => x"ec",
          1660 => x"f7",
          1661 => x"b4",
          1662 => x"33",
          1663 => x"b4",
          1664 => x"08",
          1665 => x"b4",
          1666 => x"33",
          1667 => x"b5",
          1668 => x"05",
          1669 => x"b4",
          1670 => x"08",
          1671 => x"05",
          1672 => x"08",
          1673 => x"55",
          1674 => x"82",
          1675 => x"f8",
          1676 => x"a5",
          1677 => x"b4",
          1678 => x"33",
          1679 => x"2e",
          1680 => x"b5",
          1681 => x"05",
          1682 => x"b5",
          1683 => x"05",
          1684 => x"b4",
          1685 => x"08",
          1686 => x"08",
          1687 => x"71",
          1688 => x"0b",
          1689 => x"08",
          1690 => x"82",
          1691 => x"ec",
          1692 => x"b5",
          1693 => x"3d",
          1694 => x"b4",
          1695 => x"b5",
          1696 => x"82",
          1697 => x"fd",
          1698 => x"cc",
          1699 => x"82",
          1700 => x"8c",
          1701 => x"82",
          1702 => x"88",
          1703 => x"df",
          1704 => x"b5",
          1705 => x"82",
          1706 => x"54",
          1707 => x"82",
          1708 => x"04",
          1709 => x"08",
          1710 => x"b4",
          1711 => x"0d",
          1712 => x"b5",
          1713 => x"05",
          1714 => x"b4",
          1715 => x"08",
          1716 => x"0c",
          1717 => x"08",
          1718 => x"70",
          1719 => x"72",
          1720 => x"82",
          1721 => x"f8",
          1722 => x"81",
          1723 => x"72",
          1724 => x"81",
          1725 => x"82",
          1726 => x"88",
          1727 => x"08",
          1728 => x"0c",
          1729 => x"82",
          1730 => x"f8",
          1731 => x"72",
          1732 => x"81",
          1733 => x"81",
          1734 => x"b4",
          1735 => x"34",
          1736 => x"08",
          1737 => x"70",
          1738 => x"71",
          1739 => x"51",
          1740 => x"82",
          1741 => x"f8",
          1742 => x"b5",
          1743 => x"05",
          1744 => x"b0",
          1745 => x"06",
          1746 => x"82",
          1747 => x"88",
          1748 => x"08",
          1749 => x"0c",
          1750 => x"53",
          1751 => x"b5",
          1752 => x"05",
          1753 => x"b4",
          1754 => x"33",
          1755 => x"08",
          1756 => x"82",
          1757 => x"e8",
          1758 => x"e2",
          1759 => x"82",
          1760 => x"e8",
          1761 => x"f8",
          1762 => x"80",
          1763 => x"0b",
          1764 => x"08",
          1765 => x"82",
          1766 => x"88",
          1767 => x"08",
          1768 => x"0c",
          1769 => x"53",
          1770 => x"b5",
          1771 => x"05",
          1772 => x"39",
          1773 => x"b5",
          1774 => x"05",
          1775 => x"b4",
          1776 => x"08",
          1777 => x"05",
          1778 => x"08",
          1779 => x"33",
          1780 => x"08",
          1781 => x"80",
          1782 => x"b5",
          1783 => x"05",
          1784 => x"a0",
          1785 => x"81",
          1786 => x"b4",
          1787 => x"0c",
          1788 => x"82",
          1789 => x"f8",
          1790 => x"af",
          1791 => x"38",
          1792 => x"08",
          1793 => x"53",
          1794 => x"83",
          1795 => x"80",
          1796 => x"b4",
          1797 => x"0c",
          1798 => x"88",
          1799 => x"b4",
          1800 => x"34",
          1801 => x"b5",
          1802 => x"05",
          1803 => x"73",
          1804 => x"82",
          1805 => x"f8",
          1806 => x"72",
          1807 => x"38",
          1808 => x"0b",
          1809 => x"08",
          1810 => x"82",
          1811 => x"0b",
          1812 => x"08",
          1813 => x"80",
          1814 => x"b4",
          1815 => x"0c",
          1816 => x"08",
          1817 => x"53",
          1818 => x"81",
          1819 => x"b5",
          1820 => x"05",
          1821 => x"e0",
          1822 => x"38",
          1823 => x"08",
          1824 => x"e0",
          1825 => x"72",
          1826 => x"08",
          1827 => x"82",
          1828 => x"f8",
          1829 => x"11",
          1830 => x"82",
          1831 => x"f8",
          1832 => x"b5",
          1833 => x"05",
          1834 => x"73",
          1835 => x"82",
          1836 => x"f8",
          1837 => x"11",
          1838 => x"82",
          1839 => x"f8",
          1840 => x"b5",
          1841 => x"05",
          1842 => x"89",
          1843 => x"80",
          1844 => x"b4",
          1845 => x"0c",
          1846 => x"82",
          1847 => x"f8",
          1848 => x"b5",
          1849 => x"05",
          1850 => x"72",
          1851 => x"38",
          1852 => x"b5",
          1853 => x"05",
          1854 => x"39",
          1855 => x"08",
          1856 => x"70",
          1857 => x"08",
          1858 => x"29",
          1859 => x"08",
          1860 => x"70",
          1861 => x"b4",
          1862 => x"0c",
          1863 => x"08",
          1864 => x"70",
          1865 => x"71",
          1866 => x"51",
          1867 => x"53",
          1868 => x"b5",
          1869 => x"05",
          1870 => x"39",
          1871 => x"08",
          1872 => x"53",
          1873 => x"90",
          1874 => x"b4",
          1875 => x"08",
          1876 => x"b4",
          1877 => x"0c",
          1878 => x"08",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"0c",
          1882 => x"82",
          1883 => x"ec",
          1884 => x"b5",
          1885 => x"05",
          1886 => x"a8",
          1887 => x"0d",
          1888 => x"0c",
          1889 => x"b4",
          1890 => x"b5",
          1891 => x"3d",
          1892 => x"82",
          1893 => x"f8",
          1894 => x"cc",
          1895 => x"11",
          1896 => x"2a",
          1897 => x"70",
          1898 => x"51",
          1899 => x"72",
          1900 => x"38",
          1901 => x"b5",
          1902 => x"05",
          1903 => x"39",
          1904 => x"08",
          1905 => x"53",
          1906 => x"b5",
          1907 => x"05",
          1908 => x"82",
          1909 => x"88",
          1910 => x"72",
          1911 => x"08",
          1912 => x"72",
          1913 => x"53",
          1914 => x"b0",
          1915 => x"fc",
          1916 => x"fc",
          1917 => x"b5",
          1918 => x"05",
          1919 => x"11",
          1920 => x"72",
          1921 => x"a8",
          1922 => x"80",
          1923 => x"38",
          1924 => x"b5",
          1925 => x"05",
          1926 => x"39",
          1927 => x"08",
          1928 => x"08",
          1929 => x"51",
          1930 => x"53",
          1931 => x"b5",
          1932 => x"72",
          1933 => x"38",
          1934 => x"b5",
          1935 => x"05",
          1936 => x"b4",
          1937 => x"08",
          1938 => x"b4",
          1939 => x"0c",
          1940 => x"b4",
          1941 => x"08",
          1942 => x"0c",
          1943 => x"82",
          1944 => x"04",
          1945 => x"08",
          1946 => x"b4",
          1947 => x"0d",
          1948 => x"b5",
          1949 => x"05",
          1950 => x"b4",
          1951 => x"08",
          1952 => x"70",
          1953 => x"81",
          1954 => x"06",
          1955 => x"51",
          1956 => x"2e",
          1957 => x"0b",
          1958 => x"08",
          1959 => x"80",
          1960 => x"b5",
          1961 => x"05",
          1962 => x"33",
          1963 => x"08",
          1964 => x"81",
          1965 => x"b4",
          1966 => x"0c",
          1967 => x"b5",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"82",
          1972 => x"8c",
          1973 => x"b5",
          1974 => x"05",
          1975 => x"b5",
          1976 => x"05",
          1977 => x"11",
          1978 => x"72",
          1979 => x"a8",
          1980 => x"80",
          1981 => x"38",
          1982 => x"b5",
          1983 => x"05",
          1984 => x"39",
          1985 => x"08",
          1986 => x"70",
          1987 => x"08",
          1988 => x"53",
          1989 => x"08",
          1990 => x"82",
          1991 => x"87",
          1992 => x"b5",
          1993 => x"82",
          1994 => x"02",
          1995 => x"0c",
          1996 => x"82",
          1997 => x"52",
          1998 => x"08",
          1999 => x"51",
          2000 => x"b5",
          2001 => x"82",
          2002 => x"53",
          2003 => x"82",
          2004 => x"04",
          2005 => x"08",
          2006 => x"b4",
          2007 => x"0d",
          2008 => x"08",
          2009 => x"85",
          2010 => x"81",
          2011 => x"32",
          2012 => x"51",
          2013 => x"53",
          2014 => x"8d",
          2015 => x"82",
          2016 => x"fc",
          2017 => x"cb",
          2018 => x"b4",
          2019 => x"08",
          2020 => x"70",
          2021 => x"81",
          2022 => x"51",
          2023 => x"2e",
          2024 => x"82",
          2025 => x"8c",
          2026 => x"b5",
          2027 => x"05",
          2028 => x"8c",
          2029 => x"14",
          2030 => x"38",
          2031 => x"08",
          2032 => x"70",
          2033 => x"b5",
          2034 => x"05",
          2035 => x"54",
          2036 => x"34",
          2037 => x"05",
          2038 => x"b5",
          2039 => x"05",
          2040 => x"08",
          2041 => x"12",
          2042 => x"b4",
          2043 => x"08",
          2044 => x"b4",
          2045 => x"0c",
          2046 => x"d7",
          2047 => x"b4",
          2048 => x"08",
          2049 => x"08",
          2050 => x"53",
          2051 => x"08",
          2052 => x"70",
          2053 => x"53",
          2054 => x"51",
          2055 => x"2d",
          2056 => x"08",
          2057 => x"38",
          2058 => x"08",
          2059 => x"8c",
          2060 => x"05",
          2061 => x"82",
          2062 => x"88",
          2063 => x"82",
          2064 => x"fc",
          2065 => x"53",
          2066 => x"0b",
          2067 => x"08",
          2068 => x"82",
          2069 => x"fc",
          2070 => x"b5",
          2071 => x"3d",
          2072 => x"b4",
          2073 => x"b5",
          2074 => x"82",
          2075 => x"f9",
          2076 => x"b5",
          2077 => x"05",
          2078 => x"33",
          2079 => x"70",
          2080 => x"51",
          2081 => x"80",
          2082 => x"ff",
          2083 => x"b4",
          2084 => x"0c",
          2085 => x"82",
          2086 => x"88",
          2087 => x"11",
          2088 => x"2a",
          2089 => x"51",
          2090 => x"71",
          2091 => x"c5",
          2092 => x"b4",
          2093 => x"08",
          2094 => x"08",
          2095 => x"53",
          2096 => x"33",
          2097 => x"06",
          2098 => x"85",
          2099 => x"b5",
          2100 => x"05",
          2101 => x"08",
          2102 => x"12",
          2103 => x"b4",
          2104 => x"08",
          2105 => x"70",
          2106 => x"08",
          2107 => x"51",
          2108 => x"b6",
          2109 => x"b4",
          2110 => x"08",
          2111 => x"70",
          2112 => x"81",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"82",
          2116 => x"88",
          2117 => x"08",
          2118 => x"b5",
          2119 => x"05",
          2120 => x"82",
          2121 => x"fc",
          2122 => x"38",
          2123 => x"08",
          2124 => x"82",
          2125 => x"88",
          2126 => x"53",
          2127 => x"70",
          2128 => x"52",
          2129 => x"34",
          2130 => x"b5",
          2131 => x"05",
          2132 => x"39",
          2133 => x"08",
          2134 => x"70",
          2135 => x"71",
          2136 => x"a1",
          2137 => x"b4",
          2138 => x"08",
          2139 => x"08",
          2140 => x"52",
          2141 => x"51",
          2142 => x"82",
          2143 => x"70",
          2144 => x"08",
          2145 => x"52",
          2146 => x"08",
          2147 => x"80",
          2148 => x"38",
          2149 => x"08",
          2150 => x"82",
          2151 => x"f4",
          2152 => x"b5",
          2153 => x"05",
          2154 => x"33",
          2155 => x"08",
          2156 => x"52",
          2157 => x"08",
          2158 => x"ff",
          2159 => x"06",
          2160 => x"b5",
          2161 => x"05",
          2162 => x"52",
          2163 => x"b4",
          2164 => x"34",
          2165 => x"b5",
          2166 => x"05",
          2167 => x"52",
          2168 => x"b4",
          2169 => x"34",
          2170 => x"08",
          2171 => x"52",
          2172 => x"08",
          2173 => x"85",
          2174 => x"0b",
          2175 => x"08",
          2176 => x"a6",
          2177 => x"b4",
          2178 => x"08",
          2179 => x"81",
          2180 => x"0c",
          2181 => x"08",
          2182 => x"70",
          2183 => x"70",
          2184 => x"08",
          2185 => x"51",
          2186 => x"b5",
          2187 => x"05",
          2188 => x"a8",
          2189 => x"0d",
          2190 => x"0c",
          2191 => x"b4",
          2192 => x"b5",
          2193 => x"3d",
          2194 => x"b4",
          2195 => x"08",
          2196 => x"08",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"b5",
          2200 => x"05",
          2201 => x"b4",
          2202 => x"08",
          2203 => x"a2",
          2204 => x"b4",
          2205 => x"08",
          2206 => x"08",
          2207 => x"26",
          2208 => x"82",
          2209 => x"f8",
          2210 => x"b5",
          2211 => x"05",
          2212 => x"82",
          2213 => x"fc",
          2214 => x"27",
          2215 => x"82",
          2216 => x"fc",
          2217 => x"b5",
          2218 => x"05",
          2219 => x"b5",
          2220 => x"05",
          2221 => x"b4",
          2222 => x"08",
          2223 => x"08",
          2224 => x"05",
          2225 => x"08",
          2226 => x"82",
          2227 => x"90",
          2228 => x"05",
          2229 => x"08",
          2230 => x"82",
          2231 => x"90",
          2232 => x"05",
          2233 => x"08",
          2234 => x"82",
          2235 => x"90",
          2236 => x"2e",
          2237 => x"82",
          2238 => x"fc",
          2239 => x"05",
          2240 => x"08",
          2241 => x"82",
          2242 => x"f8",
          2243 => x"05",
          2244 => x"08",
          2245 => x"82",
          2246 => x"fc",
          2247 => x"b5",
          2248 => x"05",
          2249 => x"71",
          2250 => x"ff",
          2251 => x"b5",
          2252 => x"05",
          2253 => x"82",
          2254 => x"90",
          2255 => x"b5",
          2256 => x"05",
          2257 => x"82",
          2258 => x"90",
          2259 => x"b5",
          2260 => x"05",
          2261 => x"ba",
          2262 => x"b4",
          2263 => x"08",
          2264 => x"82",
          2265 => x"f8",
          2266 => x"05",
          2267 => x"08",
          2268 => x"82",
          2269 => x"fc",
          2270 => x"52",
          2271 => x"82",
          2272 => x"fc",
          2273 => x"05",
          2274 => x"08",
          2275 => x"ff",
          2276 => x"b5",
          2277 => x"05",
          2278 => x"b5",
          2279 => x"85",
          2280 => x"b5",
          2281 => x"82",
          2282 => x"02",
          2283 => x"0c",
          2284 => x"82",
          2285 => x"88",
          2286 => x"b5",
          2287 => x"05",
          2288 => x"b4",
          2289 => x"08",
          2290 => x"82",
          2291 => x"fc",
          2292 => x"05",
          2293 => x"08",
          2294 => x"70",
          2295 => x"51",
          2296 => x"2e",
          2297 => x"39",
          2298 => x"08",
          2299 => x"ff",
          2300 => x"b4",
          2301 => x"0c",
          2302 => x"08",
          2303 => x"82",
          2304 => x"88",
          2305 => x"70",
          2306 => x"0c",
          2307 => x"0d",
          2308 => x"0c",
          2309 => x"b4",
          2310 => x"b5",
          2311 => x"3d",
          2312 => x"b4",
          2313 => x"08",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"71",
          2318 => x"b4",
          2319 => x"08",
          2320 => x"b5",
          2321 => x"05",
          2322 => x"b4",
          2323 => x"08",
          2324 => x"72",
          2325 => x"b4",
          2326 => x"08",
          2327 => x"b5",
          2328 => x"05",
          2329 => x"ff",
          2330 => x"80",
          2331 => x"ff",
          2332 => x"b5",
          2333 => x"05",
          2334 => x"b5",
          2335 => x"84",
          2336 => x"b5",
          2337 => x"82",
          2338 => x"02",
          2339 => x"0c",
          2340 => x"82",
          2341 => x"88",
          2342 => x"b5",
          2343 => x"05",
          2344 => x"b4",
          2345 => x"08",
          2346 => x"08",
          2347 => x"82",
          2348 => x"90",
          2349 => x"2e",
          2350 => x"82",
          2351 => x"90",
          2352 => x"05",
          2353 => x"08",
          2354 => x"82",
          2355 => x"90",
          2356 => x"05",
          2357 => x"08",
          2358 => x"82",
          2359 => x"90",
          2360 => x"2e",
          2361 => x"b5",
          2362 => x"05",
          2363 => x"33",
          2364 => x"08",
          2365 => x"81",
          2366 => x"b4",
          2367 => x"0c",
          2368 => x"08",
          2369 => x"52",
          2370 => x"34",
          2371 => x"08",
          2372 => x"81",
          2373 => x"b4",
          2374 => x"0c",
          2375 => x"82",
          2376 => x"88",
          2377 => x"82",
          2378 => x"51",
          2379 => x"82",
          2380 => x"04",
          2381 => x"08",
          2382 => x"b4",
          2383 => x"0d",
          2384 => x"08",
          2385 => x"80",
          2386 => x"38",
          2387 => x"08",
          2388 => x"52",
          2389 => x"b5",
          2390 => x"05",
          2391 => x"82",
          2392 => x"8c",
          2393 => x"b5",
          2394 => x"05",
          2395 => x"72",
          2396 => x"53",
          2397 => x"71",
          2398 => x"38",
          2399 => x"82",
          2400 => x"88",
          2401 => x"71",
          2402 => x"b4",
          2403 => x"08",
          2404 => x"b5",
          2405 => x"05",
          2406 => x"ff",
          2407 => x"70",
          2408 => x"0b",
          2409 => x"08",
          2410 => x"81",
          2411 => x"b5",
          2412 => x"05",
          2413 => x"82",
          2414 => x"90",
          2415 => x"b5",
          2416 => x"05",
          2417 => x"84",
          2418 => x"39",
          2419 => x"08",
          2420 => x"80",
          2421 => x"38",
          2422 => x"08",
          2423 => x"70",
          2424 => x"70",
          2425 => x"0b",
          2426 => x"08",
          2427 => x"80",
          2428 => x"b5",
          2429 => x"05",
          2430 => x"82",
          2431 => x"8c",
          2432 => x"b5",
          2433 => x"05",
          2434 => x"52",
          2435 => x"38",
          2436 => x"b5",
          2437 => x"05",
          2438 => x"82",
          2439 => x"88",
          2440 => x"33",
          2441 => x"08",
          2442 => x"70",
          2443 => x"31",
          2444 => x"b4",
          2445 => x"0c",
          2446 => x"52",
          2447 => x"80",
          2448 => x"b4",
          2449 => x"0c",
          2450 => x"08",
          2451 => x"82",
          2452 => x"85",
          2453 => x"b5",
          2454 => x"82",
          2455 => x"02",
          2456 => x"0c",
          2457 => x"82",
          2458 => x"88",
          2459 => x"b5",
          2460 => x"05",
          2461 => x"b4",
          2462 => x"08",
          2463 => x"0b",
          2464 => x"08",
          2465 => x"80",
          2466 => x"b5",
          2467 => x"05",
          2468 => x"33",
          2469 => x"08",
          2470 => x"81",
          2471 => x"b4",
          2472 => x"0c",
          2473 => x"06",
          2474 => x"80",
          2475 => x"82",
          2476 => x"8c",
          2477 => x"05",
          2478 => x"08",
          2479 => x"82",
          2480 => x"8c",
          2481 => x"2e",
          2482 => x"be",
          2483 => x"b4",
          2484 => x"08",
          2485 => x"b5",
          2486 => x"05",
          2487 => x"b4",
          2488 => x"08",
          2489 => x"08",
          2490 => x"31",
          2491 => x"b4",
          2492 => x"0c",
          2493 => x"b4",
          2494 => x"08",
          2495 => x"0c",
          2496 => x"82",
          2497 => x"04",
          2498 => x"08",
          2499 => x"b4",
          2500 => x"0d",
          2501 => x"08",
          2502 => x"82",
          2503 => x"fc",
          2504 => x"b5",
          2505 => x"05",
          2506 => x"80",
          2507 => x"b5",
          2508 => x"05",
          2509 => x"82",
          2510 => x"90",
          2511 => x"b5",
          2512 => x"05",
          2513 => x"82",
          2514 => x"90",
          2515 => x"b5",
          2516 => x"05",
          2517 => x"a9",
          2518 => x"b4",
          2519 => x"08",
          2520 => x"b5",
          2521 => x"05",
          2522 => x"71",
          2523 => x"b5",
          2524 => x"05",
          2525 => x"82",
          2526 => x"fc",
          2527 => x"be",
          2528 => x"b4",
          2529 => x"08",
          2530 => x"a8",
          2531 => x"3d",
          2532 => x"b4",
          2533 => x"b5",
          2534 => x"82",
          2535 => x"f9",
          2536 => x"0b",
          2537 => x"08",
          2538 => x"82",
          2539 => x"88",
          2540 => x"25",
          2541 => x"b5",
          2542 => x"05",
          2543 => x"b5",
          2544 => x"05",
          2545 => x"82",
          2546 => x"f4",
          2547 => x"b5",
          2548 => x"05",
          2549 => x"81",
          2550 => x"b4",
          2551 => x"0c",
          2552 => x"08",
          2553 => x"82",
          2554 => x"fc",
          2555 => x"b5",
          2556 => x"05",
          2557 => x"b9",
          2558 => x"b4",
          2559 => x"08",
          2560 => x"b4",
          2561 => x"0c",
          2562 => x"b5",
          2563 => x"05",
          2564 => x"b4",
          2565 => x"08",
          2566 => x"0b",
          2567 => x"08",
          2568 => x"82",
          2569 => x"f0",
          2570 => x"b5",
          2571 => x"05",
          2572 => x"82",
          2573 => x"8c",
          2574 => x"82",
          2575 => x"88",
          2576 => x"82",
          2577 => x"b5",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"82",
          2581 => x"fc",
          2582 => x"2e",
          2583 => x"b5",
          2584 => x"05",
          2585 => x"b5",
          2586 => x"05",
          2587 => x"b4",
          2588 => x"08",
          2589 => x"a8",
          2590 => x"3d",
          2591 => x"b4",
          2592 => x"b5",
          2593 => x"82",
          2594 => x"fb",
          2595 => x"0b",
          2596 => x"08",
          2597 => x"82",
          2598 => x"88",
          2599 => x"25",
          2600 => x"b5",
          2601 => x"05",
          2602 => x"b5",
          2603 => x"05",
          2604 => x"82",
          2605 => x"fc",
          2606 => x"b5",
          2607 => x"05",
          2608 => x"90",
          2609 => x"b4",
          2610 => x"08",
          2611 => x"b4",
          2612 => x"0c",
          2613 => x"b5",
          2614 => x"05",
          2615 => x"b5",
          2616 => x"05",
          2617 => x"a2",
          2618 => x"a8",
          2619 => x"b5",
          2620 => x"05",
          2621 => x"b5",
          2622 => x"05",
          2623 => x"90",
          2624 => x"b4",
          2625 => x"08",
          2626 => x"b4",
          2627 => x"0c",
          2628 => x"08",
          2629 => x"70",
          2630 => x"0c",
          2631 => x"0d",
          2632 => x"0c",
          2633 => x"b4",
          2634 => x"b5",
          2635 => x"3d",
          2636 => x"82",
          2637 => x"8c",
          2638 => x"82",
          2639 => x"88",
          2640 => x"80",
          2641 => x"b5",
          2642 => x"82",
          2643 => x"54",
          2644 => x"82",
          2645 => x"04",
          2646 => x"08",
          2647 => x"b4",
          2648 => x"0d",
          2649 => x"b5",
          2650 => x"05",
          2651 => x"b5",
          2652 => x"05",
          2653 => x"3f",
          2654 => x"08",
          2655 => x"a8",
          2656 => x"3d",
          2657 => x"b4",
          2658 => x"b5",
          2659 => x"82",
          2660 => x"fd",
          2661 => x"0b",
          2662 => x"08",
          2663 => x"80",
          2664 => x"b4",
          2665 => x"0c",
          2666 => x"08",
          2667 => x"82",
          2668 => x"88",
          2669 => x"b9",
          2670 => x"b4",
          2671 => x"08",
          2672 => x"38",
          2673 => x"b5",
          2674 => x"05",
          2675 => x"38",
          2676 => x"08",
          2677 => x"10",
          2678 => x"08",
          2679 => x"82",
          2680 => x"fc",
          2681 => x"82",
          2682 => x"fc",
          2683 => x"b8",
          2684 => x"b4",
          2685 => x"08",
          2686 => x"e1",
          2687 => x"b4",
          2688 => x"08",
          2689 => x"08",
          2690 => x"26",
          2691 => x"b5",
          2692 => x"05",
          2693 => x"b4",
          2694 => x"08",
          2695 => x"b4",
          2696 => x"0c",
          2697 => x"08",
          2698 => x"82",
          2699 => x"fc",
          2700 => x"82",
          2701 => x"f8",
          2702 => x"b5",
          2703 => x"05",
          2704 => x"82",
          2705 => x"fc",
          2706 => x"b5",
          2707 => x"05",
          2708 => x"82",
          2709 => x"8c",
          2710 => x"95",
          2711 => x"b4",
          2712 => x"08",
          2713 => x"38",
          2714 => x"08",
          2715 => x"70",
          2716 => x"08",
          2717 => x"51",
          2718 => x"b5",
          2719 => x"05",
          2720 => x"b5",
          2721 => x"05",
          2722 => x"b5",
          2723 => x"05",
          2724 => x"a8",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"f3",
          2733 => x"a8",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"94",
          2762 => x"71",
          2763 => x"9a",
          2764 => x"80",
          2765 => x"98",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"9a",
          2771 => x"e4",
          2772 => x"e0",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"9b",
          2778 => x"c8",
          2779 => x"b4",
          2780 => x"39",
          2781 => x"51",
          2782 => x"9b",
          2783 => x"39",
          2784 => x"51",
          2785 => x"9c",
          2786 => x"39",
          2787 => x"51",
          2788 => x"9c",
          2789 => x"39",
          2790 => x"51",
          2791 => x"9d",
          2792 => x"39",
          2793 => x"51",
          2794 => x"9d",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"cd",
          2806 => x"a8",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"a8",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"98",
          2840 => x"a8",
          2841 => x"b5",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"a8",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"58",
          2864 => x"80",
          2865 => x"7a",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"80",
          2869 => x"76",
          2870 => x"38",
          2871 => x"56",
          2872 => x"54",
          2873 => x"53",
          2874 => x"51",
          2875 => x"b5",
          2876 => x"83",
          2877 => x"77",
          2878 => x"0c",
          2879 => x"04",
          2880 => x"7f",
          2881 => x"8c",
          2882 => x"05",
          2883 => x"15",
          2884 => x"5c",
          2885 => x"5e",
          2886 => x"9e",
          2887 => x"b9",
          2888 => x"9e",
          2889 => x"dd",
          2890 => x"74",
          2891 => x"fd",
          2892 => x"2e",
          2893 => x"a0",
          2894 => x"80",
          2895 => x"18",
          2896 => x"27",
          2897 => x"22",
          2898 => x"8c",
          2899 => x"88",
          2900 => x"82",
          2901 => x"e0",
          2902 => x"15",
          2903 => x"39",
          2904 => x"72",
          2905 => x"38",
          2906 => x"82",
          2907 => x"ff",
          2908 => x"88",
          2909 => x"94",
          2910 => x"3f",
          2911 => x"a0",
          2912 => x"53",
          2913 => x"8e",
          2914 => x"52",
          2915 => x"51",
          2916 => x"3f",
          2917 => x"9e",
          2918 => x"e9",
          2919 => x"55",
          2920 => x"08",
          2921 => x"e3",
          2922 => x"ff",
          2923 => x"ac",
          2924 => x"3f",
          2925 => x"79",
          2926 => x"38",
          2927 => x"33",
          2928 => x"56",
          2929 => x"83",
          2930 => x"80",
          2931 => x"27",
          2932 => x"53",
          2933 => x"70",
          2934 => x"51",
          2935 => x"2e",
          2936 => x"80",
          2937 => x"38",
          2938 => x"08",
          2939 => x"88",
          2940 => x"fc",
          2941 => x"51",
          2942 => x"81",
          2943 => x"b6",
          2944 => x"b0",
          2945 => x"3f",
          2946 => x"1c",
          2947 => x"c0",
          2948 => x"a8",
          2949 => x"70",
          2950 => x"57",
          2951 => x"09",
          2952 => x"38",
          2953 => x"82",
          2954 => x"98",
          2955 => x"2c",
          2956 => x"70",
          2957 => x"32",
          2958 => x"72",
          2959 => x"07",
          2960 => x"58",
          2961 => x"57",
          2962 => x"d8",
          2963 => x"2e",
          2964 => x"85",
          2965 => x"8c",
          2966 => x"53",
          2967 => x"fd",
          2968 => x"53",
          2969 => x"a8",
          2970 => x"0d",
          2971 => x"0d",
          2972 => x"33",
          2973 => x"53",
          2974 => x"52",
          2975 => x"d8",
          2976 => x"80",
          2977 => x"9b",
          2978 => x"c4",
          2979 => x"d0",
          2980 => x"81",
          2981 => x"9e",
          2982 => x"b6",
          2983 => x"80",
          2984 => x"a0",
          2985 => x"3d",
          2986 => x"3d",
          2987 => x"96",
          2988 => x"a5",
          2989 => x"51",
          2990 => x"82",
          2991 => x"99",
          2992 => x"51",
          2993 => x"72",
          2994 => x"81",
          2995 => x"71",
          2996 => x"38",
          2997 => x"e5",
          2998 => x"8c",
          2999 => x"3f",
          3000 => x"d9",
          3001 => x"2a",
          3002 => x"51",
          3003 => x"2e",
          3004 => x"51",
          3005 => x"82",
          3006 => x"98",
          3007 => x"51",
          3008 => x"72",
          3009 => x"81",
          3010 => x"71",
          3011 => x"38",
          3012 => x"a9",
          3013 => x"b0",
          3014 => x"3f",
          3015 => x"9d",
          3016 => x"2a",
          3017 => x"51",
          3018 => x"2e",
          3019 => x"51",
          3020 => x"82",
          3021 => x"98",
          3022 => x"51",
          3023 => x"72",
          3024 => x"81",
          3025 => x"71",
          3026 => x"38",
          3027 => x"ed",
          3028 => x"d8",
          3029 => x"3f",
          3030 => x"e1",
          3031 => x"2a",
          3032 => x"51",
          3033 => x"2e",
          3034 => x"51",
          3035 => x"82",
          3036 => x"97",
          3037 => x"51",
          3038 => x"72",
          3039 => x"81",
          3040 => x"71",
          3041 => x"38",
          3042 => x"b1",
          3043 => x"80",
          3044 => x"3f",
          3045 => x"a5",
          3046 => x"2a",
          3047 => x"51",
          3048 => x"2e",
          3049 => x"51",
          3050 => x"82",
          3051 => x"97",
          3052 => x"51",
          3053 => x"a3",
          3054 => x"3d",
          3055 => x"3d",
          3056 => x"84",
          3057 => x"33",
          3058 => x"56",
          3059 => x"51",
          3060 => x"0b",
          3061 => x"a4",
          3062 => x"a9",
          3063 => x"82",
          3064 => x"82",
          3065 => x"80",
          3066 => x"82",
          3067 => x"30",
          3068 => x"a8",
          3069 => x"25",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"a4",
          3073 => x"82",
          3074 => x"54",
          3075 => x"09",
          3076 => x"38",
          3077 => x"53",
          3078 => x"51",
          3079 => x"3f",
          3080 => x"08",
          3081 => x"38",
          3082 => x"08",
          3083 => x"3f",
          3084 => x"cc",
          3085 => x"83",
          3086 => x"0b",
          3087 => x"b0",
          3088 => x"0b",
          3089 => x"33",
          3090 => x"2e",
          3091 => x"8c",
          3092 => x"e4",
          3093 => x"75",
          3094 => x"3f",
          3095 => x"b5",
          3096 => x"3d",
          3097 => x"3d",
          3098 => x"71",
          3099 => x"0c",
          3100 => x"52",
          3101 => x"c5",
          3102 => x"b5",
          3103 => x"ff",
          3104 => x"7e",
          3105 => x"06",
          3106 => x"3d",
          3107 => x"82",
          3108 => x"79",
          3109 => x"3f",
          3110 => x"52",
          3111 => x"51",
          3112 => x"3f",
          3113 => x"08",
          3114 => x"38",
          3115 => x"51",
          3116 => x"81",
          3117 => x"82",
          3118 => x"d9",
          3119 => x"3d",
          3120 => x"80",
          3121 => x"51",
          3122 => x"b5",
          3123 => x"05",
          3124 => x"3f",
          3125 => x"08",
          3126 => x"90",
          3127 => x"79",
          3128 => x"87",
          3129 => x"80",
          3130 => x"38",
          3131 => x"81",
          3132 => x"bd",
          3133 => x"79",
          3134 => x"bb",
          3135 => x"2e",
          3136 => x"8a",
          3137 => x"80",
          3138 => x"95",
          3139 => x"c0",
          3140 => x"38",
          3141 => x"82",
          3142 => x"a9",
          3143 => x"f9",
          3144 => x"38",
          3145 => x"24",
          3146 => x"80",
          3147 => x"fa",
          3148 => x"f8",
          3149 => x"38",
          3150 => x"79",
          3151 => x"89",
          3152 => x"81",
          3153 => x"38",
          3154 => x"2e",
          3155 => x"89",
          3156 => x"81",
          3157 => x"e7",
          3158 => x"39",
          3159 => x"80",
          3160 => x"84",
          3161 => x"cc",
          3162 => x"a8",
          3163 => x"fe",
          3164 => x"3d",
          3165 => x"53",
          3166 => x"51",
          3167 => x"82",
          3168 => x"80",
          3169 => x"38",
          3170 => x"f8",
          3171 => x"84",
          3172 => x"a0",
          3173 => x"a8",
          3174 => x"82",
          3175 => x"43",
          3176 => x"51",
          3177 => x"64",
          3178 => x"7a",
          3179 => x"ea",
          3180 => x"79",
          3181 => x"05",
          3182 => x"7b",
          3183 => x"81",
          3184 => x"3d",
          3185 => x"53",
          3186 => x"51",
          3187 => x"82",
          3188 => x"80",
          3189 => x"38",
          3190 => x"fc",
          3191 => x"84",
          3192 => x"d0",
          3193 => x"a8",
          3194 => x"fd",
          3195 => x"3d",
          3196 => x"53",
          3197 => x"51",
          3198 => x"82",
          3199 => x"80",
          3200 => x"38",
          3201 => x"51",
          3202 => x"64",
          3203 => x"27",
          3204 => x"62",
          3205 => x"81",
          3206 => x"7a",
          3207 => x"05",
          3208 => x"b5",
          3209 => x"11",
          3210 => x"05",
          3211 => x"3f",
          3212 => x"08",
          3213 => x"ff",
          3214 => x"fe",
          3215 => x"ff",
          3216 => x"d0",
          3217 => x"b5",
          3218 => x"2e",
          3219 => x"b5",
          3220 => x"11",
          3221 => x"05",
          3222 => x"3f",
          3223 => x"08",
          3224 => x"d3",
          3225 => x"c8",
          3226 => x"3f",
          3227 => x"64",
          3228 => x"62",
          3229 => x"33",
          3230 => x"79",
          3231 => x"38",
          3232 => x"54",
          3233 => x"7a",
          3234 => x"d8",
          3235 => x"c8",
          3236 => x"63",
          3237 => x"5b",
          3238 => x"a1",
          3239 => x"a7",
          3240 => x"ff",
          3241 => x"ff",
          3242 => x"d0",
          3243 => x"b5",
          3244 => x"df",
          3245 => x"94",
          3246 => x"80",
          3247 => x"82",
          3248 => x"45",
          3249 => x"82",
          3250 => x"5a",
          3251 => x"88",
          3252 => x"d4",
          3253 => x"39",
          3254 => x"33",
          3255 => x"2e",
          3256 => x"b3",
          3257 => x"ab",
          3258 => x"97",
          3259 => x"80",
          3260 => x"82",
          3261 => x"45",
          3262 => x"b4",
          3263 => x"79",
          3264 => x"38",
          3265 => x"08",
          3266 => x"82",
          3267 => x"fc",
          3268 => x"b5",
          3269 => x"11",
          3270 => x"05",
          3271 => x"3f",
          3272 => x"08",
          3273 => x"82",
          3274 => x"5a",
          3275 => x"89",
          3276 => x"d0",
          3277 => x"cc",
          3278 => x"95",
          3279 => x"80",
          3280 => x"82",
          3281 => x"44",
          3282 => x"b4",
          3283 => x"79",
          3284 => x"38",
          3285 => x"08",
          3286 => x"82",
          3287 => x"5a",
          3288 => x"88",
          3289 => x"e8",
          3290 => x"39",
          3291 => x"33",
          3292 => x"2e",
          3293 => x"b3",
          3294 => x"88",
          3295 => x"fc",
          3296 => x"44",
          3297 => x"f8",
          3298 => x"84",
          3299 => x"a4",
          3300 => x"a8",
          3301 => x"a7",
          3302 => x"5d",
          3303 => x"2e",
          3304 => x"5d",
          3305 => x"70",
          3306 => x"07",
          3307 => x"60",
          3308 => x"5b",
          3309 => x"2e",
          3310 => x"a0",
          3311 => x"88",
          3312 => x"f4",
          3313 => x"3f",
          3314 => x"54",
          3315 => x"52",
          3316 => x"ac",
          3317 => x"84",
          3318 => x"39",
          3319 => x"80",
          3320 => x"84",
          3321 => x"cc",
          3322 => x"a8",
          3323 => x"f9",
          3324 => x"3d",
          3325 => x"53",
          3326 => x"51",
          3327 => x"82",
          3328 => x"80",
          3329 => x"64",
          3330 => x"cf",
          3331 => x"34",
          3332 => x"45",
          3333 => x"fc",
          3334 => x"84",
          3335 => x"94",
          3336 => x"a8",
          3337 => x"f9",
          3338 => x"70",
          3339 => x"82",
          3340 => x"ff",
          3341 => x"80",
          3342 => x"51",
          3343 => x"7a",
          3344 => x"5a",
          3345 => x"f8",
          3346 => x"7a",
          3347 => x"b5",
          3348 => x"11",
          3349 => x"05",
          3350 => x"3f",
          3351 => x"08",
          3352 => x"38",
          3353 => x"80",
          3354 => x"7a",
          3355 => x"05",
          3356 => x"39",
          3357 => x"51",
          3358 => x"ff",
          3359 => x"3d",
          3360 => x"53",
          3361 => x"51",
          3362 => x"82",
          3363 => x"80",
          3364 => x"38",
          3365 => x"f0",
          3366 => x"84",
          3367 => x"8d",
          3368 => x"a8",
          3369 => x"a6",
          3370 => x"02",
          3371 => x"22",
          3372 => x"05",
          3373 => x"42",
          3374 => x"f0",
          3375 => x"84",
          3376 => x"e9",
          3377 => x"a8",
          3378 => x"f7",
          3379 => x"70",
          3380 => x"82",
          3381 => x"ff",
          3382 => x"80",
          3383 => x"51",
          3384 => x"7a",
          3385 => x"5a",
          3386 => x"f7",
          3387 => x"9f",
          3388 => x"61",
          3389 => x"d6",
          3390 => x"fe",
          3391 => x"ff",
          3392 => x"c5",
          3393 => x"b5",
          3394 => x"2e",
          3395 => x"5a",
          3396 => x"05",
          3397 => x"82",
          3398 => x"79",
          3399 => x"39",
          3400 => x"51",
          3401 => x"ff",
          3402 => x"3d",
          3403 => x"53",
          3404 => x"51",
          3405 => x"82",
          3406 => x"80",
          3407 => x"38",
          3408 => x"f0",
          3409 => x"84",
          3410 => x"e1",
          3411 => x"a8",
          3412 => x"a0",
          3413 => x"71",
          3414 => x"84",
          3415 => x"3d",
          3416 => x"53",
          3417 => x"51",
          3418 => x"82",
          3419 => x"e5",
          3420 => x"39",
          3421 => x"54",
          3422 => x"b0",
          3423 => x"d8",
          3424 => x"52",
          3425 => x"f6",
          3426 => x"7a",
          3427 => x"ae",
          3428 => x"38",
          3429 => x"9b",
          3430 => x"fe",
          3431 => x"ff",
          3432 => x"c4",
          3433 => x"b5",
          3434 => x"2e",
          3435 => x"61",
          3436 => x"61",
          3437 => x"ff",
          3438 => x"a2",
          3439 => x"c5",
          3440 => x"39",
          3441 => x"80",
          3442 => x"84",
          3443 => x"e4",
          3444 => x"a8",
          3445 => x"f5",
          3446 => x"52",
          3447 => x"51",
          3448 => x"3f",
          3449 => x"04",
          3450 => x"80",
          3451 => x"84",
          3452 => x"c0",
          3453 => x"a8",
          3454 => x"f5",
          3455 => x"52",
          3456 => x"51",
          3457 => x"3f",
          3458 => x"2d",
          3459 => x"08",
          3460 => x"a3",
          3461 => x"a8",
          3462 => x"a2",
          3463 => x"a7",
          3464 => x"93",
          3465 => x"90",
          3466 => x"3f",
          3467 => x"3f",
          3468 => x"82",
          3469 => x"ce",
          3470 => x"5a",
          3471 => x"91",
          3472 => x"f3",
          3473 => x"7a",
          3474 => x"80",
          3475 => x"38",
          3476 => x"5a",
          3477 => x"81",
          3478 => x"3d",
          3479 => x"51",
          3480 => x"82",
          3481 => x"5d",
          3482 => x"82",
          3483 => x"7b",
          3484 => x"38",
          3485 => x"8c",
          3486 => x"39",
          3487 => x"b0",
          3488 => x"39",
          3489 => x"56",
          3490 => x"a3",
          3491 => x"53",
          3492 => x"52",
          3493 => x"b0",
          3494 => x"a9",
          3495 => x"39",
          3496 => x"52",
          3497 => x"b0",
          3498 => x"a9",
          3499 => x"39",
          3500 => x"a3",
          3501 => x"53",
          3502 => x"52",
          3503 => x"b0",
          3504 => x"a8",
          3505 => x"39",
          3506 => x"53",
          3507 => x"52",
          3508 => x"b0",
          3509 => x"a8",
          3510 => x"cc",
          3511 => x"b3",
          3512 => x"b5",
          3513 => x"56",
          3514 => x"54",
          3515 => x"53",
          3516 => x"52",
          3517 => x"b0",
          3518 => x"b9",
          3519 => x"a8",
          3520 => x"a8",
          3521 => x"30",
          3522 => x"80",
          3523 => x"5c",
          3524 => x"7b",
          3525 => x"38",
          3526 => x"7b",
          3527 => x"80",
          3528 => x"81",
          3529 => x"ff",
          3530 => x"7b",
          3531 => x"7e",
          3532 => x"81",
          3533 => x"79",
          3534 => x"ff",
          3535 => x"06",
          3536 => x"82",
          3537 => x"cc",
          3538 => x"eb",
          3539 => x"0d",
          3540 => x"b5",
          3541 => x"c0",
          3542 => x"08",
          3543 => x"84",
          3544 => x"51",
          3545 => x"82",
          3546 => x"90",
          3547 => x"55",
          3548 => x"80",
          3549 => x"e3",
          3550 => x"82",
          3551 => x"07",
          3552 => x"c0",
          3553 => x"08",
          3554 => x"84",
          3555 => x"51",
          3556 => x"82",
          3557 => x"90",
          3558 => x"55",
          3559 => x"80",
          3560 => x"e3",
          3561 => x"82",
          3562 => x"07",
          3563 => x"80",
          3564 => x"c0",
          3565 => x"8c",
          3566 => x"87",
          3567 => x"0c",
          3568 => x"51",
          3569 => x"80",
          3570 => x"80",
          3571 => x"83",
          3572 => x"99",
          3573 => x"5c",
          3574 => x"05",
          3575 => x"0c",
          3576 => x"93",
          3577 => x"a4",
          3578 => x"99",
          3579 => x"a4",
          3580 => x"3f",
          3581 => x"51",
          3582 => x"80",
          3583 => x"92",
          3584 => x"51",
          3585 => x"f0",
          3586 => x"04",
          3587 => x"80",
          3588 => x"71",
          3589 => x"87",
          3590 => x"b5",
          3591 => x"ff",
          3592 => x"ff",
          3593 => x"72",
          3594 => x"38",
          3595 => x"a8",
          3596 => x"0d",
          3597 => x"0d",
          3598 => x"54",
          3599 => x"52",
          3600 => x"2e",
          3601 => x"72",
          3602 => x"a0",
          3603 => x"06",
          3604 => x"13",
          3605 => x"72",
          3606 => x"a2",
          3607 => x"06",
          3608 => x"13",
          3609 => x"72",
          3610 => x"2e",
          3611 => x"9f",
          3612 => x"81",
          3613 => x"72",
          3614 => x"70",
          3615 => x"38",
          3616 => x"80",
          3617 => x"73",
          3618 => x"39",
          3619 => x"80",
          3620 => x"54",
          3621 => x"83",
          3622 => x"70",
          3623 => x"38",
          3624 => x"80",
          3625 => x"54",
          3626 => x"09",
          3627 => x"38",
          3628 => x"a2",
          3629 => x"70",
          3630 => x"07",
          3631 => x"70",
          3632 => x"38",
          3633 => x"81",
          3634 => x"71",
          3635 => x"51",
          3636 => x"a8",
          3637 => x"0d",
          3638 => x"0d",
          3639 => x"08",
          3640 => x"38",
          3641 => x"05",
          3642 => x"ff",
          3643 => x"82",
          3644 => x"85",
          3645 => x"83",
          3646 => x"72",
          3647 => x"0c",
          3648 => x"04",
          3649 => x"76",
          3650 => x"ff",
          3651 => x"81",
          3652 => x"26",
          3653 => x"83",
          3654 => x"05",
          3655 => x"70",
          3656 => x"8a",
          3657 => x"33",
          3658 => x"70",
          3659 => x"fe",
          3660 => x"33",
          3661 => x"70",
          3662 => x"f2",
          3663 => x"33",
          3664 => x"70",
          3665 => x"e6",
          3666 => x"22",
          3667 => x"74",
          3668 => x"80",
          3669 => x"13",
          3670 => x"52",
          3671 => x"26",
          3672 => x"81",
          3673 => x"98",
          3674 => x"22",
          3675 => x"bc",
          3676 => x"33",
          3677 => x"b8",
          3678 => x"33",
          3679 => x"b4",
          3680 => x"33",
          3681 => x"b0",
          3682 => x"33",
          3683 => x"ac",
          3684 => x"33",
          3685 => x"a8",
          3686 => x"c0",
          3687 => x"73",
          3688 => x"a0",
          3689 => x"87",
          3690 => x"0c",
          3691 => x"82",
          3692 => x"86",
          3693 => x"f3",
          3694 => x"5b",
          3695 => x"9c",
          3696 => x"0c",
          3697 => x"bc",
          3698 => x"7b",
          3699 => x"98",
          3700 => x"79",
          3701 => x"87",
          3702 => x"08",
          3703 => x"1c",
          3704 => x"98",
          3705 => x"79",
          3706 => x"87",
          3707 => x"08",
          3708 => x"1c",
          3709 => x"98",
          3710 => x"79",
          3711 => x"87",
          3712 => x"08",
          3713 => x"1c",
          3714 => x"98",
          3715 => x"79",
          3716 => x"80",
          3717 => x"83",
          3718 => x"59",
          3719 => x"ff",
          3720 => x"1b",
          3721 => x"1b",
          3722 => x"1b",
          3723 => x"1b",
          3724 => x"1b",
          3725 => x"83",
          3726 => x"52",
          3727 => x"51",
          3728 => x"3f",
          3729 => x"04",
          3730 => x"02",
          3731 => x"82",
          3732 => x"70",
          3733 => x"58",
          3734 => x"c0",
          3735 => x"75",
          3736 => x"38",
          3737 => x"94",
          3738 => x"70",
          3739 => x"81",
          3740 => x"52",
          3741 => x"8c",
          3742 => x"2a",
          3743 => x"51",
          3744 => x"38",
          3745 => x"70",
          3746 => x"51",
          3747 => x"8d",
          3748 => x"2a",
          3749 => x"51",
          3750 => x"be",
          3751 => x"ff",
          3752 => x"c0",
          3753 => x"70",
          3754 => x"38",
          3755 => x"90",
          3756 => x"0c",
          3757 => x"a8",
          3758 => x"0d",
          3759 => x"0d",
          3760 => x"33",
          3761 => x"9f",
          3762 => x"52",
          3763 => x"c8",
          3764 => x"0d",
          3765 => x"0d",
          3766 => x"33",
          3767 => x"2e",
          3768 => x"87",
          3769 => x"8d",
          3770 => x"82",
          3771 => x"70",
          3772 => x"58",
          3773 => x"94",
          3774 => x"80",
          3775 => x"87",
          3776 => x"53",
          3777 => x"96",
          3778 => x"06",
          3779 => x"72",
          3780 => x"38",
          3781 => x"70",
          3782 => x"53",
          3783 => x"74",
          3784 => x"81",
          3785 => x"72",
          3786 => x"38",
          3787 => x"70",
          3788 => x"53",
          3789 => x"38",
          3790 => x"06",
          3791 => x"94",
          3792 => x"80",
          3793 => x"87",
          3794 => x"54",
          3795 => x"80",
          3796 => x"a8",
          3797 => x"0d",
          3798 => x"0d",
          3799 => x"74",
          3800 => x"ff",
          3801 => x"57",
          3802 => x"80",
          3803 => x"81",
          3804 => x"15",
          3805 => x"33",
          3806 => x"06",
          3807 => x"58",
          3808 => x"84",
          3809 => x"2e",
          3810 => x"c0",
          3811 => x"70",
          3812 => x"2a",
          3813 => x"53",
          3814 => x"80",
          3815 => x"71",
          3816 => x"81",
          3817 => x"70",
          3818 => x"81",
          3819 => x"06",
          3820 => x"80",
          3821 => x"71",
          3822 => x"81",
          3823 => x"70",
          3824 => x"74",
          3825 => x"51",
          3826 => x"80",
          3827 => x"2e",
          3828 => x"c0",
          3829 => x"77",
          3830 => x"17",
          3831 => x"81",
          3832 => x"53",
          3833 => x"86",
          3834 => x"b5",
          3835 => x"3d",
          3836 => x"3d",
          3837 => x"c8",
          3838 => x"ff",
          3839 => x"87",
          3840 => x"51",
          3841 => x"86",
          3842 => x"94",
          3843 => x"08",
          3844 => x"70",
          3845 => x"51",
          3846 => x"2e",
          3847 => x"81",
          3848 => x"87",
          3849 => x"52",
          3850 => x"86",
          3851 => x"94",
          3852 => x"08",
          3853 => x"06",
          3854 => x"0c",
          3855 => x"0d",
          3856 => x"3f",
          3857 => x"08",
          3858 => x"82",
          3859 => x"04",
          3860 => x"82",
          3861 => x"70",
          3862 => x"52",
          3863 => x"94",
          3864 => x"80",
          3865 => x"87",
          3866 => x"52",
          3867 => x"82",
          3868 => x"06",
          3869 => x"ff",
          3870 => x"2e",
          3871 => x"81",
          3872 => x"87",
          3873 => x"52",
          3874 => x"86",
          3875 => x"94",
          3876 => x"08",
          3877 => x"70",
          3878 => x"53",
          3879 => x"b5",
          3880 => x"3d",
          3881 => x"3d",
          3882 => x"9e",
          3883 => x"9c",
          3884 => x"51",
          3885 => x"2e",
          3886 => x"87",
          3887 => x"08",
          3888 => x"0c",
          3889 => x"a8",
          3890 => x"d0",
          3891 => x"9e",
          3892 => x"b3",
          3893 => x"c0",
          3894 => x"82",
          3895 => x"87",
          3896 => x"08",
          3897 => x"0c",
          3898 => x"a0",
          3899 => x"e0",
          3900 => x"9e",
          3901 => x"b3",
          3902 => x"c0",
          3903 => x"82",
          3904 => x"87",
          3905 => x"08",
          3906 => x"0c",
          3907 => x"b8",
          3908 => x"f0",
          3909 => x"9e",
          3910 => x"b3",
          3911 => x"c0",
          3912 => x"82",
          3913 => x"87",
          3914 => x"08",
          3915 => x"0c",
          3916 => x"80",
          3917 => x"82",
          3918 => x"87",
          3919 => x"08",
          3920 => x"0c",
          3921 => x"88",
          3922 => x"88",
          3923 => x"9e",
          3924 => x"b4",
          3925 => x"0b",
          3926 => x"34",
          3927 => x"c0",
          3928 => x"70",
          3929 => x"06",
          3930 => x"70",
          3931 => x"38",
          3932 => x"82",
          3933 => x"80",
          3934 => x"9e",
          3935 => x"88",
          3936 => x"51",
          3937 => x"80",
          3938 => x"81",
          3939 => x"b4",
          3940 => x"0b",
          3941 => x"90",
          3942 => x"80",
          3943 => x"52",
          3944 => x"2e",
          3945 => x"52",
          3946 => x"93",
          3947 => x"87",
          3948 => x"08",
          3949 => x"80",
          3950 => x"52",
          3951 => x"83",
          3952 => x"71",
          3953 => x"34",
          3954 => x"c0",
          3955 => x"70",
          3956 => x"06",
          3957 => x"70",
          3958 => x"38",
          3959 => x"82",
          3960 => x"80",
          3961 => x"9e",
          3962 => x"90",
          3963 => x"51",
          3964 => x"80",
          3965 => x"81",
          3966 => x"b4",
          3967 => x"0b",
          3968 => x"90",
          3969 => x"80",
          3970 => x"52",
          3971 => x"2e",
          3972 => x"52",
          3973 => x"97",
          3974 => x"87",
          3975 => x"08",
          3976 => x"80",
          3977 => x"52",
          3978 => x"83",
          3979 => x"71",
          3980 => x"34",
          3981 => x"c0",
          3982 => x"70",
          3983 => x"06",
          3984 => x"70",
          3985 => x"38",
          3986 => x"82",
          3987 => x"80",
          3988 => x"9e",
          3989 => x"80",
          3990 => x"51",
          3991 => x"80",
          3992 => x"81",
          3993 => x"b4",
          3994 => x"0b",
          3995 => x"90",
          3996 => x"80",
          3997 => x"52",
          3998 => x"83",
          3999 => x"71",
          4000 => x"34",
          4001 => x"90",
          4002 => x"80",
          4003 => x"2a",
          4004 => x"70",
          4005 => x"34",
          4006 => x"c0",
          4007 => x"70",
          4008 => x"51",
          4009 => x"80",
          4010 => x"81",
          4011 => x"b4",
          4012 => x"c0",
          4013 => x"70",
          4014 => x"70",
          4015 => x"51",
          4016 => x"b4",
          4017 => x"0b",
          4018 => x"90",
          4019 => x"06",
          4020 => x"70",
          4021 => x"38",
          4022 => x"82",
          4023 => x"87",
          4024 => x"08",
          4025 => x"51",
          4026 => x"b4",
          4027 => x"3d",
          4028 => x"3d",
          4029 => x"e0",
          4030 => x"89",
          4031 => x"90",
          4032 => x"80",
          4033 => x"82",
          4034 => x"ff",
          4035 => x"82",
          4036 => x"ff",
          4037 => x"82",
          4038 => x"54",
          4039 => x"94",
          4040 => x"ec",
          4041 => x"f0",
          4042 => x"52",
          4043 => x"51",
          4044 => x"3f",
          4045 => x"33",
          4046 => x"2e",
          4047 => x"b3",
          4048 => x"b3",
          4049 => x"54",
          4050 => x"bc",
          4051 => x"88",
          4052 => x"94",
          4053 => x"80",
          4054 => x"82",
          4055 => x"82",
          4056 => x"11",
          4057 => x"a5",
          4058 => x"94",
          4059 => x"b4",
          4060 => x"73",
          4061 => x"38",
          4062 => x"08",
          4063 => x"08",
          4064 => x"82",
          4065 => x"ff",
          4066 => x"82",
          4067 => x"54",
          4068 => x"94",
          4069 => x"dc",
          4070 => x"e0",
          4071 => x"52",
          4072 => x"51",
          4073 => x"3f",
          4074 => x"33",
          4075 => x"2e",
          4076 => x"b4",
          4077 => x"82",
          4078 => x"ff",
          4079 => x"82",
          4080 => x"54",
          4081 => x"8e",
          4082 => x"a0",
          4083 => x"a6",
          4084 => x"94",
          4085 => x"b4",
          4086 => x"73",
          4087 => x"38",
          4088 => x"33",
          4089 => x"ec",
          4090 => x"ec",
          4091 => x"91",
          4092 => x"80",
          4093 => x"82",
          4094 => x"ff",
          4095 => x"82",
          4096 => x"54",
          4097 => x"89",
          4098 => x"a0",
          4099 => x"f5",
          4100 => x"98",
          4101 => x"80",
          4102 => x"82",
          4103 => x"ff",
          4104 => x"82",
          4105 => x"54",
          4106 => x"89",
          4107 => x"b8",
          4108 => x"d1",
          4109 => x"9a",
          4110 => x"80",
          4111 => x"82",
          4112 => x"ff",
          4113 => x"82",
          4114 => x"ff",
          4115 => x"82",
          4116 => x"52",
          4117 => x"51",
          4118 => x"3f",
          4119 => x"08",
          4120 => x"84",
          4121 => x"f0",
          4122 => x"fc",
          4123 => x"a8",
          4124 => x"92",
          4125 => x"a8",
          4126 => x"ba",
          4127 => x"b4",
          4128 => x"82",
          4129 => x"ff",
          4130 => x"82",
          4131 => x"56",
          4132 => x"52",
          4133 => x"8d",
          4134 => x"a8",
          4135 => x"c0",
          4136 => x"31",
          4137 => x"b5",
          4138 => x"82",
          4139 => x"ff",
          4140 => x"82",
          4141 => x"54",
          4142 => x"a9",
          4143 => x"88",
          4144 => x"84",
          4145 => x"51",
          4146 => x"82",
          4147 => x"bd",
          4148 => x"76",
          4149 => x"54",
          4150 => x"08",
          4151 => x"b0",
          4152 => x"f4",
          4153 => x"92",
          4154 => x"80",
          4155 => x"82",
          4156 => x"56",
          4157 => x"52",
          4158 => x"a9",
          4159 => x"a8",
          4160 => x"c0",
          4161 => x"31",
          4162 => x"b5",
          4163 => x"82",
          4164 => x"ff",
          4165 => x"82",
          4166 => x"ff",
          4167 => x"87",
          4168 => x"fe",
          4169 => x"92",
          4170 => x"05",
          4171 => x"26",
          4172 => x"84",
          4173 => x"90",
          4174 => x"08",
          4175 => x"88",
          4176 => x"82",
          4177 => x"97",
          4178 => x"98",
          4179 => x"82",
          4180 => x"8b",
          4181 => x"a4",
          4182 => x"82",
          4183 => x"ff",
          4184 => x"84",
          4185 => x"71",
          4186 => x"04",
          4187 => x"c0",
          4188 => x"04",
          4189 => x"08",
          4190 => x"84",
          4191 => x"3d",
          4192 => x"2b",
          4193 => x"79",
          4194 => x"98",
          4195 => x"13",
          4196 => x"51",
          4197 => x"51",
          4198 => x"82",
          4199 => x"33",
          4200 => x"74",
          4201 => x"82",
          4202 => x"08",
          4203 => x"05",
          4204 => x"71",
          4205 => x"52",
          4206 => x"09",
          4207 => x"38",
          4208 => x"82",
          4209 => x"85",
          4210 => x"fc",
          4211 => x"02",
          4212 => x"05",
          4213 => x"54",
          4214 => x"80",
          4215 => x"88",
          4216 => x"c3",
          4217 => x"ff",
          4218 => x"88",
          4219 => x"b7",
          4220 => x"ff",
          4221 => x"73",
          4222 => x"ff",
          4223 => x"39",
          4224 => x"b7",
          4225 => x"73",
          4226 => x"0d",
          4227 => x"0d",
          4228 => x"05",
          4229 => x"02",
          4230 => x"05",
          4231 => x"80",
          4232 => x"29",
          4233 => x"05",
          4234 => x"59",
          4235 => x"59",
          4236 => x"86",
          4237 => x"9a",
          4238 => x"b5",
          4239 => x"84",
          4240 => x"a8",
          4241 => x"70",
          4242 => x"5a",
          4243 => x"82",
          4244 => x"75",
          4245 => x"80",
          4246 => x"29",
          4247 => x"05",
          4248 => x"56",
          4249 => x"2e",
          4250 => x"53",
          4251 => x"51",
          4252 => x"82",
          4253 => x"81",
          4254 => x"82",
          4255 => x"74",
          4256 => x"55",
          4257 => x"87",
          4258 => x"82",
          4259 => x"77",
          4260 => x"38",
          4261 => x"08",
          4262 => x"2e",
          4263 => x"b4",
          4264 => x"74",
          4265 => x"3d",
          4266 => x"76",
          4267 => x"75",
          4268 => x"c1",
          4269 => x"fc",
          4270 => x"51",
          4271 => x"3f",
          4272 => x"08",
          4273 => x"9e",
          4274 => x"0d",
          4275 => x"0d",
          4276 => x"53",
          4277 => x"08",
          4278 => x"2e",
          4279 => x"51",
          4280 => x"80",
          4281 => x"14",
          4282 => x"54",
          4283 => x"e6",
          4284 => x"82",
          4285 => x"82",
          4286 => x"52",
          4287 => x"95",
          4288 => x"80",
          4289 => x"82",
          4290 => x"51",
          4291 => x"80",
          4292 => x"fc",
          4293 => x"0d",
          4294 => x"0d",
          4295 => x"52",
          4296 => x"08",
          4297 => x"eb",
          4298 => x"a8",
          4299 => x"38",
          4300 => x"08",
          4301 => x"52",
          4302 => x"52",
          4303 => x"b9",
          4304 => x"a8",
          4305 => x"b9",
          4306 => x"c0",
          4307 => x"b5",
          4308 => x"80",
          4309 => x"a8",
          4310 => x"38",
          4311 => x"08",
          4312 => x"17",
          4313 => x"74",
          4314 => x"76",
          4315 => x"82",
          4316 => x"57",
          4317 => x"3f",
          4318 => x"09",
          4319 => x"b0",
          4320 => x"0d",
          4321 => x"0d",
          4322 => x"ad",
          4323 => x"5a",
          4324 => x"58",
          4325 => x"b4",
          4326 => x"80",
          4327 => x"82",
          4328 => x"81",
          4329 => x"0b",
          4330 => x"08",
          4331 => x"f8",
          4332 => x"70",
          4333 => x"8a",
          4334 => x"b5",
          4335 => x"2e",
          4336 => x"51",
          4337 => x"3f",
          4338 => x"08",
          4339 => x"55",
          4340 => x"b5",
          4341 => x"8e",
          4342 => x"a8",
          4343 => x"70",
          4344 => x"80",
          4345 => x"09",
          4346 => x"72",
          4347 => x"51",
          4348 => x"77",
          4349 => x"73",
          4350 => x"82",
          4351 => x"8c",
          4352 => x"51",
          4353 => x"3f",
          4354 => x"08",
          4355 => x"38",
          4356 => x"51",
          4357 => x"3f",
          4358 => x"09",
          4359 => x"38",
          4360 => x"51",
          4361 => x"3f",
          4362 => x"be",
          4363 => x"3d",
          4364 => x"b5",
          4365 => x"34",
          4366 => x"82",
          4367 => x"a9",
          4368 => x"f6",
          4369 => x"7e",
          4370 => x"72",
          4371 => x"5a",
          4372 => x"2e",
          4373 => x"a2",
          4374 => x"78",
          4375 => x"76",
          4376 => x"81",
          4377 => x"70",
          4378 => x"58",
          4379 => x"2e",
          4380 => x"86",
          4381 => x"26",
          4382 => x"54",
          4383 => x"82",
          4384 => x"70",
          4385 => x"ff",
          4386 => x"82",
          4387 => x"53",
          4388 => x"08",
          4389 => x"3f",
          4390 => x"08",
          4391 => x"84",
          4392 => x"74",
          4393 => x"38",
          4394 => x"88",
          4395 => x"fc",
          4396 => x"39",
          4397 => x"8c",
          4398 => x"53",
          4399 => x"ff",
          4400 => x"82",
          4401 => x"80",
          4402 => x"ff",
          4403 => x"52",
          4404 => x"b1",
          4405 => x"a8",
          4406 => x"06",
          4407 => x"38",
          4408 => x"39",
          4409 => x"81",
          4410 => x"54",
          4411 => x"ff",
          4412 => x"54",
          4413 => x"a8",
          4414 => x"0d",
          4415 => x"0d",
          4416 => x"b2",
          4417 => x"3d",
          4418 => x"5a",
          4419 => x"3d",
          4420 => x"80",
          4421 => x"fc",
          4422 => x"73",
          4423 => x"73",
          4424 => x"33",
          4425 => x"83",
          4426 => x"76",
          4427 => x"bc",
          4428 => x"76",
          4429 => x"73",
          4430 => x"ad",
          4431 => x"97",
          4432 => x"b5",
          4433 => x"b4",
          4434 => x"b5",
          4435 => x"2e",
          4436 => x"93",
          4437 => x"82",
          4438 => x"51",
          4439 => x"3f",
          4440 => x"08",
          4441 => x"38",
          4442 => x"51",
          4443 => x"3f",
          4444 => x"82",
          4445 => x"5b",
          4446 => x"08",
          4447 => x"52",
          4448 => x"52",
          4449 => x"f1",
          4450 => x"a8",
          4451 => x"b5",
          4452 => x"2e",
          4453 => x"80",
          4454 => x"b5",
          4455 => x"ff",
          4456 => x"82",
          4457 => x"55",
          4458 => x"b5",
          4459 => x"a9",
          4460 => x"a8",
          4461 => x"70",
          4462 => x"80",
          4463 => x"53",
          4464 => x"06",
          4465 => x"f8",
          4466 => x"1b",
          4467 => x"06",
          4468 => x"7b",
          4469 => x"80",
          4470 => x"2e",
          4471 => x"ff",
          4472 => x"39",
          4473 => x"f8",
          4474 => x"38",
          4475 => x"08",
          4476 => x"38",
          4477 => x"8f",
          4478 => x"d4",
          4479 => x"a8",
          4480 => x"70",
          4481 => x"59",
          4482 => x"ee",
          4483 => x"ff",
          4484 => x"d4",
          4485 => x"2b",
          4486 => x"82",
          4487 => x"70",
          4488 => x"97",
          4489 => x"2c",
          4490 => x"29",
          4491 => x"05",
          4492 => x"70",
          4493 => x"51",
          4494 => x"51",
          4495 => x"81",
          4496 => x"2e",
          4497 => x"77",
          4498 => x"38",
          4499 => x"0a",
          4500 => x"0a",
          4501 => x"2c",
          4502 => x"75",
          4503 => x"38",
          4504 => x"52",
          4505 => x"96",
          4506 => x"a8",
          4507 => x"06",
          4508 => x"2e",
          4509 => x"82",
          4510 => x"81",
          4511 => x"74",
          4512 => x"29",
          4513 => x"05",
          4514 => x"70",
          4515 => x"56",
          4516 => x"95",
          4517 => x"76",
          4518 => x"77",
          4519 => x"3f",
          4520 => x"08",
          4521 => x"54",
          4522 => x"d3",
          4523 => x"75",
          4524 => x"ca",
          4525 => x"55",
          4526 => x"d4",
          4527 => x"2b",
          4528 => x"82",
          4529 => x"70",
          4530 => x"98",
          4531 => x"11",
          4532 => x"82",
          4533 => x"33",
          4534 => x"51",
          4535 => x"55",
          4536 => x"09",
          4537 => x"92",
          4538 => x"bc",
          4539 => x"0c",
          4540 => x"cc",
          4541 => x"0b",
          4542 => x"34",
          4543 => x"82",
          4544 => x"75",
          4545 => x"34",
          4546 => x"34",
          4547 => x"7e",
          4548 => x"26",
          4549 => x"73",
          4550 => x"95",
          4551 => x"73",
          4552 => x"cc",
          4553 => x"73",
          4554 => x"cb",
          4555 => x"d8",
          4556 => x"75",
          4557 => x"74",
          4558 => x"98",
          4559 => x"73",
          4560 => x"38",
          4561 => x"73",
          4562 => x"34",
          4563 => x"0a",
          4564 => x"0a",
          4565 => x"2c",
          4566 => x"33",
          4567 => x"df",
          4568 => x"dc",
          4569 => x"56",
          4570 => x"cc",
          4571 => x"1a",
          4572 => x"33",
          4573 => x"cc",
          4574 => x"73",
          4575 => x"38",
          4576 => x"73",
          4577 => x"34",
          4578 => x"33",
          4579 => x"0a",
          4580 => x"0a",
          4581 => x"2c",
          4582 => x"33",
          4583 => x"56",
          4584 => x"a3",
          4585 => x"70",
          4586 => x"ff",
          4587 => x"74",
          4588 => x"29",
          4589 => x"05",
          4590 => x"82",
          4591 => x"56",
          4592 => x"75",
          4593 => x"82",
          4594 => x"70",
          4595 => x"98",
          4596 => x"d8",
          4597 => x"56",
          4598 => x"25",
          4599 => x"88",
          4600 => x"c3",
          4601 => x"80",
          4602 => x"80",
          4603 => x"98",
          4604 => x"d8",
          4605 => x"55",
          4606 => x"e3",
          4607 => x"39",
          4608 => x"80",
          4609 => x"34",
          4610 => x"53",
          4611 => x"a2",
          4612 => x"b7",
          4613 => x"39",
          4614 => x"33",
          4615 => x"06",
          4616 => x"80",
          4617 => x"38",
          4618 => x"33",
          4619 => x"73",
          4620 => x"34",
          4621 => x"73",
          4622 => x"34",
          4623 => x"ad",
          4624 => x"cc",
          4625 => x"98",
          4626 => x"2c",
          4627 => x"33",
          4628 => x"57",
          4629 => x"a8",
          4630 => x"54",
          4631 => x"74",
          4632 => x"51",
          4633 => x"3f",
          4634 => x"0a",
          4635 => x"0a",
          4636 => x"2c",
          4637 => x"33",
          4638 => x"75",
          4639 => x"38",
          4640 => x"ad",
          4641 => x"cc",
          4642 => x"98",
          4643 => x"2c",
          4644 => x"33",
          4645 => x"57",
          4646 => x"fa",
          4647 => x"51",
          4648 => x"3f",
          4649 => x"0a",
          4650 => x"0a",
          4651 => x"2c",
          4652 => x"33",
          4653 => x"75",
          4654 => x"38",
          4655 => x"82",
          4656 => x"7a",
          4657 => x"74",
          4658 => x"ff",
          4659 => x"82",
          4660 => x"79",
          4661 => x"3f",
          4662 => x"08",
          4663 => x"54",
          4664 => x"82",
          4665 => x"54",
          4666 => x"8f",
          4667 => x"73",
          4668 => x"f2",
          4669 => x"39",
          4670 => x"80",
          4671 => x"dc",
          4672 => x"82",
          4673 => x"79",
          4674 => x"0c",
          4675 => x"04",
          4676 => x"33",
          4677 => x"2e",
          4678 => x"88",
          4679 => x"87",
          4680 => x"dc",
          4681 => x"54",
          4682 => x"dc",
          4683 => x"ff",
          4684 => x"39",
          4685 => x"33",
          4686 => x"33",
          4687 => x"75",
          4688 => x"38",
          4689 => x"73",
          4690 => x"34",
          4691 => x"70",
          4692 => x"81",
          4693 => x"51",
          4694 => x"25",
          4695 => x"1a",
          4696 => x"33",
          4697 => x"33",
          4698 => x"bb",
          4699 => x"80",
          4700 => x"80",
          4701 => x"98",
          4702 => x"d8",
          4703 => x"55",
          4704 => x"da",
          4705 => x"ff",
          4706 => x"82",
          4707 => x"70",
          4708 => x"98",
          4709 => x"d8",
          4710 => x"56",
          4711 => x"24",
          4712 => x"88",
          4713 => x"ff",
          4714 => x"80",
          4715 => x"80",
          4716 => x"98",
          4717 => x"d8",
          4718 => x"55",
          4719 => x"e3",
          4720 => x"39",
          4721 => x"33",
          4722 => x"06",
          4723 => x"33",
          4724 => x"74",
          4725 => x"9f",
          4726 => x"54",
          4727 => x"dc",
          4728 => x"70",
          4729 => x"ff",
          4730 => x"82",
          4731 => x"70",
          4732 => x"82",
          4733 => x"58",
          4734 => x"75",
          4735 => x"f7",
          4736 => x"cc",
          4737 => x"52",
          4738 => x"51",
          4739 => x"80",
          4740 => x"dc",
          4741 => x"82",
          4742 => x"f7",
          4743 => x"b0",
          4744 => x"f4",
          4745 => x"80",
          4746 => x"74",
          4747 => x"f7",
          4748 => x"a8",
          4749 => x"d8",
          4750 => x"a8",
          4751 => x"06",
          4752 => x"74",
          4753 => x"ff",
          4754 => x"93",
          4755 => x"39",
          4756 => x"82",
          4757 => x"fc",
          4758 => x"54",
          4759 => x"a7",
          4760 => x"ff",
          4761 => x"82",
          4762 => x"82",
          4763 => x"82",
          4764 => x"81",
          4765 => x"05",
          4766 => x"79",
          4767 => x"87",
          4768 => x"54",
          4769 => x"73",
          4770 => x"80",
          4771 => x"38",
          4772 => x"b2",
          4773 => x"39",
          4774 => x"09",
          4775 => x"38",
          4776 => x"08",
          4777 => x"2e",
          4778 => x"51",
          4779 => x"3f",
          4780 => x"08",
          4781 => x"34",
          4782 => x"08",
          4783 => x"81",
          4784 => x"52",
          4785 => x"b3",
          4786 => x"c3",
          4787 => x"29",
          4788 => x"05",
          4789 => x"54",
          4790 => x"ab",
          4791 => x"ff",
          4792 => x"82",
          4793 => x"82",
          4794 => x"82",
          4795 => x"81",
          4796 => x"05",
          4797 => x"79",
          4798 => x"8b",
          4799 => x"54",
          4800 => x"06",
          4801 => x"74",
          4802 => x"34",
          4803 => x"82",
          4804 => x"82",
          4805 => x"52",
          4806 => x"af",
          4807 => x"39",
          4808 => x"33",
          4809 => x"06",
          4810 => x"33",
          4811 => x"74",
          4812 => x"c3",
          4813 => x"54",
          4814 => x"dc",
          4815 => x"70",
          4816 => x"ff",
          4817 => x"f5",
          4818 => x"cc",
          4819 => x"73",
          4820 => x"a3",
          4821 => x"ff",
          4822 => x"82",
          4823 => x"ff",
          4824 => x"82",
          4825 => x"f5",
          4826 => x"3d",
          4827 => x"f4",
          4828 => x"a0",
          4829 => x"0b",
          4830 => x"23",
          4831 => x"80",
          4832 => x"f4",
          4833 => x"80",
          4834 => x"a0",
          4835 => x"58",
          4836 => x"81",
          4837 => x"15",
          4838 => x"a0",
          4839 => x"84",
          4840 => x"85",
          4841 => x"b5",
          4842 => x"77",
          4843 => x"76",
          4844 => x"82",
          4845 => x"82",
          4846 => x"ff",
          4847 => x"80",
          4848 => x"ff",
          4849 => x"88",
          4850 => x"55",
          4851 => x"17",
          4852 => x"17",
          4853 => x"9c",
          4854 => x"29",
          4855 => x"08",
          4856 => x"51",
          4857 => x"82",
          4858 => x"83",
          4859 => x"3d",
          4860 => x"3d",
          4861 => x"81",
          4862 => x"27",
          4863 => x"12",
          4864 => x"11",
          4865 => x"ff",
          4866 => x"51",
          4867 => x"a8",
          4868 => x"0d",
          4869 => x"0d",
          4870 => x"22",
          4871 => x"aa",
          4872 => x"05",
          4873 => x"08",
          4874 => x"71",
          4875 => x"2b",
          4876 => x"33",
          4877 => x"71",
          4878 => x"02",
          4879 => x"05",
          4880 => x"ff",
          4881 => x"70",
          4882 => x"51",
          4883 => x"5b",
          4884 => x"54",
          4885 => x"34",
          4886 => x"34",
          4887 => x"08",
          4888 => x"2a",
          4889 => x"82",
          4890 => x"83",
          4891 => x"b5",
          4892 => x"17",
          4893 => x"12",
          4894 => x"2b",
          4895 => x"2b",
          4896 => x"06",
          4897 => x"52",
          4898 => x"83",
          4899 => x"70",
          4900 => x"54",
          4901 => x"12",
          4902 => x"ff",
          4903 => x"83",
          4904 => x"b5",
          4905 => x"56",
          4906 => x"72",
          4907 => x"89",
          4908 => x"fb",
          4909 => x"b5",
          4910 => x"84",
          4911 => x"22",
          4912 => x"72",
          4913 => x"33",
          4914 => x"71",
          4915 => x"83",
          4916 => x"5b",
          4917 => x"52",
          4918 => x"12",
          4919 => x"33",
          4920 => x"07",
          4921 => x"54",
          4922 => x"70",
          4923 => x"73",
          4924 => x"82",
          4925 => x"70",
          4926 => x"33",
          4927 => x"71",
          4928 => x"83",
          4929 => x"59",
          4930 => x"05",
          4931 => x"87",
          4932 => x"88",
          4933 => x"88",
          4934 => x"56",
          4935 => x"13",
          4936 => x"13",
          4937 => x"a0",
          4938 => x"33",
          4939 => x"71",
          4940 => x"70",
          4941 => x"06",
          4942 => x"53",
          4943 => x"53",
          4944 => x"70",
          4945 => x"87",
          4946 => x"fa",
          4947 => x"a2",
          4948 => x"b5",
          4949 => x"83",
          4950 => x"70",
          4951 => x"33",
          4952 => x"07",
          4953 => x"15",
          4954 => x"12",
          4955 => x"2b",
          4956 => x"07",
          4957 => x"55",
          4958 => x"57",
          4959 => x"80",
          4960 => x"38",
          4961 => x"ab",
          4962 => x"a0",
          4963 => x"70",
          4964 => x"33",
          4965 => x"71",
          4966 => x"74",
          4967 => x"81",
          4968 => x"88",
          4969 => x"83",
          4970 => x"f8",
          4971 => x"54",
          4972 => x"58",
          4973 => x"74",
          4974 => x"52",
          4975 => x"34",
          4976 => x"34",
          4977 => x"08",
          4978 => x"33",
          4979 => x"71",
          4980 => x"83",
          4981 => x"59",
          4982 => x"05",
          4983 => x"12",
          4984 => x"2b",
          4985 => x"ff",
          4986 => x"88",
          4987 => x"52",
          4988 => x"74",
          4989 => x"15",
          4990 => x"0d",
          4991 => x"0d",
          4992 => x"08",
          4993 => x"9e",
          4994 => x"83",
          4995 => x"82",
          4996 => x"12",
          4997 => x"2b",
          4998 => x"07",
          4999 => x"52",
          5000 => x"05",
          5001 => x"13",
          5002 => x"2b",
          5003 => x"05",
          5004 => x"71",
          5005 => x"2a",
          5006 => x"53",
          5007 => x"34",
          5008 => x"34",
          5009 => x"08",
          5010 => x"33",
          5011 => x"71",
          5012 => x"83",
          5013 => x"59",
          5014 => x"05",
          5015 => x"83",
          5016 => x"88",
          5017 => x"88",
          5018 => x"56",
          5019 => x"13",
          5020 => x"13",
          5021 => x"a0",
          5022 => x"11",
          5023 => x"33",
          5024 => x"07",
          5025 => x"0c",
          5026 => x"3d",
          5027 => x"3d",
          5028 => x"b5",
          5029 => x"83",
          5030 => x"ff",
          5031 => x"53",
          5032 => x"a7",
          5033 => x"a0",
          5034 => x"2b",
          5035 => x"11",
          5036 => x"33",
          5037 => x"71",
          5038 => x"75",
          5039 => x"81",
          5040 => x"98",
          5041 => x"2b",
          5042 => x"40",
          5043 => x"58",
          5044 => x"72",
          5045 => x"38",
          5046 => x"52",
          5047 => x"9d",
          5048 => x"39",
          5049 => x"85",
          5050 => x"8b",
          5051 => x"2b",
          5052 => x"79",
          5053 => x"51",
          5054 => x"76",
          5055 => x"75",
          5056 => x"56",
          5057 => x"34",
          5058 => x"08",
          5059 => x"12",
          5060 => x"33",
          5061 => x"07",
          5062 => x"54",
          5063 => x"53",
          5064 => x"34",
          5065 => x"34",
          5066 => x"08",
          5067 => x"0b",
          5068 => x"80",
          5069 => x"34",
          5070 => x"08",
          5071 => x"14",
          5072 => x"14",
          5073 => x"a0",
          5074 => x"33",
          5075 => x"71",
          5076 => x"70",
          5077 => x"07",
          5078 => x"53",
          5079 => x"54",
          5080 => x"72",
          5081 => x"8b",
          5082 => x"ff",
          5083 => x"52",
          5084 => x"08",
          5085 => x"f2",
          5086 => x"2e",
          5087 => x"51",
          5088 => x"83",
          5089 => x"f5",
          5090 => x"7e",
          5091 => x"e2",
          5092 => x"a8",
          5093 => x"ff",
          5094 => x"a0",
          5095 => x"33",
          5096 => x"71",
          5097 => x"70",
          5098 => x"58",
          5099 => x"ff",
          5100 => x"2e",
          5101 => x"75",
          5102 => x"70",
          5103 => x"33",
          5104 => x"07",
          5105 => x"ff",
          5106 => x"70",
          5107 => x"06",
          5108 => x"52",
          5109 => x"59",
          5110 => x"27",
          5111 => x"80",
          5112 => x"75",
          5113 => x"84",
          5114 => x"16",
          5115 => x"2b",
          5116 => x"75",
          5117 => x"81",
          5118 => x"85",
          5119 => x"59",
          5120 => x"83",
          5121 => x"a0",
          5122 => x"33",
          5123 => x"71",
          5124 => x"70",
          5125 => x"06",
          5126 => x"56",
          5127 => x"75",
          5128 => x"81",
          5129 => x"79",
          5130 => x"cc",
          5131 => x"74",
          5132 => x"c4",
          5133 => x"2e",
          5134 => x"89",
          5135 => x"f8",
          5136 => x"ac",
          5137 => x"80",
          5138 => x"75",
          5139 => x"3f",
          5140 => x"08",
          5141 => x"11",
          5142 => x"33",
          5143 => x"71",
          5144 => x"53",
          5145 => x"74",
          5146 => x"70",
          5147 => x"06",
          5148 => x"5c",
          5149 => x"78",
          5150 => x"76",
          5151 => x"57",
          5152 => x"34",
          5153 => x"08",
          5154 => x"71",
          5155 => x"86",
          5156 => x"12",
          5157 => x"2b",
          5158 => x"2a",
          5159 => x"53",
          5160 => x"73",
          5161 => x"75",
          5162 => x"82",
          5163 => x"70",
          5164 => x"33",
          5165 => x"71",
          5166 => x"83",
          5167 => x"5d",
          5168 => x"05",
          5169 => x"15",
          5170 => x"15",
          5171 => x"a0",
          5172 => x"71",
          5173 => x"33",
          5174 => x"71",
          5175 => x"70",
          5176 => x"5a",
          5177 => x"54",
          5178 => x"34",
          5179 => x"34",
          5180 => x"08",
          5181 => x"54",
          5182 => x"a8",
          5183 => x"0d",
          5184 => x"0d",
          5185 => x"b5",
          5186 => x"38",
          5187 => x"71",
          5188 => x"2e",
          5189 => x"51",
          5190 => x"82",
          5191 => x"53",
          5192 => x"a8",
          5193 => x"0d",
          5194 => x"0d",
          5195 => x"5c",
          5196 => x"40",
          5197 => x"08",
          5198 => x"81",
          5199 => x"f4",
          5200 => x"8e",
          5201 => x"ff",
          5202 => x"b5",
          5203 => x"83",
          5204 => x"8b",
          5205 => x"fc",
          5206 => x"54",
          5207 => x"7e",
          5208 => x"3f",
          5209 => x"08",
          5210 => x"06",
          5211 => x"08",
          5212 => x"83",
          5213 => x"ff",
          5214 => x"83",
          5215 => x"70",
          5216 => x"33",
          5217 => x"07",
          5218 => x"70",
          5219 => x"06",
          5220 => x"fc",
          5221 => x"29",
          5222 => x"81",
          5223 => x"88",
          5224 => x"90",
          5225 => x"4e",
          5226 => x"52",
          5227 => x"41",
          5228 => x"5b",
          5229 => x"8f",
          5230 => x"ff",
          5231 => x"31",
          5232 => x"ff",
          5233 => x"82",
          5234 => x"17",
          5235 => x"2b",
          5236 => x"29",
          5237 => x"81",
          5238 => x"98",
          5239 => x"2b",
          5240 => x"45",
          5241 => x"73",
          5242 => x"38",
          5243 => x"70",
          5244 => x"06",
          5245 => x"7b",
          5246 => x"38",
          5247 => x"73",
          5248 => x"81",
          5249 => x"78",
          5250 => x"3f",
          5251 => x"ff",
          5252 => x"e5",
          5253 => x"38",
          5254 => x"89",
          5255 => x"f6",
          5256 => x"a5",
          5257 => x"55",
          5258 => x"80",
          5259 => x"1d",
          5260 => x"83",
          5261 => x"88",
          5262 => x"57",
          5263 => x"3f",
          5264 => x"51",
          5265 => x"82",
          5266 => x"83",
          5267 => x"7e",
          5268 => x"70",
          5269 => x"b5",
          5270 => x"84",
          5271 => x"59",
          5272 => x"3f",
          5273 => x"08",
          5274 => x"75",
          5275 => x"06",
          5276 => x"85",
          5277 => x"54",
          5278 => x"80",
          5279 => x"51",
          5280 => x"82",
          5281 => x"1d",
          5282 => x"83",
          5283 => x"88",
          5284 => x"43",
          5285 => x"3f",
          5286 => x"51",
          5287 => x"82",
          5288 => x"83",
          5289 => x"7e",
          5290 => x"70",
          5291 => x"b5",
          5292 => x"84",
          5293 => x"59",
          5294 => x"3f",
          5295 => x"08",
          5296 => x"60",
          5297 => x"55",
          5298 => x"ff",
          5299 => x"a9",
          5300 => x"52",
          5301 => x"3f",
          5302 => x"08",
          5303 => x"a8",
          5304 => x"93",
          5305 => x"73",
          5306 => x"a8",
          5307 => x"a3",
          5308 => x"51",
          5309 => x"7a",
          5310 => x"27",
          5311 => x"53",
          5312 => x"51",
          5313 => x"7a",
          5314 => x"82",
          5315 => x"05",
          5316 => x"f6",
          5317 => x"54",
          5318 => x"a8",
          5319 => x"0d",
          5320 => x"0d",
          5321 => x"70",
          5322 => x"d5",
          5323 => x"a8",
          5324 => x"b5",
          5325 => x"2e",
          5326 => x"53",
          5327 => x"b5",
          5328 => x"ff",
          5329 => x"74",
          5330 => x"0c",
          5331 => x"04",
          5332 => x"02",
          5333 => x"51",
          5334 => x"72",
          5335 => x"82",
          5336 => x"33",
          5337 => x"b5",
          5338 => x"3d",
          5339 => x"3d",
          5340 => x"05",
          5341 => x"05",
          5342 => x"56",
          5343 => x"72",
          5344 => x"e0",
          5345 => x"2b",
          5346 => x"8c",
          5347 => x"88",
          5348 => x"2e",
          5349 => x"88",
          5350 => x"0c",
          5351 => x"8c",
          5352 => x"71",
          5353 => x"87",
          5354 => x"0c",
          5355 => x"08",
          5356 => x"51",
          5357 => x"2e",
          5358 => x"c0",
          5359 => x"51",
          5360 => x"71",
          5361 => x"80",
          5362 => x"92",
          5363 => x"98",
          5364 => x"70",
          5365 => x"38",
          5366 => x"a4",
          5367 => x"b5",
          5368 => x"51",
          5369 => x"a8",
          5370 => x"0d",
          5371 => x"0d",
          5372 => x"02",
          5373 => x"05",
          5374 => x"58",
          5375 => x"52",
          5376 => x"3f",
          5377 => x"08",
          5378 => x"54",
          5379 => x"be",
          5380 => x"75",
          5381 => x"c0",
          5382 => x"87",
          5383 => x"12",
          5384 => x"84",
          5385 => x"40",
          5386 => x"85",
          5387 => x"98",
          5388 => x"7d",
          5389 => x"0c",
          5390 => x"85",
          5391 => x"06",
          5392 => x"71",
          5393 => x"38",
          5394 => x"71",
          5395 => x"05",
          5396 => x"19",
          5397 => x"a2",
          5398 => x"71",
          5399 => x"38",
          5400 => x"83",
          5401 => x"38",
          5402 => x"8a",
          5403 => x"98",
          5404 => x"71",
          5405 => x"c0",
          5406 => x"52",
          5407 => x"87",
          5408 => x"80",
          5409 => x"81",
          5410 => x"c0",
          5411 => x"53",
          5412 => x"82",
          5413 => x"71",
          5414 => x"1a",
          5415 => x"84",
          5416 => x"19",
          5417 => x"06",
          5418 => x"79",
          5419 => x"38",
          5420 => x"80",
          5421 => x"87",
          5422 => x"26",
          5423 => x"73",
          5424 => x"06",
          5425 => x"2e",
          5426 => x"52",
          5427 => x"82",
          5428 => x"8f",
          5429 => x"f3",
          5430 => x"62",
          5431 => x"05",
          5432 => x"57",
          5433 => x"83",
          5434 => x"52",
          5435 => x"3f",
          5436 => x"08",
          5437 => x"54",
          5438 => x"2e",
          5439 => x"81",
          5440 => x"74",
          5441 => x"c0",
          5442 => x"87",
          5443 => x"12",
          5444 => x"84",
          5445 => x"5f",
          5446 => x"0b",
          5447 => x"8c",
          5448 => x"0c",
          5449 => x"80",
          5450 => x"70",
          5451 => x"81",
          5452 => x"54",
          5453 => x"8c",
          5454 => x"81",
          5455 => x"7c",
          5456 => x"58",
          5457 => x"70",
          5458 => x"52",
          5459 => x"8a",
          5460 => x"98",
          5461 => x"71",
          5462 => x"c0",
          5463 => x"52",
          5464 => x"87",
          5465 => x"80",
          5466 => x"81",
          5467 => x"c0",
          5468 => x"53",
          5469 => x"82",
          5470 => x"71",
          5471 => x"19",
          5472 => x"81",
          5473 => x"ff",
          5474 => x"19",
          5475 => x"78",
          5476 => x"38",
          5477 => x"80",
          5478 => x"87",
          5479 => x"26",
          5480 => x"73",
          5481 => x"06",
          5482 => x"2e",
          5483 => x"52",
          5484 => x"82",
          5485 => x"8f",
          5486 => x"fa",
          5487 => x"02",
          5488 => x"05",
          5489 => x"05",
          5490 => x"71",
          5491 => x"57",
          5492 => x"82",
          5493 => x"81",
          5494 => x"54",
          5495 => x"38",
          5496 => x"c0",
          5497 => x"81",
          5498 => x"2e",
          5499 => x"71",
          5500 => x"38",
          5501 => x"87",
          5502 => x"11",
          5503 => x"80",
          5504 => x"80",
          5505 => x"83",
          5506 => x"38",
          5507 => x"72",
          5508 => x"2a",
          5509 => x"51",
          5510 => x"80",
          5511 => x"87",
          5512 => x"08",
          5513 => x"38",
          5514 => x"8c",
          5515 => x"96",
          5516 => x"0c",
          5517 => x"8c",
          5518 => x"08",
          5519 => x"51",
          5520 => x"38",
          5521 => x"56",
          5522 => x"80",
          5523 => x"85",
          5524 => x"77",
          5525 => x"83",
          5526 => x"75",
          5527 => x"b5",
          5528 => x"3d",
          5529 => x"3d",
          5530 => x"11",
          5531 => x"71",
          5532 => x"82",
          5533 => x"53",
          5534 => x"0d",
          5535 => x"0d",
          5536 => x"33",
          5537 => x"71",
          5538 => x"88",
          5539 => x"14",
          5540 => x"07",
          5541 => x"33",
          5542 => x"b5",
          5543 => x"53",
          5544 => x"52",
          5545 => x"04",
          5546 => x"73",
          5547 => x"92",
          5548 => x"52",
          5549 => x"81",
          5550 => x"70",
          5551 => x"70",
          5552 => x"3d",
          5553 => x"3d",
          5554 => x"52",
          5555 => x"70",
          5556 => x"34",
          5557 => x"51",
          5558 => x"81",
          5559 => x"70",
          5560 => x"70",
          5561 => x"05",
          5562 => x"88",
          5563 => x"72",
          5564 => x"0d",
          5565 => x"0d",
          5566 => x"54",
          5567 => x"80",
          5568 => x"71",
          5569 => x"53",
          5570 => x"81",
          5571 => x"ff",
          5572 => x"39",
          5573 => x"04",
          5574 => x"75",
          5575 => x"52",
          5576 => x"70",
          5577 => x"34",
          5578 => x"70",
          5579 => x"3d",
          5580 => x"3d",
          5581 => x"79",
          5582 => x"74",
          5583 => x"56",
          5584 => x"81",
          5585 => x"71",
          5586 => x"16",
          5587 => x"52",
          5588 => x"86",
          5589 => x"2e",
          5590 => x"82",
          5591 => x"86",
          5592 => x"fe",
          5593 => x"76",
          5594 => x"39",
          5595 => x"8a",
          5596 => x"51",
          5597 => x"71",
          5598 => x"33",
          5599 => x"0c",
          5600 => x"04",
          5601 => x"b5",
          5602 => x"80",
          5603 => x"a8",
          5604 => x"3d",
          5605 => x"80",
          5606 => x"33",
          5607 => x"7a",
          5608 => x"38",
          5609 => x"16",
          5610 => x"16",
          5611 => x"17",
          5612 => x"fa",
          5613 => x"b5",
          5614 => x"2e",
          5615 => x"b7",
          5616 => x"a8",
          5617 => x"34",
          5618 => x"70",
          5619 => x"31",
          5620 => x"59",
          5621 => x"77",
          5622 => x"82",
          5623 => x"74",
          5624 => x"81",
          5625 => x"81",
          5626 => x"53",
          5627 => x"16",
          5628 => x"e3",
          5629 => x"81",
          5630 => x"b5",
          5631 => x"3d",
          5632 => x"3d",
          5633 => x"56",
          5634 => x"74",
          5635 => x"2e",
          5636 => x"51",
          5637 => x"82",
          5638 => x"57",
          5639 => x"08",
          5640 => x"54",
          5641 => x"16",
          5642 => x"33",
          5643 => x"3f",
          5644 => x"08",
          5645 => x"38",
          5646 => x"57",
          5647 => x"0c",
          5648 => x"a8",
          5649 => x"0d",
          5650 => x"0d",
          5651 => x"57",
          5652 => x"82",
          5653 => x"58",
          5654 => x"08",
          5655 => x"76",
          5656 => x"83",
          5657 => x"06",
          5658 => x"84",
          5659 => x"78",
          5660 => x"81",
          5661 => x"38",
          5662 => x"82",
          5663 => x"52",
          5664 => x"52",
          5665 => x"3f",
          5666 => x"52",
          5667 => x"51",
          5668 => x"84",
          5669 => x"d2",
          5670 => x"fc",
          5671 => x"8a",
          5672 => x"52",
          5673 => x"51",
          5674 => x"90",
          5675 => x"84",
          5676 => x"fc",
          5677 => x"17",
          5678 => x"a0",
          5679 => x"86",
          5680 => x"08",
          5681 => x"b0",
          5682 => x"55",
          5683 => x"81",
          5684 => x"f8",
          5685 => x"84",
          5686 => x"53",
          5687 => x"17",
          5688 => x"d7",
          5689 => x"a8",
          5690 => x"83",
          5691 => x"77",
          5692 => x"0c",
          5693 => x"04",
          5694 => x"77",
          5695 => x"12",
          5696 => x"55",
          5697 => x"56",
          5698 => x"8d",
          5699 => x"22",
          5700 => x"ac",
          5701 => x"57",
          5702 => x"b5",
          5703 => x"3d",
          5704 => x"3d",
          5705 => x"70",
          5706 => x"57",
          5707 => x"81",
          5708 => x"98",
          5709 => x"81",
          5710 => x"74",
          5711 => x"72",
          5712 => x"f5",
          5713 => x"24",
          5714 => x"81",
          5715 => x"81",
          5716 => x"83",
          5717 => x"38",
          5718 => x"76",
          5719 => x"70",
          5720 => x"16",
          5721 => x"74",
          5722 => x"96",
          5723 => x"a8",
          5724 => x"38",
          5725 => x"06",
          5726 => x"33",
          5727 => x"89",
          5728 => x"08",
          5729 => x"54",
          5730 => x"fc",
          5731 => x"b5",
          5732 => x"fe",
          5733 => x"ff",
          5734 => x"11",
          5735 => x"2b",
          5736 => x"81",
          5737 => x"2a",
          5738 => x"51",
          5739 => x"e2",
          5740 => x"ff",
          5741 => x"da",
          5742 => x"2a",
          5743 => x"05",
          5744 => x"fc",
          5745 => x"b5",
          5746 => x"c6",
          5747 => x"83",
          5748 => x"05",
          5749 => x"f9",
          5750 => x"b5",
          5751 => x"ff",
          5752 => x"ae",
          5753 => x"2a",
          5754 => x"05",
          5755 => x"fc",
          5756 => x"b5",
          5757 => x"38",
          5758 => x"83",
          5759 => x"05",
          5760 => x"f8",
          5761 => x"b5",
          5762 => x"0a",
          5763 => x"39",
          5764 => x"82",
          5765 => x"89",
          5766 => x"f8",
          5767 => x"7c",
          5768 => x"56",
          5769 => x"77",
          5770 => x"38",
          5771 => x"08",
          5772 => x"38",
          5773 => x"72",
          5774 => x"9d",
          5775 => x"24",
          5776 => x"81",
          5777 => x"82",
          5778 => x"83",
          5779 => x"38",
          5780 => x"76",
          5781 => x"70",
          5782 => x"18",
          5783 => x"76",
          5784 => x"9e",
          5785 => x"a8",
          5786 => x"b5",
          5787 => x"d9",
          5788 => x"ff",
          5789 => x"05",
          5790 => x"81",
          5791 => x"54",
          5792 => x"80",
          5793 => x"77",
          5794 => x"f0",
          5795 => x"8f",
          5796 => x"51",
          5797 => x"34",
          5798 => x"17",
          5799 => x"2a",
          5800 => x"05",
          5801 => x"fa",
          5802 => x"b5",
          5803 => x"82",
          5804 => x"81",
          5805 => x"83",
          5806 => x"b4",
          5807 => x"2a",
          5808 => x"8f",
          5809 => x"2a",
          5810 => x"f0",
          5811 => x"06",
          5812 => x"72",
          5813 => x"ec",
          5814 => x"2a",
          5815 => x"05",
          5816 => x"fa",
          5817 => x"b5",
          5818 => x"82",
          5819 => x"80",
          5820 => x"83",
          5821 => x"52",
          5822 => x"fe",
          5823 => x"b4",
          5824 => x"a4",
          5825 => x"76",
          5826 => x"17",
          5827 => x"75",
          5828 => x"3f",
          5829 => x"08",
          5830 => x"a8",
          5831 => x"77",
          5832 => x"77",
          5833 => x"fc",
          5834 => x"b4",
          5835 => x"51",
          5836 => x"c9",
          5837 => x"a8",
          5838 => x"06",
          5839 => x"72",
          5840 => x"3f",
          5841 => x"17",
          5842 => x"b5",
          5843 => x"3d",
          5844 => x"3d",
          5845 => x"7e",
          5846 => x"56",
          5847 => x"75",
          5848 => x"74",
          5849 => x"27",
          5850 => x"80",
          5851 => x"ff",
          5852 => x"75",
          5853 => x"3f",
          5854 => x"08",
          5855 => x"a8",
          5856 => x"38",
          5857 => x"54",
          5858 => x"81",
          5859 => x"39",
          5860 => x"08",
          5861 => x"39",
          5862 => x"51",
          5863 => x"82",
          5864 => x"58",
          5865 => x"08",
          5866 => x"c7",
          5867 => x"a8",
          5868 => x"d2",
          5869 => x"a8",
          5870 => x"cf",
          5871 => x"74",
          5872 => x"fc",
          5873 => x"b5",
          5874 => x"38",
          5875 => x"fe",
          5876 => x"08",
          5877 => x"74",
          5878 => x"38",
          5879 => x"17",
          5880 => x"33",
          5881 => x"73",
          5882 => x"77",
          5883 => x"26",
          5884 => x"80",
          5885 => x"b5",
          5886 => x"3d",
          5887 => x"3d",
          5888 => x"71",
          5889 => x"5b",
          5890 => x"8c",
          5891 => x"77",
          5892 => x"38",
          5893 => x"78",
          5894 => x"81",
          5895 => x"79",
          5896 => x"f9",
          5897 => x"55",
          5898 => x"a8",
          5899 => x"e0",
          5900 => x"a8",
          5901 => x"b5",
          5902 => x"2e",
          5903 => x"98",
          5904 => x"b5",
          5905 => x"82",
          5906 => x"58",
          5907 => x"70",
          5908 => x"80",
          5909 => x"38",
          5910 => x"09",
          5911 => x"e2",
          5912 => x"56",
          5913 => x"76",
          5914 => x"82",
          5915 => x"7a",
          5916 => x"3f",
          5917 => x"b5",
          5918 => x"2e",
          5919 => x"86",
          5920 => x"a8",
          5921 => x"b5",
          5922 => x"70",
          5923 => x"07",
          5924 => x"7c",
          5925 => x"a8",
          5926 => x"51",
          5927 => x"81",
          5928 => x"b5",
          5929 => x"2e",
          5930 => x"17",
          5931 => x"74",
          5932 => x"73",
          5933 => x"27",
          5934 => x"58",
          5935 => x"80",
          5936 => x"56",
          5937 => x"98",
          5938 => x"26",
          5939 => x"56",
          5940 => x"81",
          5941 => x"52",
          5942 => x"c6",
          5943 => x"a8",
          5944 => x"b8",
          5945 => x"82",
          5946 => x"81",
          5947 => x"06",
          5948 => x"b5",
          5949 => x"82",
          5950 => x"09",
          5951 => x"72",
          5952 => x"70",
          5953 => x"51",
          5954 => x"80",
          5955 => x"78",
          5956 => x"06",
          5957 => x"73",
          5958 => x"39",
          5959 => x"52",
          5960 => x"f7",
          5961 => x"a8",
          5962 => x"a8",
          5963 => x"82",
          5964 => x"07",
          5965 => x"55",
          5966 => x"2e",
          5967 => x"80",
          5968 => x"75",
          5969 => x"76",
          5970 => x"3f",
          5971 => x"08",
          5972 => x"38",
          5973 => x"0c",
          5974 => x"fe",
          5975 => x"08",
          5976 => x"74",
          5977 => x"ff",
          5978 => x"0c",
          5979 => x"81",
          5980 => x"84",
          5981 => x"39",
          5982 => x"81",
          5983 => x"8c",
          5984 => x"8c",
          5985 => x"a8",
          5986 => x"39",
          5987 => x"55",
          5988 => x"a8",
          5989 => x"0d",
          5990 => x"0d",
          5991 => x"55",
          5992 => x"82",
          5993 => x"58",
          5994 => x"b5",
          5995 => x"d8",
          5996 => x"74",
          5997 => x"3f",
          5998 => x"08",
          5999 => x"08",
          6000 => x"59",
          6001 => x"77",
          6002 => x"70",
          6003 => x"c8",
          6004 => x"84",
          6005 => x"56",
          6006 => x"58",
          6007 => x"97",
          6008 => x"75",
          6009 => x"52",
          6010 => x"51",
          6011 => x"82",
          6012 => x"80",
          6013 => x"8a",
          6014 => x"32",
          6015 => x"72",
          6016 => x"2a",
          6017 => x"56",
          6018 => x"a8",
          6019 => x"0d",
          6020 => x"0d",
          6021 => x"08",
          6022 => x"74",
          6023 => x"26",
          6024 => x"74",
          6025 => x"72",
          6026 => x"74",
          6027 => x"88",
          6028 => x"73",
          6029 => x"33",
          6030 => x"27",
          6031 => x"16",
          6032 => x"9b",
          6033 => x"2a",
          6034 => x"88",
          6035 => x"58",
          6036 => x"80",
          6037 => x"16",
          6038 => x"0c",
          6039 => x"8a",
          6040 => x"89",
          6041 => x"72",
          6042 => x"38",
          6043 => x"51",
          6044 => x"82",
          6045 => x"54",
          6046 => x"08",
          6047 => x"38",
          6048 => x"b5",
          6049 => x"8b",
          6050 => x"08",
          6051 => x"08",
          6052 => x"82",
          6053 => x"74",
          6054 => x"cb",
          6055 => x"75",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"73",
          6059 => x"98",
          6060 => x"82",
          6061 => x"2e",
          6062 => x"39",
          6063 => x"39",
          6064 => x"13",
          6065 => x"74",
          6066 => x"16",
          6067 => x"18",
          6068 => x"77",
          6069 => x"0c",
          6070 => x"04",
          6071 => x"7a",
          6072 => x"12",
          6073 => x"59",
          6074 => x"80",
          6075 => x"86",
          6076 => x"98",
          6077 => x"14",
          6078 => x"55",
          6079 => x"81",
          6080 => x"83",
          6081 => x"77",
          6082 => x"81",
          6083 => x"0c",
          6084 => x"55",
          6085 => x"76",
          6086 => x"17",
          6087 => x"74",
          6088 => x"9b",
          6089 => x"39",
          6090 => x"ff",
          6091 => x"2a",
          6092 => x"81",
          6093 => x"52",
          6094 => x"e6",
          6095 => x"a8",
          6096 => x"55",
          6097 => x"b5",
          6098 => x"80",
          6099 => x"55",
          6100 => x"08",
          6101 => x"f4",
          6102 => x"08",
          6103 => x"08",
          6104 => x"38",
          6105 => x"77",
          6106 => x"84",
          6107 => x"39",
          6108 => x"52",
          6109 => x"86",
          6110 => x"a8",
          6111 => x"55",
          6112 => x"08",
          6113 => x"c4",
          6114 => x"82",
          6115 => x"81",
          6116 => x"81",
          6117 => x"a8",
          6118 => x"b0",
          6119 => x"a8",
          6120 => x"51",
          6121 => x"82",
          6122 => x"a0",
          6123 => x"15",
          6124 => x"75",
          6125 => x"3f",
          6126 => x"08",
          6127 => x"76",
          6128 => x"77",
          6129 => x"9c",
          6130 => x"55",
          6131 => x"a8",
          6132 => x"0d",
          6133 => x"0d",
          6134 => x"08",
          6135 => x"80",
          6136 => x"fc",
          6137 => x"b5",
          6138 => x"82",
          6139 => x"80",
          6140 => x"b5",
          6141 => x"98",
          6142 => x"78",
          6143 => x"3f",
          6144 => x"08",
          6145 => x"a8",
          6146 => x"38",
          6147 => x"08",
          6148 => x"70",
          6149 => x"58",
          6150 => x"2e",
          6151 => x"83",
          6152 => x"82",
          6153 => x"55",
          6154 => x"81",
          6155 => x"07",
          6156 => x"2e",
          6157 => x"16",
          6158 => x"2e",
          6159 => x"88",
          6160 => x"82",
          6161 => x"56",
          6162 => x"51",
          6163 => x"82",
          6164 => x"54",
          6165 => x"08",
          6166 => x"9b",
          6167 => x"2e",
          6168 => x"83",
          6169 => x"73",
          6170 => x"0c",
          6171 => x"04",
          6172 => x"76",
          6173 => x"54",
          6174 => x"82",
          6175 => x"83",
          6176 => x"76",
          6177 => x"53",
          6178 => x"2e",
          6179 => x"90",
          6180 => x"51",
          6181 => x"82",
          6182 => x"90",
          6183 => x"53",
          6184 => x"a8",
          6185 => x"0d",
          6186 => x"0d",
          6187 => x"83",
          6188 => x"54",
          6189 => x"55",
          6190 => x"3f",
          6191 => x"51",
          6192 => x"2e",
          6193 => x"8b",
          6194 => x"2a",
          6195 => x"51",
          6196 => x"86",
          6197 => x"f7",
          6198 => x"7d",
          6199 => x"75",
          6200 => x"98",
          6201 => x"2e",
          6202 => x"98",
          6203 => x"78",
          6204 => x"3f",
          6205 => x"08",
          6206 => x"a8",
          6207 => x"38",
          6208 => x"70",
          6209 => x"73",
          6210 => x"58",
          6211 => x"8b",
          6212 => x"bf",
          6213 => x"ff",
          6214 => x"53",
          6215 => x"34",
          6216 => x"08",
          6217 => x"e5",
          6218 => x"81",
          6219 => x"2e",
          6220 => x"70",
          6221 => x"57",
          6222 => x"9e",
          6223 => x"2e",
          6224 => x"b5",
          6225 => x"df",
          6226 => x"72",
          6227 => x"81",
          6228 => x"76",
          6229 => x"2e",
          6230 => x"52",
          6231 => x"fc",
          6232 => x"a8",
          6233 => x"b5",
          6234 => x"38",
          6235 => x"fe",
          6236 => x"39",
          6237 => x"16",
          6238 => x"b5",
          6239 => x"3d",
          6240 => x"3d",
          6241 => x"08",
          6242 => x"52",
          6243 => x"c5",
          6244 => x"a8",
          6245 => x"b5",
          6246 => x"38",
          6247 => x"52",
          6248 => x"de",
          6249 => x"a8",
          6250 => x"b5",
          6251 => x"38",
          6252 => x"b5",
          6253 => x"9c",
          6254 => x"ea",
          6255 => x"53",
          6256 => x"9c",
          6257 => x"ea",
          6258 => x"0b",
          6259 => x"74",
          6260 => x"0c",
          6261 => x"04",
          6262 => x"75",
          6263 => x"12",
          6264 => x"53",
          6265 => x"9a",
          6266 => x"a8",
          6267 => x"9c",
          6268 => x"e5",
          6269 => x"0b",
          6270 => x"85",
          6271 => x"fa",
          6272 => x"7a",
          6273 => x"0b",
          6274 => x"98",
          6275 => x"2e",
          6276 => x"80",
          6277 => x"55",
          6278 => x"17",
          6279 => x"33",
          6280 => x"51",
          6281 => x"2e",
          6282 => x"85",
          6283 => x"06",
          6284 => x"e5",
          6285 => x"2e",
          6286 => x"8b",
          6287 => x"70",
          6288 => x"34",
          6289 => x"71",
          6290 => x"05",
          6291 => x"15",
          6292 => x"27",
          6293 => x"15",
          6294 => x"80",
          6295 => x"34",
          6296 => x"52",
          6297 => x"88",
          6298 => x"17",
          6299 => x"52",
          6300 => x"3f",
          6301 => x"08",
          6302 => x"12",
          6303 => x"3f",
          6304 => x"08",
          6305 => x"98",
          6306 => x"da",
          6307 => x"a8",
          6308 => x"23",
          6309 => x"04",
          6310 => x"7f",
          6311 => x"5b",
          6312 => x"33",
          6313 => x"73",
          6314 => x"38",
          6315 => x"80",
          6316 => x"38",
          6317 => x"8c",
          6318 => x"08",
          6319 => x"aa",
          6320 => x"41",
          6321 => x"33",
          6322 => x"73",
          6323 => x"81",
          6324 => x"81",
          6325 => x"dc",
          6326 => x"70",
          6327 => x"07",
          6328 => x"73",
          6329 => x"88",
          6330 => x"70",
          6331 => x"73",
          6332 => x"38",
          6333 => x"ab",
          6334 => x"52",
          6335 => x"91",
          6336 => x"a8",
          6337 => x"98",
          6338 => x"61",
          6339 => x"5a",
          6340 => x"a0",
          6341 => x"e7",
          6342 => x"70",
          6343 => x"79",
          6344 => x"73",
          6345 => x"81",
          6346 => x"38",
          6347 => x"33",
          6348 => x"ae",
          6349 => x"70",
          6350 => x"82",
          6351 => x"51",
          6352 => x"54",
          6353 => x"79",
          6354 => x"74",
          6355 => x"57",
          6356 => x"af",
          6357 => x"70",
          6358 => x"51",
          6359 => x"dc",
          6360 => x"73",
          6361 => x"38",
          6362 => x"82",
          6363 => x"19",
          6364 => x"54",
          6365 => x"82",
          6366 => x"54",
          6367 => x"78",
          6368 => x"81",
          6369 => x"54",
          6370 => x"81",
          6371 => x"af",
          6372 => x"77",
          6373 => x"70",
          6374 => x"25",
          6375 => x"07",
          6376 => x"51",
          6377 => x"2e",
          6378 => x"39",
          6379 => x"80",
          6380 => x"33",
          6381 => x"73",
          6382 => x"81",
          6383 => x"81",
          6384 => x"dc",
          6385 => x"70",
          6386 => x"07",
          6387 => x"73",
          6388 => x"b5",
          6389 => x"2e",
          6390 => x"83",
          6391 => x"76",
          6392 => x"07",
          6393 => x"2e",
          6394 => x"8b",
          6395 => x"77",
          6396 => x"30",
          6397 => x"71",
          6398 => x"53",
          6399 => x"55",
          6400 => x"38",
          6401 => x"5c",
          6402 => x"75",
          6403 => x"73",
          6404 => x"38",
          6405 => x"06",
          6406 => x"11",
          6407 => x"75",
          6408 => x"3f",
          6409 => x"08",
          6410 => x"38",
          6411 => x"33",
          6412 => x"54",
          6413 => x"e6",
          6414 => x"b5",
          6415 => x"2e",
          6416 => x"ff",
          6417 => x"74",
          6418 => x"38",
          6419 => x"75",
          6420 => x"17",
          6421 => x"57",
          6422 => x"a7",
          6423 => x"82",
          6424 => x"e5",
          6425 => x"b5",
          6426 => x"38",
          6427 => x"54",
          6428 => x"89",
          6429 => x"70",
          6430 => x"57",
          6431 => x"54",
          6432 => x"81",
          6433 => x"f7",
          6434 => x"7e",
          6435 => x"2e",
          6436 => x"33",
          6437 => x"e5",
          6438 => x"06",
          6439 => x"7a",
          6440 => x"a0",
          6441 => x"38",
          6442 => x"55",
          6443 => x"84",
          6444 => x"39",
          6445 => x"8b",
          6446 => x"7b",
          6447 => x"7a",
          6448 => x"3f",
          6449 => x"08",
          6450 => x"a8",
          6451 => x"38",
          6452 => x"52",
          6453 => x"aa",
          6454 => x"a8",
          6455 => x"b5",
          6456 => x"c2",
          6457 => x"08",
          6458 => x"55",
          6459 => x"ff",
          6460 => x"15",
          6461 => x"54",
          6462 => x"34",
          6463 => x"70",
          6464 => x"81",
          6465 => x"58",
          6466 => x"8b",
          6467 => x"74",
          6468 => x"3f",
          6469 => x"08",
          6470 => x"38",
          6471 => x"51",
          6472 => x"ff",
          6473 => x"ab",
          6474 => x"55",
          6475 => x"bb",
          6476 => x"2e",
          6477 => x"80",
          6478 => x"85",
          6479 => x"06",
          6480 => x"58",
          6481 => x"80",
          6482 => x"75",
          6483 => x"73",
          6484 => x"b5",
          6485 => x"0b",
          6486 => x"80",
          6487 => x"39",
          6488 => x"54",
          6489 => x"85",
          6490 => x"75",
          6491 => x"81",
          6492 => x"73",
          6493 => x"1b",
          6494 => x"2a",
          6495 => x"51",
          6496 => x"80",
          6497 => x"90",
          6498 => x"ff",
          6499 => x"05",
          6500 => x"f5",
          6501 => x"b5",
          6502 => x"1c",
          6503 => x"39",
          6504 => x"a8",
          6505 => x"0d",
          6506 => x"0d",
          6507 => x"7b",
          6508 => x"73",
          6509 => x"55",
          6510 => x"2e",
          6511 => x"75",
          6512 => x"57",
          6513 => x"26",
          6514 => x"ba",
          6515 => x"70",
          6516 => x"ba",
          6517 => x"06",
          6518 => x"73",
          6519 => x"70",
          6520 => x"51",
          6521 => x"89",
          6522 => x"82",
          6523 => x"ff",
          6524 => x"56",
          6525 => x"2e",
          6526 => x"80",
          6527 => x"e0",
          6528 => x"08",
          6529 => x"76",
          6530 => x"58",
          6531 => x"81",
          6532 => x"ff",
          6533 => x"53",
          6534 => x"26",
          6535 => x"13",
          6536 => x"06",
          6537 => x"9f",
          6538 => x"99",
          6539 => x"e0",
          6540 => x"ff",
          6541 => x"72",
          6542 => x"2a",
          6543 => x"72",
          6544 => x"06",
          6545 => x"ff",
          6546 => x"30",
          6547 => x"70",
          6548 => x"07",
          6549 => x"9f",
          6550 => x"54",
          6551 => x"80",
          6552 => x"81",
          6553 => x"59",
          6554 => x"25",
          6555 => x"8b",
          6556 => x"24",
          6557 => x"76",
          6558 => x"78",
          6559 => x"82",
          6560 => x"51",
          6561 => x"a8",
          6562 => x"0d",
          6563 => x"0d",
          6564 => x"0b",
          6565 => x"ff",
          6566 => x"0c",
          6567 => x"51",
          6568 => x"84",
          6569 => x"a8",
          6570 => x"38",
          6571 => x"51",
          6572 => x"82",
          6573 => x"83",
          6574 => x"54",
          6575 => x"82",
          6576 => x"09",
          6577 => x"e3",
          6578 => x"b4",
          6579 => x"57",
          6580 => x"2e",
          6581 => x"83",
          6582 => x"74",
          6583 => x"70",
          6584 => x"25",
          6585 => x"51",
          6586 => x"38",
          6587 => x"2e",
          6588 => x"b5",
          6589 => x"82",
          6590 => x"80",
          6591 => x"e0",
          6592 => x"b5",
          6593 => x"82",
          6594 => x"80",
          6595 => x"85",
          6596 => x"a4",
          6597 => x"16",
          6598 => x"3f",
          6599 => x"08",
          6600 => x"a8",
          6601 => x"83",
          6602 => x"74",
          6603 => x"0c",
          6604 => x"04",
          6605 => x"61",
          6606 => x"80",
          6607 => x"58",
          6608 => x"0c",
          6609 => x"e1",
          6610 => x"a8",
          6611 => x"56",
          6612 => x"b5",
          6613 => x"86",
          6614 => x"b5",
          6615 => x"29",
          6616 => x"05",
          6617 => x"53",
          6618 => x"80",
          6619 => x"38",
          6620 => x"76",
          6621 => x"74",
          6622 => x"72",
          6623 => x"38",
          6624 => x"51",
          6625 => x"82",
          6626 => x"81",
          6627 => x"81",
          6628 => x"72",
          6629 => x"80",
          6630 => x"38",
          6631 => x"70",
          6632 => x"53",
          6633 => x"86",
          6634 => x"a7",
          6635 => x"34",
          6636 => x"34",
          6637 => x"14",
          6638 => x"b2",
          6639 => x"a8",
          6640 => x"06",
          6641 => x"54",
          6642 => x"72",
          6643 => x"76",
          6644 => x"38",
          6645 => x"70",
          6646 => x"53",
          6647 => x"85",
          6648 => x"70",
          6649 => x"5b",
          6650 => x"82",
          6651 => x"81",
          6652 => x"76",
          6653 => x"81",
          6654 => x"38",
          6655 => x"56",
          6656 => x"83",
          6657 => x"70",
          6658 => x"80",
          6659 => x"83",
          6660 => x"dc",
          6661 => x"b5",
          6662 => x"76",
          6663 => x"05",
          6664 => x"16",
          6665 => x"56",
          6666 => x"d7",
          6667 => x"8d",
          6668 => x"72",
          6669 => x"54",
          6670 => x"57",
          6671 => x"95",
          6672 => x"73",
          6673 => x"3f",
          6674 => x"08",
          6675 => x"57",
          6676 => x"89",
          6677 => x"56",
          6678 => x"d7",
          6679 => x"76",
          6680 => x"f1",
          6681 => x"76",
          6682 => x"e9",
          6683 => x"51",
          6684 => x"82",
          6685 => x"83",
          6686 => x"53",
          6687 => x"2e",
          6688 => x"84",
          6689 => x"ca",
          6690 => x"da",
          6691 => x"a8",
          6692 => x"ff",
          6693 => x"8d",
          6694 => x"14",
          6695 => x"3f",
          6696 => x"08",
          6697 => x"15",
          6698 => x"14",
          6699 => x"34",
          6700 => x"33",
          6701 => x"81",
          6702 => x"54",
          6703 => x"72",
          6704 => x"91",
          6705 => x"ff",
          6706 => x"29",
          6707 => x"33",
          6708 => x"72",
          6709 => x"72",
          6710 => x"38",
          6711 => x"06",
          6712 => x"2e",
          6713 => x"56",
          6714 => x"80",
          6715 => x"da",
          6716 => x"b5",
          6717 => x"82",
          6718 => x"88",
          6719 => x"8f",
          6720 => x"56",
          6721 => x"38",
          6722 => x"51",
          6723 => x"82",
          6724 => x"83",
          6725 => x"55",
          6726 => x"80",
          6727 => x"da",
          6728 => x"b5",
          6729 => x"80",
          6730 => x"da",
          6731 => x"b5",
          6732 => x"ff",
          6733 => x"8d",
          6734 => x"2e",
          6735 => x"88",
          6736 => x"14",
          6737 => x"05",
          6738 => x"75",
          6739 => x"38",
          6740 => x"52",
          6741 => x"51",
          6742 => x"3f",
          6743 => x"08",
          6744 => x"a8",
          6745 => x"82",
          6746 => x"b5",
          6747 => x"ff",
          6748 => x"26",
          6749 => x"57",
          6750 => x"f5",
          6751 => x"82",
          6752 => x"f5",
          6753 => x"81",
          6754 => x"8d",
          6755 => x"2e",
          6756 => x"82",
          6757 => x"16",
          6758 => x"16",
          6759 => x"70",
          6760 => x"7a",
          6761 => x"0c",
          6762 => x"83",
          6763 => x"06",
          6764 => x"de",
          6765 => x"ae",
          6766 => x"a8",
          6767 => x"ff",
          6768 => x"56",
          6769 => x"38",
          6770 => x"38",
          6771 => x"51",
          6772 => x"82",
          6773 => x"a8",
          6774 => x"82",
          6775 => x"39",
          6776 => x"80",
          6777 => x"38",
          6778 => x"15",
          6779 => x"53",
          6780 => x"8d",
          6781 => x"15",
          6782 => x"76",
          6783 => x"51",
          6784 => x"13",
          6785 => x"8d",
          6786 => x"15",
          6787 => x"c5",
          6788 => x"90",
          6789 => x"0b",
          6790 => x"ff",
          6791 => x"15",
          6792 => x"2e",
          6793 => x"81",
          6794 => x"e4",
          6795 => x"b6",
          6796 => x"a8",
          6797 => x"ff",
          6798 => x"81",
          6799 => x"06",
          6800 => x"81",
          6801 => x"51",
          6802 => x"82",
          6803 => x"80",
          6804 => x"b5",
          6805 => x"15",
          6806 => x"14",
          6807 => x"3f",
          6808 => x"08",
          6809 => x"06",
          6810 => x"d4",
          6811 => x"81",
          6812 => x"38",
          6813 => x"d8",
          6814 => x"b5",
          6815 => x"8b",
          6816 => x"2e",
          6817 => x"b3",
          6818 => x"14",
          6819 => x"3f",
          6820 => x"08",
          6821 => x"e4",
          6822 => x"81",
          6823 => x"84",
          6824 => x"d7",
          6825 => x"b5",
          6826 => x"15",
          6827 => x"14",
          6828 => x"3f",
          6829 => x"08",
          6830 => x"76",
          6831 => x"cc",
          6832 => x"05",
          6833 => x"cc",
          6834 => x"86",
          6835 => x"0b",
          6836 => x"80",
          6837 => x"b5",
          6838 => x"3d",
          6839 => x"3d",
          6840 => x"89",
          6841 => x"2e",
          6842 => x"08",
          6843 => x"2e",
          6844 => x"33",
          6845 => x"2e",
          6846 => x"13",
          6847 => x"22",
          6848 => x"76",
          6849 => x"06",
          6850 => x"13",
          6851 => x"c0",
          6852 => x"a8",
          6853 => x"52",
          6854 => x"71",
          6855 => x"55",
          6856 => x"53",
          6857 => x"0c",
          6858 => x"b5",
          6859 => x"3d",
          6860 => x"3d",
          6861 => x"05",
          6862 => x"89",
          6863 => x"52",
          6864 => x"3f",
          6865 => x"0b",
          6866 => x"08",
          6867 => x"82",
          6868 => x"84",
          6869 => x"e0",
          6870 => x"55",
          6871 => x"2e",
          6872 => x"74",
          6873 => x"73",
          6874 => x"38",
          6875 => x"78",
          6876 => x"54",
          6877 => x"92",
          6878 => x"89",
          6879 => x"84",
          6880 => x"b0",
          6881 => x"a8",
          6882 => x"82",
          6883 => x"88",
          6884 => x"eb",
          6885 => x"02",
          6886 => x"e7",
          6887 => x"59",
          6888 => x"80",
          6889 => x"38",
          6890 => x"70",
          6891 => x"d0",
          6892 => x"3d",
          6893 => x"58",
          6894 => x"82",
          6895 => x"55",
          6896 => x"08",
          6897 => x"7a",
          6898 => x"8c",
          6899 => x"56",
          6900 => x"82",
          6901 => x"55",
          6902 => x"08",
          6903 => x"80",
          6904 => x"70",
          6905 => x"57",
          6906 => x"83",
          6907 => x"77",
          6908 => x"73",
          6909 => x"ab",
          6910 => x"2e",
          6911 => x"84",
          6912 => x"06",
          6913 => x"51",
          6914 => x"82",
          6915 => x"55",
          6916 => x"b2",
          6917 => x"06",
          6918 => x"b8",
          6919 => x"2a",
          6920 => x"51",
          6921 => x"2e",
          6922 => x"55",
          6923 => x"77",
          6924 => x"74",
          6925 => x"77",
          6926 => x"81",
          6927 => x"73",
          6928 => x"af",
          6929 => x"7a",
          6930 => x"3f",
          6931 => x"08",
          6932 => x"b2",
          6933 => x"8e",
          6934 => x"ea",
          6935 => x"a0",
          6936 => x"34",
          6937 => x"52",
          6938 => x"bd",
          6939 => x"62",
          6940 => x"d4",
          6941 => x"54",
          6942 => x"15",
          6943 => x"2e",
          6944 => x"7a",
          6945 => x"51",
          6946 => x"75",
          6947 => x"d4",
          6948 => x"be",
          6949 => x"a8",
          6950 => x"b5",
          6951 => x"ca",
          6952 => x"74",
          6953 => x"02",
          6954 => x"70",
          6955 => x"81",
          6956 => x"56",
          6957 => x"86",
          6958 => x"82",
          6959 => x"81",
          6960 => x"06",
          6961 => x"80",
          6962 => x"75",
          6963 => x"73",
          6964 => x"38",
          6965 => x"92",
          6966 => x"7a",
          6967 => x"3f",
          6968 => x"08",
          6969 => x"8c",
          6970 => x"55",
          6971 => x"08",
          6972 => x"77",
          6973 => x"81",
          6974 => x"73",
          6975 => x"38",
          6976 => x"07",
          6977 => x"11",
          6978 => x"0c",
          6979 => x"0c",
          6980 => x"52",
          6981 => x"3f",
          6982 => x"08",
          6983 => x"08",
          6984 => x"63",
          6985 => x"5a",
          6986 => x"82",
          6987 => x"82",
          6988 => x"8c",
          6989 => x"7a",
          6990 => x"17",
          6991 => x"23",
          6992 => x"34",
          6993 => x"1a",
          6994 => x"9c",
          6995 => x"0b",
          6996 => x"77",
          6997 => x"81",
          6998 => x"73",
          6999 => x"8d",
          7000 => x"a8",
          7001 => x"81",
          7002 => x"b5",
          7003 => x"1a",
          7004 => x"22",
          7005 => x"7b",
          7006 => x"a8",
          7007 => x"78",
          7008 => x"3f",
          7009 => x"08",
          7010 => x"a8",
          7011 => x"83",
          7012 => x"82",
          7013 => x"ff",
          7014 => x"06",
          7015 => x"55",
          7016 => x"56",
          7017 => x"76",
          7018 => x"51",
          7019 => x"27",
          7020 => x"70",
          7021 => x"5a",
          7022 => x"76",
          7023 => x"74",
          7024 => x"83",
          7025 => x"73",
          7026 => x"38",
          7027 => x"51",
          7028 => x"82",
          7029 => x"85",
          7030 => x"8e",
          7031 => x"2a",
          7032 => x"08",
          7033 => x"0c",
          7034 => x"79",
          7035 => x"73",
          7036 => x"0c",
          7037 => x"04",
          7038 => x"60",
          7039 => x"40",
          7040 => x"80",
          7041 => x"3d",
          7042 => x"78",
          7043 => x"3f",
          7044 => x"08",
          7045 => x"a8",
          7046 => x"91",
          7047 => x"74",
          7048 => x"38",
          7049 => x"c4",
          7050 => x"33",
          7051 => x"87",
          7052 => x"2e",
          7053 => x"95",
          7054 => x"91",
          7055 => x"56",
          7056 => x"81",
          7057 => x"34",
          7058 => x"a0",
          7059 => x"08",
          7060 => x"31",
          7061 => x"27",
          7062 => x"5c",
          7063 => x"82",
          7064 => x"19",
          7065 => x"ff",
          7066 => x"74",
          7067 => x"7e",
          7068 => x"ff",
          7069 => x"2a",
          7070 => x"79",
          7071 => x"87",
          7072 => x"08",
          7073 => x"98",
          7074 => x"78",
          7075 => x"3f",
          7076 => x"08",
          7077 => x"27",
          7078 => x"74",
          7079 => x"a3",
          7080 => x"1a",
          7081 => x"08",
          7082 => x"d4",
          7083 => x"b5",
          7084 => x"2e",
          7085 => x"82",
          7086 => x"1a",
          7087 => x"59",
          7088 => x"2e",
          7089 => x"77",
          7090 => x"11",
          7091 => x"55",
          7092 => x"85",
          7093 => x"31",
          7094 => x"76",
          7095 => x"81",
          7096 => x"ca",
          7097 => x"b5",
          7098 => x"d7",
          7099 => x"11",
          7100 => x"74",
          7101 => x"38",
          7102 => x"77",
          7103 => x"78",
          7104 => x"84",
          7105 => x"16",
          7106 => x"08",
          7107 => x"2b",
          7108 => x"cf",
          7109 => x"89",
          7110 => x"39",
          7111 => x"0c",
          7112 => x"83",
          7113 => x"80",
          7114 => x"55",
          7115 => x"83",
          7116 => x"9c",
          7117 => x"7e",
          7118 => x"3f",
          7119 => x"08",
          7120 => x"75",
          7121 => x"08",
          7122 => x"1f",
          7123 => x"7c",
          7124 => x"3f",
          7125 => x"7e",
          7126 => x"0c",
          7127 => x"1b",
          7128 => x"1c",
          7129 => x"fd",
          7130 => x"56",
          7131 => x"a8",
          7132 => x"0d",
          7133 => x"0d",
          7134 => x"64",
          7135 => x"58",
          7136 => x"90",
          7137 => x"52",
          7138 => x"d2",
          7139 => x"a8",
          7140 => x"b5",
          7141 => x"38",
          7142 => x"55",
          7143 => x"86",
          7144 => x"83",
          7145 => x"18",
          7146 => x"2a",
          7147 => x"51",
          7148 => x"56",
          7149 => x"83",
          7150 => x"39",
          7151 => x"19",
          7152 => x"83",
          7153 => x"0b",
          7154 => x"81",
          7155 => x"39",
          7156 => x"7c",
          7157 => x"74",
          7158 => x"38",
          7159 => x"7b",
          7160 => x"ec",
          7161 => x"08",
          7162 => x"06",
          7163 => x"81",
          7164 => x"8a",
          7165 => x"05",
          7166 => x"06",
          7167 => x"bf",
          7168 => x"38",
          7169 => x"55",
          7170 => x"7a",
          7171 => x"98",
          7172 => x"77",
          7173 => x"3f",
          7174 => x"08",
          7175 => x"a8",
          7176 => x"82",
          7177 => x"81",
          7178 => x"38",
          7179 => x"ff",
          7180 => x"98",
          7181 => x"18",
          7182 => x"74",
          7183 => x"7e",
          7184 => x"08",
          7185 => x"2e",
          7186 => x"8d",
          7187 => x"ce",
          7188 => x"b5",
          7189 => x"ee",
          7190 => x"08",
          7191 => x"d1",
          7192 => x"b5",
          7193 => x"2e",
          7194 => x"82",
          7195 => x"1b",
          7196 => x"5a",
          7197 => x"2e",
          7198 => x"78",
          7199 => x"11",
          7200 => x"55",
          7201 => x"85",
          7202 => x"31",
          7203 => x"76",
          7204 => x"81",
          7205 => x"c8",
          7206 => x"b5",
          7207 => x"a6",
          7208 => x"11",
          7209 => x"56",
          7210 => x"27",
          7211 => x"80",
          7212 => x"08",
          7213 => x"2b",
          7214 => x"b4",
          7215 => x"b5",
          7216 => x"80",
          7217 => x"34",
          7218 => x"56",
          7219 => x"8c",
          7220 => x"19",
          7221 => x"38",
          7222 => x"b6",
          7223 => x"a8",
          7224 => x"38",
          7225 => x"12",
          7226 => x"9c",
          7227 => x"18",
          7228 => x"06",
          7229 => x"31",
          7230 => x"76",
          7231 => x"7b",
          7232 => x"08",
          7233 => x"cd",
          7234 => x"b5",
          7235 => x"b6",
          7236 => x"7c",
          7237 => x"08",
          7238 => x"1f",
          7239 => x"cb",
          7240 => x"55",
          7241 => x"16",
          7242 => x"31",
          7243 => x"7f",
          7244 => x"94",
          7245 => x"70",
          7246 => x"8c",
          7247 => x"58",
          7248 => x"76",
          7249 => x"75",
          7250 => x"19",
          7251 => x"39",
          7252 => x"80",
          7253 => x"74",
          7254 => x"80",
          7255 => x"b5",
          7256 => x"3d",
          7257 => x"3d",
          7258 => x"3d",
          7259 => x"70",
          7260 => x"ea",
          7261 => x"a8",
          7262 => x"b5",
          7263 => x"fb",
          7264 => x"33",
          7265 => x"70",
          7266 => x"55",
          7267 => x"2e",
          7268 => x"a0",
          7269 => x"78",
          7270 => x"3f",
          7271 => x"08",
          7272 => x"a8",
          7273 => x"38",
          7274 => x"8b",
          7275 => x"07",
          7276 => x"8b",
          7277 => x"16",
          7278 => x"52",
          7279 => x"dd",
          7280 => x"16",
          7281 => x"15",
          7282 => x"3f",
          7283 => x"0a",
          7284 => x"51",
          7285 => x"76",
          7286 => x"51",
          7287 => x"78",
          7288 => x"83",
          7289 => x"51",
          7290 => x"82",
          7291 => x"90",
          7292 => x"bf",
          7293 => x"73",
          7294 => x"76",
          7295 => x"0c",
          7296 => x"04",
          7297 => x"76",
          7298 => x"fe",
          7299 => x"b5",
          7300 => x"82",
          7301 => x"9c",
          7302 => x"fc",
          7303 => x"51",
          7304 => x"82",
          7305 => x"53",
          7306 => x"08",
          7307 => x"b5",
          7308 => x"0c",
          7309 => x"a8",
          7310 => x"0d",
          7311 => x"0d",
          7312 => x"e6",
          7313 => x"52",
          7314 => x"b5",
          7315 => x"8b",
          7316 => x"a8",
          7317 => x"f4",
          7318 => x"71",
          7319 => x"0c",
          7320 => x"04",
          7321 => x"80",
          7322 => x"d0",
          7323 => x"3d",
          7324 => x"3f",
          7325 => x"08",
          7326 => x"a8",
          7327 => x"38",
          7328 => x"52",
          7329 => x"05",
          7330 => x"3f",
          7331 => x"08",
          7332 => x"a8",
          7333 => x"02",
          7334 => x"33",
          7335 => x"55",
          7336 => x"25",
          7337 => x"7a",
          7338 => x"54",
          7339 => x"a2",
          7340 => x"84",
          7341 => x"06",
          7342 => x"73",
          7343 => x"38",
          7344 => x"70",
          7345 => x"a8",
          7346 => x"a8",
          7347 => x"0c",
          7348 => x"b5",
          7349 => x"2e",
          7350 => x"83",
          7351 => x"74",
          7352 => x"0c",
          7353 => x"04",
          7354 => x"6f",
          7355 => x"80",
          7356 => x"53",
          7357 => x"b8",
          7358 => x"3d",
          7359 => x"3f",
          7360 => x"08",
          7361 => x"a8",
          7362 => x"38",
          7363 => x"7c",
          7364 => x"47",
          7365 => x"54",
          7366 => x"81",
          7367 => x"52",
          7368 => x"52",
          7369 => x"3f",
          7370 => x"08",
          7371 => x"a8",
          7372 => x"38",
          7373 => x"51",
          7374 => x"82",
          7375 => x"57",
          7376 => x"08",
          7377 => x"69",
          7378 => x"da",
          7379 => x"b5",
          7380 => x"76",
          7381 => x"d5",
          7382 => x"b5",
          7383 => x"82",
          7384 => x"82",
          7385 => x"52",
          7386 => x"eb",
          7387 => x"a8",
          7388 => x"b5",
          7389 => x"38",
          7390 => x"51",
          7391 => x"73",
          7392 => x"08",
          7393 => x"76",
          7394 => x"d6",
          7395 => x"b5",
          7396 => x"82",
          7397 => x"80",
          7398 => x"76",
          7399 => x"81",
          7400 => x"82",
          7401 => x"39",
          7402 => x"38",
          7403 => x"bc",
          7404 => x"51",
          7405 => x"76",
          7406 => x"11",
          7407 => x"51",
          7408 => x"73",
          7409 => x"38",
          7410 => x"55",
          7411 => x"16",
          7412 => x"56",
          7413 => x"38",
          7414 => x"73",
          7415 => x"90",
          7416 => x"2e",
          7417 => x"16",
          7418 => x"ff",
          7419 => x"ff",
          7420 => x"58",
          7421 => x"74",
          7422 => x"75",
          7423 => x"18",
          7424 => x"58",
          7425 => x"fe",
          7426 => x"7b",
          7427 => x"06",
          7428 => x"18",
          7429 => x"58",
          7430 => x"80",
          7431 => x"f4",
          7432 => x"29",
          7433 => x"05",
          7434 => x"33",
          7435 => x"56",
          7436 => x"2e",
          7437 => x"16",
          7438 => x"33",
          7439 => x"73",
          7440 => x"16",
          7441 => x"26",
          7442 => x"55",
          7443 => x"91",
          7444 => x"54",
          7445 => x"70",
          7446 => x"34",
          7447 => x"ec",
          7448 => x"70",
          7449 => x"34",
          7450 => x"09",
          7451 => x"38",
          7452 => x"39",
          7453 => x"19",
          7454 => x"33",
          7455 => x"05",
          7456 => x"78",
          7457 => x"80",
          7458 => x"82",
          7459 => x"9e",
          7460 => x"f7",
          7461 => x"7d",
          7462 => x"05",
          7463 => x"57",
          7464 => x"3f",
          7465 => x"08",
          7466 => x"a8",
          7467 => x"38",
          7468 => x"53",
          7469 => x"38",
          7470 => x"54",
          7471 => x"92",
          7472 => x"33",
          7473 => x"70",
          7474 => x"54",
          7475 => x"38",
          7476 => x"15",
          7477 => x"70",
          7478 => x"58",
          7479 => x"82",
          7480 => x"8a",
          7481 => x"89",
          7482 => x"53",
          7483 => x"b7",
          7484 => x"ff",
          7485 => x"e8",
          7486 => x"b5",
          7487 => x"15",
          7488 => x"53",
          7489 => x"e8",
          7490 => x"b5",
          7491 => x"26",
          7492 => x"30",
          7493 => x"70",
          7494 => x"77",
          7495 => x"18",
          7496 => x"51",
          7497 => x"88",
          7498 => x"73",
          7499 => x"52",
          7500 => x"ca",
          7501 => x"a8",
          7502 => x"b5",
          7503 => x"2e",
          7504 => x"82",
          7505 => x"ff",
          7506 => x"38",
          7507 => x"08",
          7508 => x"73",
          7509 => x"73",
          7510 => x"9c",
          7511 => x"27",
          7512 => x"75",
          7513 => x"16",
          7514 => x"17",
          7515 => x"33",
          7516 => x"70",
          7517 => x"55",
          7518 => x"80",
          7519 => x"73",
          7520 => x"cc",
          7521 => x"b5",
          7522 => x"82",
          7523 => x"94",
          7524 => x"a8",
          7525 => x"39",
          7526 => x"51",
          7527 => x"82",
          7528 => x"54",
          7529 => x"be",
          7530 => x"27",
          7531 => x"53",
          7532 => x"08",
          7533 => x"73",
          7534 => x"ff",
          7535 => x"15",
          7536 => x"16",
          7537 => x"ff",
          7538 => x"80",
          7539 => x"73",
          7540 => x"c6",
          7541 => x"b5",
          7542 => x"38",
          7543 => x"16",
          7544 => x"80",
          7545 => x"0b",
          7546 => x"81",
          7547 => x"75",
          7548 => x"b5",
          7549 => x"58",
          7550 => x"54",
          7551 => x"74",
          7552 => x"73",
          7553 => x"90",
          7554 => x"c0",
          7555 => x"90",
          7556 => x"83",
          7557 => x"72",
          7558 => x"38",
          7559 => x"08",
          7560 => x"77",
          7561 => x"80",
          7562 => x"b5",
          7563 => x"3d",
          7564 => x"3d",
          7565 => x"89",
          7566 => x"2e",
          7567 => x"80",
          7568 => x"fc",
          7569 => x"3d",
          7570 => x"e1",
          7571 => x"b5",
          7572 => x"82",
          7573 => x"80",
          7574 => x"76",
          7575 => x"75",
          7576 => x"3f",
          7577 => x"08",
          7578 => x"a8",
          7579 => x"38",
          7580 => x"70",
          7581 => x"57",
          7582 => x"a2",
          7583 => x"33",
          7584 => x"70",
          7585 => x"55",
          7586 => x"2e",
          7587 => x"16",
          7588 => x"51",
          7589 => x"82",
          7590 => x"88",
          7591 => x"54",
          7592 => x"84",
          7593 => x"52",
          7594 => x"e5",
          7595 => x"a8",
          7596 => x"84",
          7597 => x"06",
          7598 => x"55",
          7599 => x"80",
          7600 => x"80",
          7601 => x"54",
          7602 => x"a8",
          7603 => x"0d",
          7604 => x"0d",
          7605 => x"fc",
          7606 => x"52",
          7607 => x"3f",
          7608 => x"08",
          7609 => x"b5",
          7610 => x"0c",
          7611 => x"04",
          7612 => x"77",
          7613 => x"fc",
          7614 => x"53",
          7615 => x"de",
          7616 => x"a8",
          7617 => x"b5",
          7618 => x"df",
          7619 => x"38",
          7620 => x"08",
          7621 => x"cd",
          7622 => x"b5",
          7623 => x"80",
          7624 => x"b5",
          7625 => x"73",
          7626 => x"3f",
          7627 => x"08",
          7628 => x"a8",
          7629 => x"09",
          7630 => x"38",
          7631 => x"39",
          7632 => x"08",
          7633 => x"52",
          7634 => x"b3",
          7635 => x"73",
          7636 => x"3f",
          7637 => x"08",
          7638 => x"30",
          7639 => x"9f",
          7640 => x"b5",
          7641 => x"51",
          7642 => x"72",
          7643 => x"0c",
          7644 => x"04",
          7645 => x"65",
          7646 => x"89",
          7647 => x"96",
          7648 => x"df",
          7649 => x"b5",
          7650 => x"82",
          7651 => x"b2",
          7652 => x"75",
          7653 => x"3f",
          7654 => x"08",
          7655 => x"a8",
          7656 => x"02",
          7657 => x"33",
          7658 => x"55",
          7659 => x"25",
          7660 => x"55",
          7661 => x"80",
          7662 => x"76",
          7663 => x"d4",
          7664 => x"82",
          7665 => x"94",
          7666 => x"f0",
          7667 => x"65",
          7668 => x"53",
          7669 => x"05",
          7670 => x"51",
          7671 => x"82",
          7672 => x"5b",
          7673 => x"08",
          7674 => x"7c",
          7675 => x"08",
          7676 => x"fe",
          7677 => x"08",
          7678 => x"55",
          7679 => x"91",
          7680 => x"0c",
          7681 => x"81",
          7682 => x"39",
          7683 => x"c7",
          7684 => x"a8",
          7685 => x"55",
          7686 => x"2e",
          7687 => x"bf",
          7688 => x"5f",
          7689 => x"92",
          7690 => x"51",
          7691 => x"82",
          7692 => x"ff",
          7693 => x"82",
          7694 => x"81",
          7695 => x"82",
          7696 => x"30",
          7697 => x"a8",
          7698 => x"25",
          7699 => x"19",
          7700 => x"5a",
          7701 => x"08",
          7702 => x"38",
          7703 => x"a4",
          7704 => x"b5",
          7705 => x"58",
          7706 => x"77",
          7707 => x"7d",
          7708 => x"bf",
          7709 => x"b5",
          7710 => x"82",
          7711 => x"80",
          7712 => x"70",
          7713 => x"ff",
          7714 => x"56",
          7715 => x"2e",
          7716 => x"9e",
          7717 => x"51",
          7718 => x"3f",
          7719 => x"08",
          7720 => x"06",
          7721 => x"80",
          7722 => x"19",
          7723 => x"54",
          7724 => x"14",
          7725 => x"c5",
          7726 => x"a8",
          7727 => x"06",
          7728 => x"80",
          7729 => x"19",
          7730 => x"54",
          7731 => x"06",
          7732 => x"79",
          7733 => x"78",
          7734 => x"79",
          7735 => x"84",
          7736 => x"07",
          7737 => x"84",
          7738 => x"82",
          7739 => x"92",
          7740 => x"f9",
          7741 => x"8a",
          7742 => x"53",
          7743 => x"e3",
          7744 => x"b5",
          7745 => x"82",
          7746 => x"81",
          7747 => x"17",
          7748 => x"81",
          7749 => x"17",
          7750 => x"2a",
          7751 => x"51",
          7752 => x"55",
          7753 => x"81",
          7754 => x"17",
          7755 => x"8c",
          7756 => x"81",
          7757 => x"9b",
          7758 => x"a8",
          7759 => x"17",
          7760 => x"51",
          7761 => x"82",
          7762 => x"74",
          7763 => x"56",
          7764 => x"98",
          7765 => x"76",
          7766 => x"c6",
          7767 => x"a8",
          7768 => x"09",
          7769 => x"38",
          7770 => x"b5",
          7771 => x"2e",
          7772 => x"85",
          7773 => x"a3",
          7774 => x"38",
          7775 => x"b5",
          7776 => x"15",
          7777 => x"38",
          7778 => x"53",
          7779 => x"08",
          7780 => x"c3",
          7781 => x"b5",
          7782 => x"94",
          7783 => x"18",
          7784 => x"33",
          7785 => x"54",
          7786 => x"34",
          7787 => x"85",
          7788 => x"18",
          7789 => x"74",
          7790 => x"0c",
          7791 => x"04",
          7792 => x"82",
          7793 => x"ff",
          7794 => x"a1",
          7795 => x"e4",
          7796 => x"a8",
          7797 => x"b5",
          7798 => x"f5",
          7799 => x"a1",
          7800 => x"95",
          7801 => x"58",
          7802 => x"82",
          7803 => x"55",
          7804 => x"08",
          7805 => x"02",
          7806 => x"33",
          7807 => x"70",
          7808 => x"55",
          7809 => x"73",
          7810 => x"75",
          7811 => x"80",
          7812 => x"bd",
          7813 => x"d6",
          7814 => x"81",
          7815 => x"87",
          7816 => x"ad",
          7817 => x"78",
          7818 => x"3f",
          7819 => x"08",
          7820 => x"70",
          7821 => x"55",
          7822 => x"2e",
          7823 => x"78",
          7824 => x"a8",
          7825 => x"08",
          7826 => x"38",
          7827 => x"b5",
          7828 => x"76",
          7829 => x"70",
          7830 => x"b5",
          7831 => x"a8",
          7832 => x"b5",
          7833 => x"e9",
          7834 => x"a8",
          7835 => x"51",
          7836 => x"82",
          7837 => x"55",
          7838 => x"08",
          7839 => x"55",
          7840 => x"82",
          7841 => x"84",
          7842 => x"82",
          7843 => x"80",
          7844 => x"51",
          7845 => x"82",
          7846 => x"82",
          7847 => x"30",
          7848 => x"a8",
          7849 => x"25",
          7850 => x"75",
          7851 => x"38",
          7852 => x"8f",
          7853 => x"75",
          7854 => x"c1",
          7855 => x"b5",
          7856 => x"74",
          7857 => x"51",
          7858 => x"3f",
          7859 => x"08",
          7860 => x"b5",
          7861 => x"3d",
          7862 => x"3d",
          7863 => x"99",
          7864 => x"52",
          7865 => x"d8",
          7866 => x"b5",
          7867 => x"82",
          7868 => x"82",
          7869 => x"5e",
          7870 => x"3d",
          7871 => x"cf",
          7872 => x"b5",
          7873 => x"82",
          7874 => x"86",
          7875 => x"82",
          7876 => x"b5",
          7877 => x"2e",
          7878 => x"82",
          7879 => x"80",
          7880 => x"70",
          7881 => x"06",
          7882 => x"54",
          7883 => x"38",
          7884 => x"52",
          7885 => x"52",
          7886 => x"3f",
          7887 => x"08",
          7888 => x"82",
          7889 => x"83",
          7890 => x"82",
          7891 => x"81",
          7892 => x"06",
          7893 => x"54",
          7894 => x"08",
          7895 => x"81",
          7896 => x"81",
          7897 => x"39",
          7898 => x"38",
          7899 => x"08",
          7900 => x"c4",
          7901 => x"b5",
          7902 => x"82",
          7903 => x"81",
          7904 => x"53",
          7905 => x"19",
          7906 => x"8c",
          7907 => x"ae",
          7908 => x"34",
          7909 => x"0b",
          7910 => x"82",
          7911 => x"52",
          7912 => x"51",
          7913 => x"3f",
          7914 => x"b4",
          7915 => x"c9",
          7916 => x"53",
          7917 => x"53",
          7918 => x"51",
          7919 => x"3f",
          7920 => x"0b",
          7921 => x"34",
          7922 => x"80",
          7923 => x"51",
          7924 => x"78",
          7925 => x"83",
          7926 => x"51",
          7927 => x"82",
          7928 => x"54",
          7929 => x"08",
          7930 => x"88",
          7931 => x"64",
          7932 => x"ff",
          7933 => x"75",
          7934 => x"78",
          7935 => x"3f",
          7936 => x"0b",
          7937 => x"78",
          7938 => x"83",
          7939 => x"51",
          7940 => x"3f",
          7941 => x"08",
          7942 => x"80",
          7943 => x"76",
          7944 => x"ae",
          7945 => x"b5",
          7946 => x"3d",
          7947 => x"3d",
          7948 => x"84",
          7949 => x"f1",
          7950 => x"a8",
          7951 => x"05",
          7952 => x"51",
          7953 => x"82",
          7954 => x"55",
          7955 => x"08",
          7956 => x"78",
          7957 => x"08",
          7958 => x"70",
          7959 => x"b8",
          7960 => x"a8",
          7961 => x"b5",
          7962 => x"b9",
          7963 => x"9b",
          7964 => x"a0",
          7965 => x"55",
          7966 => x"38",
          7967 => x"3d",
          7968 => x"3d",
          7969 => x"51",
          7970 => x"3f",
          7971 => x"52",
          7972 => x"52",
          7973 => x"dd",
          7974 => x"08",
          7975 => x"cb",
          7976 => x"b5",
          7977 => x"82",
          7978 => x"95",
          7979 => x"2e",
          7980 => x"88",
          7981 => x"3d",
          7982 => x"38",
          7983 => x"e5",
          7984 => x"a8",
          7985 => x"09",
          7986 => x"b8",
          7987 => x"c9",
          7988 => x"b5",
          7989 => x"82",
          7990 => x"81",
          7991 => x"56",
          7992 => x"3d",
          7993 => x"52",
          7994 => x"ff",
          7995 => x"02",
          7996 => x"8b",
          7997 => x"16",
          7998 => x"2a",
          7999 => x"51",
          8000 => x"89",
          8001 => x"07",
          8002 => x"17",
          8003 => x"81",
          8004 => x"34",
          8005 => x"70",
          8006 => x"81",
          8007 => x"55",
          8008 => x"80",
          8009 => x"64",
          8010 => x"38",
          8011 => x"51",
          8012 => x"82",
          8013 => x"52",
          8014 => x"b7",
          8015 => x"55",
          8016 => x"08",
          8017 => x"dd",
          8018 => x"a8",
          8019 => x"51",
          8020 => x"3f",
          8021 => x"08",
          8022 => x"11",
          8023 => x"82",
          8024 => x"80",
          8025 => x"16",
          8026 => x"ae",
          8027 => x"06",
          8028 => x"53",
          8029 => x"51",
          8030 => x"78",
          8031 => x"83",
          8032 => x"39",
          8033 => x"08",
          8034 => x"51",
          8035 => x"82",
          8036 => x"55",
          8037 => x"08",
          8038 => x"51",
          8039 => x"3f",
          8040 => x"08",
          8041 => x"b5",
          8042 => x"3d",
          8043 => x"3d",
          8044 => x"db",
          8045 => x"84",
          8046 => x"05",
          8047 => x"82",
          8048 => x"d0",
          8049 => x"3d",
          8050 => x"3f",
          8051 => x"08",
          8052 => x"a8",
          8053 => x"38",
          8054 => x"52",
          8055 => x"05",
          8056 => x"3f",
          8057 => x"08",
          8058 => x"a8",
          8059 => x"02",
          8060 => x"33",
          8061 => x"54",
          8062 => x"aa",
          8063 => x"06",
          8064 => x"8b",
          8065 => x"06",
          8066 => x"07",
          8067 => x"56",
          8068 => x"34",
          8069 => x"0b",
          8070 => x"78",
          8071 => x"a9",
          8072 => x"a8",
          8073 => x"82",
          8074 => x"95",
          8075 => x"ef",
          8076 => x"56",
          8077 => x"3d",
          8078 => x"94",
          8079 => x"f4",
          8080 => x"a8",
          8081 => x"b5",
          8082 => x"cb",
          8083 => x"63",
          8084 => x"d4",
          8085 => x"c0",
          8086 => x"a8",
          8087 => x"b5",
          8088 => x"38",
          8089 => x"05",
          8090 => x"06",
          8091 => x"73",
          8092 => x"16",
          8093 => x"22",
          8094 => x"07",
          8095 => x"1f",
          8096 => x"c2",
          8097 => x"81",
          8098 => x"34",
          8099 => x"b3",
          8100 => x"b5",
          8101 => x"74",
          8102 => x"0c",
          8103 => x"04",
          8104 => x"69",
          8105 => x"80",
          8106 => x"d0",
          8107 => x"3d",
          8108 => x"3f",
          8109 => x"08",
          8110 => x"08",
          8111 => x"b5",
          8112 => x"80",
          8113 => x"57",
          8114 => x"81",
          8115 => x"70",
          8116 => x"55",
          8117 => x"80",
          8118 => x"5d",
          8119 => x"52",
          8120 => x"52",
          8121 => x"a9",
          8122 => x"a8",
          8123 => x"b5",
          8124 => x"d1",
          8125 => x"73",
          8126 => x"3f",
          8127 => x"08",
          8128 => x"a8",
          8129 => x"82",
          8130 => x"82",
          8131 => x"65",
          8132 => x"78",
          8133 => x"7b",
          8134 => x"55",
          8135 => x"34",
          8136 => x"8a",
          8137 => x"38",
          8138 => x"1a",
          8139 => x"34",
          8140 => x"9e",
          8141 => x"70",
          8142 => x"51",
          8143 => x"a0",
          8144 => x"8e",
          8145 => x"2e",
          8146 => x"86",
          8147 => x"34",
          8148 => x"30",
          8149 => x"80",
          8150 => x"7a",
          8151 => x"c1",
          8152 => x"2e",
          8153 => x"a0",
          8154 => x"51",
          8155 => x"3f",
          8156 => x"08",
          8157 => x"a8",
          8158 => x"7b",
          8159 => x"55",
          8160 => x"73",
          8161 => x"38",
          8162 => x"73",
          8163 => x"38",
          8164 => x"15",
          8165 => x"ff",
          8166 => x"82",
          8167 => x"7b",
          8168 => x"b5",
          8169 => x"3d",
          8170 => x"3d",
          8171 => x"9c",
          8172 => x"05",
          8173 => x"51",
          8174 => x"82",
          8175 => x"82",
          8176 => x"56",
          8177 => x"a8",
          8178 => x"38",
          8179 => x"52",
          8180 => x"52",
          8181 => x"c0",
          8182 => x"70",
          8183 => x"ff",
          8184 => x"55",
          8185 => x"27",
          8186 => x"78",
          8187 => x"ff",
          8188 => x"05",
          8189 => x"55",
          8190 => x"3f",
          8191 => x"08",
          8192 => x"38",
          8193 => x"70",
          8194 => x"ff",
          8195 => x"82",
          8196 => x"80",
          8197 => x"74",
          8198 => x"07",
          8199 => x"4e",
          8200 => x"82",
          8201 => x"55",
          8202 => x"70",
          8203 => x"06",
          8204 => x"99",
          8205 => x"e0",
          8206 => x"ff",
          8207 => x"54",
          8208 => x"27",
          8209 => x"ad",
          8210 => x"55",
          8211 => x"a3",
          8212 => x"82",
          8213 => x"ff",
          8214 => x"82",
          8215 => x"93",
          8216 => x"75",
          8217 => x"76",
          8218 => x"38",
          8219 => x"77",
          8220 => x"86",
          8221 => x"39",
          8222 => x"27",
          8223 => x"88",
          8224 => x"78",
          8225 => x"5a",
          8226 => x"57",
          8227 => x"81",
          8228 => x"81",
          8229 => x"33",
          8230 => x"06",
          8231 => x"57",
          8232 => x"fe",
          8233 => x"3d",
          8234 => x"55",
          8235 => x"2e",
          8236 => x"76",
          8237 => x"38",
          8238 => x"55",
          8239 => x"33",
          8240 => x"a0",
          8241 => x"06",
          8242 => x"17",
          8243 => x"38",
          8244 => x"43",
          8245 => x"3d",
          8246 => x"ff",
          8247 => x"82",
          8248 => x"54",
          8249 => x"08",
          8250 => x"81",
          8251 => x"ff",
          8252 => x"82",
          8253 => x"54",
          8254 => x"08",
          8255 => x"80",
          8256 => x"54",
          8257 => x"80",
          8258 => x"b5",
          8259 => x"2e",
          8260 => x"80",
          8261 => x"54",
          8262 => x"80",
          8263 => x"52",
          8264 => x"bd",
          8265 => x"b5",
          8266 => x"82",
          8267 => x"b1",
          8268 => x"82",
          8269 => x"52",
          8270 => x"ab",
          8271 => x"54",
          8272 => x"15",
          8273 => x"78",
          8274 => x"ff",
          8275 => x"79",
          8276 => x"83",
          8277 => x"51",
          8278 => x"3f",
          8279 => x"08",
          8280 => x"74",
          8281 => x"0c",
          8282 => x"04",
          8283 => x"60",
          8284 => x"05",
          8285 => x"33",
          8286 => x"05",
          8287 => x"40",
          8288 => x"da",
          8289 => x"a8",
          8290 => x"b5",
          8291 => x"bd",
          8292 => x"33",
          8293 => x"b5",
          8294 => x"2e",
          8295 => x"1a",
          8296 => x"90",
          8297 => x"33",
          8298 => x"70",
          8299 => x"55",
          8300 => x"38",
          8301 => x"97",
          8302 => x"82",
          8303 => x"58",
          8304 => x"7e",
          8305 => x"70",
          8306 => x"55",
          8307 => x"56",
          8308 => x"d1",
          8309 => x"7d",
          8310 => x"70",
          8311 => x"2a",
          8312 => x"08",
          8313 => x"08",
          8314 => x"5d",
          8315 => x"77",
          8316 => x"98",
          8317 => x"26",
          8318 => x"57",
          8319 => x"59",
          8320 => x"52",
          8321 => x"ae",
          8322 => x"15",
          8323 => x"98",
          8324 => x"26",
          8325 => x"55",
          8326 => x"08",
          8327 => x"99",
          8328 => x"a8",
          8329 => x"ff",
          8330 => x"b5",
          8331 => x"38",
          8332 => x"75",
          8333 => x"81",
          8334 => x"93",
          8335 => x"80",
          8336 => x"2e",
          8337 => x"ff",
          8338 => x"58",
          8339 => x"7d",
          8340 => x"38",
          8341 => x"55",
          8342 => x"b4",
          8343 => x"56",
          8344 => x"09",
          8345 => x"38",
          8346 => x"53",
          8347 => x"51",
          8348 => x"3f",
          8349 => x"08",
          8350 => x"a8",
          8351 => x"38",
          8352 => x"ff",
          8353 => x"5c",
          8354 => x"84",
          8355 => x"5c",
          8356 => x"12",
          8357 => x"80",
          8358 => x"78",
          8359 => x"7c",
          8360 => x"90",
          8361 => x"c0",
          8362 => x"90",
          8363 => x"15",
          8364 => x"90",
          8365 => x"54",
          8366 => x"91",
          8367 => x"31",
          8368 => x"84",
          8369 => x"07",
          8370 => x"16",
          8371 => x"73",
          8372 => x"0c",
          8373 => x"04",
          8374 => x"6b",
          8375 => x"05",
          8376 => x"33",
          8377 => x"5a",
          8378 => x"bd",
          8379 => x"80",
          8380 => x"a8",
          8381 => x"f8",
          8382 => x"a8",
          8383 => x"82",
          8384 => x"70",
          8385 => x"74",
          8386 => x"38",
          8387 => x"82",
          8388 => x"81",
          8389 => x"81",
          8390 => x"ff",
          8391 => x"82",
          8392 => x"81",
          8393 => x"81",
          8394 => x"83",
          8395 => x"c0",
          8396 => x"2a",
          8397 => x"51",
          8398 => x"74",
          8399 => x"99",
          8400 => x"53",
          8401 => x"51",
          8402 => x"3f",
          8403 => x"08",
          8404 => x"55",
          8405 => x"92",
          8406 => x"80",
          8407 => x"38",
          8408 => x"06",
          8409 => x"2e",
          8410 => x"48",
          8411 => x"87",
          8412 => x"79",
          8413 => x"78",
          8414 => x"26",
          8415 => x"19",
          8416 => x"74",
          8417 => x"38",
          8418 => x"e4",
          8419 => x"2a",
          8420 => x"70",
          8421 => x"59",
          8422 => x"7a",
          8423 => x"56",
          8424 => x"80",
          8425 => x"51",
          8426 => x"74",
          8427 => x"99",
          8428 => x"53",
          8429 => x"51",
          8430 => x"3f",
          8431 => x"b5",
          8432 => x"ac",
          8433 => x"2a",
          8434 => x"82",
          8435 => x"43",
          8436 => x"83",
          8437 => x"66",
          8438 => x"60",
          8439 => x"90",
          8440 => x"31",
          8441 => x"80",
          8442 => x"8a",
          8443 => x"56",
          8444 => x"26",
          8445 => x"77",
          8446 => x"81",
          8447 => x"74",
          8448 => x"38",
          8449 => x"55",
          8450 => x"83",
          8451 => x"81",
          8452 => x"80",
          8453 => x"38",
          8454 => x"55",
          8455 => x"5e",
          8456 => x"89",
          8457 => x"5a",
          8458 => x"09",
          8459 => x"e1",
          8460 => x"38",
          8461 => x"57",
          8462 => x"b0",
          8463 => x"5a",
          8464 => x"9d",
          8465 => x"26",
          8466 => x"b0",
          8467 => x"10",
          8468 => x"22",
          8469 => x"74",
          8470 => x"38",
          8471 => x"ee",
          8472 => x"66",
          8473 => x"bd",
          8474 => x"a8",
          8475 => x"84",
          8476 => x"89",
          8477 => x"a0",
          8478 => x"82",
          8479 => x"fc",
          8480 => x"56",
          8481 => x"f0",
          8482 => x"80",
          8483 => x"d3",
          8484 => x"38",
          8485 => x"57",
          8486 => x"b0",
          8487 => x"5a",
          8488 => x"9d",
          8489 => x"26",
          8490 => x"b0",
          8491 => x"10",
          8492 => x"22",
          8493 => x"74",
          8494 => x"38",
          8495 => x"ee",
          8496 => x"66",
          8497 => x"dd",
          8498 => x"a8",
          8499 => x"05",
          8500 => x"a8",
          8501 => x"26",
          8502 => x"0b",
          8503 => x"08",
          8504 => x"a8",
          8505 => x"11",
          8506 => x"05",
          8507 => x"83",
          8508 => x"2a",
          8509 => x"a0",
          8510 => x"7d",
          8511 => x"69",
          8512 => x"05",
          8513 => x"72",
          8514 => x"5c",
          8515 => x"59",
          8516 => x"2e",
          8517 => x"89",
          8518 => x"60",
          8519 => x"84",
          8520 => x"5d",
          8521 => x"18",
          8522 => x"68",
          8523 => x"74",
          8524 => x"af",
          8525 => x"31",
          8526 => x"53",
          8527 => x"52",
          8528 => x"e1",
          8529 => x"a8",
          8530 => x"83",
          8531 => x"06",
          8532 => x"b5",
          8533 => x"ff",
          8534 => x"dd",
          8535 => x"83",
          8536 => x"2a",
          8537 => x"be",
          8538 => x"39",
          8539 => x"09",
          8540 => x"c5",
          8541 => x"f5",
          8542 => x"a8",
          8543 => x"38",
          8544 => x"79",
          8545 => x"80",
          8546 => x"38",
          8547 => x"96",
          8548 => x"06",
          8549 => x"2e",
          8550 => x"5e",
          8551 => x"82",
          8552 => x"9f",
          8553 => x"38",
          8554 => x"38",
          8555 => x"81",
          8556 => x"fc",
          8557 => x"ab",
          8558 => x"7d",
          8559 => x"81",
          8560 => x"7d",
          8561 => x"78",
          8562 => x"74",
          8563 => x"8e",
          8564 => x"9c",
          8565 => x"53",
          8566 => x"51",
          8567 => x"3f",
          8568 => x"ae",
          8569 => x"51",
          8570 => x"3f",
          8571 => x"8b",
          8572 => x"a1",
          8573 => x"8d",
          8574 => x"83",
          8575 => x"52",
          8576 => x"ff",
          8577 => x"81",
          8578 => x"34",
          8579 => x"70",
          8580 => x"2a",
          8581 => x"54",
          8582 => x"1b",
          8583 => x"88",
          8584 => x"74",
          8585 => x"26",
          8586 => x"83",
          8587 => x"52",
          8588 => x"ff",
          8589 => x"8a",
          8590 => x"a0",
          8591 => x"a1",
          8592 => x"0b",
          8593 => x"bf",
          8594 => x"51",
          8595 => x"3f",
          8596 => x"9a",
          8597 => x"a0",
          8598 => x"52",
          8599 => x"ff",
          8600 => x"7d",
          8601 => x"81",
          8602 => x"38",
          8603 => x"0a",
          8604 => x"1b",
          8605 => x"ce",
          8606 => x"a4",
          8607 => x"a0",
          8608 => x"52",
          8609 => x"ff",
          8610 => x"81",
          8611 => x"51",
          8612 => x"3f",
          8613 => x"1b",
          8614 => x"8c",
          8615 => x"0b",
          8616 => x"34",
          8617 => x"c2",
          8618 => x"53",
          8619 => x"52",
          8620 => x"51",
          8621 => x"88",
          8622 => x"a7",
          8623 => x"a0",
          8624 => x"83",
          8625 => x"52",
          8626 => x"ff",
          8627 => x"ff",
          8628 => x"1c",
          8629 => x"a6",
          8630 => x"53",
          8631 => x"52",
          8632 => x"ff",
          8633 => x"82",
          8634 => x"83",
          8635 => x"52",
          8636 => x"b4",
          8637 => x"60",
          8638 => x"7e",
          8639 => x"d7",
          8640 => x"82",
          8641 => x"83",
          8642 => x"83",
          8643 => x"06",
          8644 => x"75",
          8645 => x"05",
          8646 => x"7e",
          8647 => x"b7",
          8648 => x"53",
          8649 => x"51",
          8650 => x"3f",
          8651 => x"a4",
          8652 => x"51",
          8653 => x"3f",
          8654 => x"e4",
          8655 => x"e4",
          8656 => x"9f",
          8657 => x"18",
          8658 => x"1b",
          8659 => x"f6",
          8660 => x"83",
          8661 => x"ff",
          8662 => x"82",
          8663 => x"78",
          8664 => x"c4",
          8665 => x"60",
          8666 => x"7a",
          8667 => x"ff",
          8668 => x"75",
          8669 => x"53",
          8670 => x"51",
          8671 => x"3f",
          8672 => x"52",
          8673 => x"9f",
          8674 => x"56",
          8675 => x"83",
          8676 => x"06",
          8677 => x"52",
          8678 => x"9e",
          8679 => x"52",
          8680 => x"ff",
          8681 => x"f0",
          8682 => x"1b",
          8683 => x"87",
          8684 => x"55",
          8685 => x"83",
          8686 => x"74",
          8687 => x"ff",
          8688 => x"7c",
          8689 => x"74",
          8690 => x"38",
          8691 => x"54",
          8692 => x"52",
          8693 => x"99",
          8694 => x"b5",
          8695 => x"87",
          8696 => x"53",
          8697 => x"08",
          8698 => x"ff",
          8699 => x"76",
          8700 => x"31",
          8701 => x"cd",
          8702 => x"58",
          8703 => x"ff",
          8704 => x"55",
          8705 => x"83",
          8706 => x"61",
          8707 => x"26",
          8708 => x"57",
          8709 => x"53",
          8710 => x"51",
          8711 => x"3f",
          8712 => x"08",
          8713 => x"76",
          8714 => x"31",
          8715 => x"db",
          8716 => x"7d",
          8717 => x"38",
          8718 => x"83",
          8719 => x"8a",
          8720 => x"7d",
          8721 => x"38",
          8722 => x"81",
          8723 => x"80",
          8724 => x"80",
          8725 => x"7a",
          8726 => x"bc",
          8727 => x"d5",
          8728 => x"ff",
          8729 => x"83",
          8730 => x"77",
          8731 => x"0b",
          8732 => x"81",
          8733 => x"34",
          8734 => x"34",
          8735 => x"34",
          8736 => x"56",
          8737 => x"52",
          8738 => x"c1",
          8739 => x"0b",
          8740 => x"82",
          8741 => x"82",
          8742 => x"56",
          8743 => x"34",
          8744 => x"08",
          8745 => x"60",
          8746 => x"1b",
          8747 => x"96",
          8748 => x"83",
          8749 => x"ff",
          8750 => x"81",
          8751 => x"7a",
          8752 => x"ff",
          8753 => x"81",
          8754 => x"a8",
          8755 => x"80",
          8756 => x"7e",
          8757 => x"e3",
          8758 => x"82",
          8759 => x"90",
          8760 => x"8e",
          8761 => x"81",
          8762 => x"82",
          8763 => x"56",
          8764 => x"a8",
          8765 => x"0d",
          8766 => x"0d",
          8767 => x"59",
          8768 => x"ff",
          8769 => x"57",
          8770 => x"b4",
          8771 => x"f8",
          8772 => x"81",
          8773 => x"52",
          8774 => x"dc",
          8775 => x"2e",
          8776 => x"9c",
          8777 => x"33",
          8778 => x"2e",
          8779 => x"76",
          8780 => x"58",
          8781 => x"57",
          8782 => x"09",
          8783 => x"38",
          8784 => x"78",
          8785 => x"38",
          8786 => x"82",
          8787 => x"8d",
          8788 => x"f7",
          8789 => x"02",
          8790 => x"05",
          8791 => x"77",
          8792 => x"81",
          8793 => x"8d",
          8794 => x"e7",
          8795 => x"08",
          8796 => x"24",
          8797 => x"17",
          8798 => x"8c",
          8799 => x"77",
          8800 => x"16",
          8801 => x"25",
          8802 => x"3d",
          8803 => x"75",
          8804 => x"52",
          8805 => x"cb",
          8806 => x"76",
          8807 => x"70",
          8808 => x"2a",
          8809 => x"51",
          8810 => x"84",
          8811 => x"19",
          8812 => x"8b",
          8813 => x"f9",
          8814 => x"84",
          8815 => x"56",
          8816 => x"a7",
          8817 => x"fc",
          8818 => x"53",
          8819 => x"75",
          8820 => x"a1",
          8821 => x"a8",
          8822 => x"84",
          8823 => x"2e",
          8824 => x"87",
          8825 => x"08",
          8826 => x"ff",
          8827 => x"b5",
          8828 => x"3d",
          8829 => x"3d",
          8830 => x"80",
          8831 => x"52",
          8832 => x"9a",
          8833 => x"74",
          8834 => x"0d",
          8835 => x"0d",
          8836 => x"05",
          8837 => x"86",
          8838 => x"54",
          8839 => x"73",
          8840 => x"fe",
          8841 => x"51",
          8842 => x"98",
          8843 => x"00",
          8844 => x"ff",
          8845 => x"00",
          8846 => x"ff",
          8847 => x"ff",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"69",
          8985 => x"00",
          8986 => x"69",
          8987 => x"6c",
          8988 => x"69",
          8989 => x"00",
          8990 => x"6c",
          8991 => x"00",
          8992 => x"65",
          8993 => x"00",
          8994 => x"63",
          8995 => x"72",
          8996 => x"63",
          8997 => x"00",
          8998 => x"64",
          8999 => x"00",
          9000 => x"64",
          9001 => x"00",
          9002 => x"65",
          9003 => x"65",
          9004 => x"65",
          9005 => x"69",
          9006 => x"69",
          9007 => x"66",
          9008 => x"66",
          9009 => x"61",
          9010 => x"00",
          9011 => x"6d",
          9012 => x"65",
          9013 => x"72",
          9014 => x"65",
          9015 => x"00",
          9016 => x"6e",
          9017 => x"00",
          9018 => x"65",
          9019 => x"00",
          9020 => x"62",
          9021 => x"63",
          9022 => x"62",
          9023 => x"63",
          9024 => x"69",
          9025 => x"00",
          9026 => x"64",
          9027 => x"69",
          9028 => x"45",
          9029 => x"72",
          9030 => x"6e",
          9031 => x"6e",
          9032 => x"65",
          9033 => x"72",
          9034 => x"00",
          9035 => x"69",
          9036 => x"6e",
          9037 => x"72",
          9038 => x"79",
          9039 => x"00",
          9040 => x"6f",
          9041 => x"6c",
          9042 => x"6f",
          9043 => x"2e",
          9044 => x"6f",
          9045 => x"74",
          9046 => x"6f",
          9047 => x"2e",
          9048 => x"6e",
          9049 => x"69",
          9050 => x"69",
          9051 => x"61",
          9052 => x"0a",
          9053 => x"63",
          9054 => x"73",
          9055 => x"6e",
          9056 => x"2e",
          9057 => x"69",
          9058 => x"61",
          9059 => x"61",
          9060 => x"65",
          9061 => x"74",
          9062 => x"00",
          9063 => x"69",
          9064 => x"68",
          9065 => x"6c",
          9066 => x"6e",
          9067 => x"69",
          9068 => x"00",
          9069 => x"44",
          9070 => x"20",
          9071 => x"74",
          9072 => x"72",
          9073 => x"63",
          9074 => x"2e",
          9075 => x"72",
          9076 => x"20",
          9077 => x"62",
          9078 => x"69",
          9079 => x"6e",
          9080 => x"69",
          9081 => x"00",
          9082 => x"69",
          9083 => x"6e",
          9084 => x"65",
          9085 => x"6c",
          9086 => x"0a",
          9087 => x"6f",
          9088 => x"6d",
          9089 => x"69",
          9090 => x"20",
          9091 => x"65",
          9092 => x"74",
          9093 => x"66",
          9094 => x"64",
          9095 => x"20",
          9096 => x"6b",
          9097 => x"00",
          9098 => x"6f",
          9099 => x"74",
          9100 => x"6f",
          9101 => x"64",
          9102 => x"00",
          9103 => x"69",
          9104 => x"75",
          9105 => x"6f",
          9106 => x"61",
          9107 => x"6e",
          9108 => x"6e",
          9109 => x"6c",
          9110 => x"0a",
          9111 => x"69",
          9112 => x"69",
          9113 => x"6f",
          9114 => x"64",
          9115 => x"00",
          9116 => x"6e",
          9117 => x"66",
          9118 => x"65",
          9119 => x"6d",
          9120 => x"72",
          9121 => x"00",
          9122 => x"6f",
          9123 => x"61",
          9124 => x"6f",
          9125 => x"20",
          9126 => x"65",
          9127 => x"00",
          9128 => x"61",
          9129 => x"65",
          9130 => x"73",
          9131 => x"63",
          9132 => x"65",
          9133 => x"0a",
          9134 => x"75",
          9135 => x"73",
          9136 => x"00",
          9137 => x"6e",
          9138 => x"77",
          9139 => x"72",
          9140 => x"2e",
          9141 => x"25",
          9142 => x"62",
          9143 => x"73",
          9144 => x"20",
          9145 => x"25",
          9146 => x"62",
          9147 => x"73",
          9148 => x"63",
          9149 => x"00",
          9150 => x"65",
          9151 => x"00",
          9152 => x"30",
          9153 => x"00",
          9154 => x"20",
          9155 => x"30",
          9156 => x"00",
          9157 => x"20",
          9158 => x"20",
          9159 => x"00",
          9160 => x"30",
          9161 => x"00",
          9162 => x"20",
          9163 => x"7c",
          9164 => x"0d",
          9165 => x"4f",
          9166 => x"2a",
          9167 => x"73",
          9168 => x"00",
          9169 => x"32",
          9170 => x"2f",
          9171 => x"30",
          9172 => x"31",
          9173 => x"00",
          9174 => x"5a",
          9175 => x"20",
          9176 => x"20",
          9177 => x"78",
          9178 => x"73",
          9179 => x"20",
          9180 => x"0a",
          9181 => x"50",
          9182 => x"6e",
          9183 => x"72",
          9184 => x"20",
          9185 => x"64",
          9186 => x"0a",
          9187 => x"69",
          9188 => x"20",
          9189 => x"65",
          9190 => x"70",
          9191 => x"00",
          9192 => x"53",
          9193 => x"6e",
          9194 => x"72",
          9195 => x"0a",
          9196 => x"4f",
          9197 => x"20",
          9198 => x"69",
          9199 => x"72",
          9200 => x"74",
          9201 => x"4f",
          9202 => x"20",
          9203 => x"69",
          9204 => x"72",
          9205 => x"74",
          9206 => x"41",
          9207 => x"20",
          9208 => x"69",
          9209 => x"72",
          9210 => x"74",
          9211 => x"41",
          9212 => x"20",
          9213 => x"69",
          9214 => x"72",
          9215 => x"74",
          9216 => x"41",
          9217 => x"20",
          9218 => x"69",
          9219 => x"72",
          9220 => x"74",
          9221 => x"41",
          9222 => x"20",
          9223 => x"69",
          9224 => x"72",
          9225 => x"74",
          9226 => x"65",
          9227 => x"6e",
          9228 => x"70",
          9229 => x"6d",
          9230 => x"2e",
          9231 => x"00",
          9232 => x"6e",
          9233 => x"69",
          9234 => x"74",
          9235 => x"72",
          9236 => x"0a",
          9237 => x"75",
          9238 => x"78",
          9239 => x"62",
          9240 => x"00",
          9241 => x"4f",
          9242 => x"73",
          9243 => x"3a",
          9244 => x"61",
          9245 => x"64",
          9246 => x"20",
          9247 => x"74",
          9248 => x"69",
          9249 => x"73",
          9250 => x"61",
          9251 => x"30",
          9252 => x"6c",
          9253 => x"65",
          9254 => x"69",
          9255 => x"61",
          9256 => x"6c",
          9257 => x"00",
          9258 => x"20",
          9259 => x"6c",
          9260 => x"69",
          9261 => x"2e",
          9262 => x"00",
          9263 => x"6f",
          9264 => x"6e",
          9265 => x"2e",
          9266 => x"6f",
          9267 => x"72",
          9268 => x"2e",
          9269 => x"00",
          9270 => x"30",
          9271 => x"28",
          9272 => x"78",
          9273 => x"25",
          9274 => x"78",
          9275 => x"38",
          9276 => x"00",
          9277 => x"75",
          9278 => x"4d",
          9279 => x"72",
          9280 => x"00",
          9281 => x"43",
          9282 => x"6c",
          9283 => x"2e",
          9284 => x"30",
          9285 => x"25",
          9286 => x"2d",
          9287 => x"3f",
          9288 => x"00",
          9289 => x"30",
          9290 => x"25",
          9291 => x"2d",
          9292 => x"30",
          9293 => x"25",
          9294 => x"2d",
          9295 => x"78",
          9296 => x"74",
          9297 => x"20",
          9298 => x"65",
          9299 => x"25",
          9300 => x"20",
          9301 => x"0a",
          9302 => x"61",
          9303 => x"6e",
          9304 => x"6f",
          9305 => x"40",
          9306 => x"38",
          9307 => x"2e",
          9308 => x"00",
          9309 => x"61",
          9310 => x"72",
          9311 => x"72",
          9312 => x"20",
          9313 => x"65",
          9314 => x"64",
          9315 => x"00",
          9316 => x"65",
          9317 => x"72",
          9318 => x"67",
          9319 => x"70",
          9320 => x"61",
          9321 => x"6e",
          9322 => x"0a",
          9323 => x"6f",
          9324 => x"72",
          9325 => x"6f",
          9326 => x"67",
          9327 => x"0a",
          9328 => x"50",
          9329 => x"69",
          9330 => x"64",
          9331 => x"73",
          9332 => x"2e",
          9333 => x"00",
          9334 => x"64",
          9335 => x"73",
          9336 => x"00",
          9337 => x"64",
          9338 => x"73",
          9339 => x"61",
          9340 => x"6f",
          9341 => x"6e",
          9342 => x"00",
          9343 => x"45",
          9344 => x"20",
          9345 => x"52",
          9346 => x"50",
          9347 => x"54",
          9348 => x"45",
          9349 => x"20",
          9350 => x"52",
          9351 => x"50",
          9352 => x"54",
          9353 => x"75",
          9354 => x"6e",
          9355 => x"2e",
          9356 => x"6e",
          9357 => x"69",
          9358 => x"69",
          9359 => x"72",
          9360 => x"74",
          9361 => x"2e",
          9362 => x"64",
          9363 => x"2f",
          9364 => x"25",
          9365 => x"64",
          9366 => x"2e",
          9367 => x"64",
          9368 => x"6f",
          9369 => x"6f",
          9370 => x"67",
          9371 => x"74",
          9372 => x"00",
          9373 => x"28",
          9374 => x"6d",
          9375 => x"43",
          9376 => x"6e",
          9377 => x"29",
          9378 => x"0a",
          9379 => x"69",
          9380 => x"20",
          9381 => x"6c",
          9382 => x"6e",
          9383 => x"3a",
          9384 => x"20",
          9385 => x"42",
          9386 => x"52",
          9387 => x"20",
          9388 => x"38",
          9389 => x"30",
          9390 => x"2e",
          9391 => x"20",
          9392 => x"44",
          9393 => x"20",
          9394 => x"20",
          9395 => x"38",
          9396 => x"30",
          9397 => x"2e",
          9398 => x"20",
          9399 => x"4e",
          9400 => x"42",
          9401 => x"20",
          9402 => x"38",
          9403 => x"30",
          9404 => x"2e",
          9405 => x"20",
          9406 => x"52",
          9407 => x"20",
          9408 => x"20",
          9409 => x"38",
          9410 => x"30",
          9411 => x"2e",
          9412 => x"20",
          9413 => x"41",
          9414 => x"20",
          9415 => x"20",
          9416 => x"38",
          9417 => x"30",
          9418 => x"2e",
          9419 => x"20",
          9420 => x"44",
          9421 => x"52",
          9422 => x"20",
          9423 => x"76",
          9424 => x"73",
          9425 => x"30",
          9426 => x"2e",
          9427 => x"20",
          9428 => x"49",
          9429 => x"31",
          9430 => x"20",
          9431 => x"6d",
          9432 => x"20",
          9433 => x"30",
          9434 => x"2e",
          9435 => x"20",
          9436 => x"4e",
          9437 => x"43",
          9438 => x"20",
          9439 => x"61",
          9440 => x"6c",
          9441 => x"30",
          9442 => x"2e",
          9443 => x"20",
          9444 => x"49",
          9445 => x"4f",
          9446 => x"42",
          9447 => x"00",
          9448 => x"20",
          9449 => x"42",
          9450 => x"43",
          9451 => x"20",
          9452 => x"4f",
          9453 => x"0a",
          9454 => x"20",
          9455 => x"53",
          9456 => x"00",
          9457 => x"20",
          9458 => x"50",
          9459 => x"00",
          9460 => x"64",
          9461 => x"73",
          9462 => x"3a",
          9463 => x"20",
          9464 => x"50",
          9465 => x"65",
          9466 => x"20",
          9467 => x"74",
          9468 => x"41",
          9469 => x"65",
          9470 => x"3d",
          9471 => x"38",
          9472 => x"00",
          9473 => x"20",
          9474 => x"50",
          9475 => x"65",
          9476 => x"79",
          9477 => x"61",
          9478 => x"41",
          9479 => x"65",
          9480 => x"3d",
          9481 => x"38",
          9482 => x"00",
          9483 => x"20",
          9484 => x"74",
          9485 => x"20",
          9486 => x"72",
          9487 => x"64",
          9488 => x"73",
          9489 => x"20",
          9490 => x"3d",
          9491 => x"38",
          9492 => x"00",
          9493 => x"69",
          9494 => x"0a",
          9495 => x"20",
          9496 => x"50",
          9497 => x"64",
          9498 => x"20",
          9499 => x"20",
          9500 => x"20",
          9501 => x"20",
          9502 => x"3d",
          9503 => x"34",
          9504 => x"00",
          9505 => x"20",
          9506 => x"79",
          9507 => x"6d",
          9508 => x"6f",
          9509 => x"46",
          9510 => x"20",
          9511 => x"20",
          9512 => x"3d",
          9513 => x"2e",
          9514 => x"64",
          9515 => x"0a",
          9516 => x"20",
          9517 => x"44",
          9518 => x"20",
          9519 => x"63",
          9520 => x"72",
          9521 => x"20",
          9522 => x"20",
          9523 => x"3d",
          9524 => x"2e",
          9525 => x"64",
          9526 => x"0a",
          9527 => x"20",
          9528 => x"69",
          9529 => x"6f",
          9530 => x"53",
          9531 => x"4d",
          9532 => x"6f",
          9533 => x"46",
          9534 => x"3d",
          9535 => x"2e",
          9536 => x"64",
          9537 => x"0a",
          9538 => x"6d",
          9539 => x"00",
          9540 => x"65",
          9541 => x"6d",
          9542 => x"6c",
          9543 => x"00",
          9544 => x"56",
          9545 => x"56",
          9546 => x"6e",
          9547 => x"6e",
          9548 => x"77",
          9549 => x"00",
          9550 => x"00",
          9551 => x"00",
          9552 => x"00",
          9553 => x"00",
          9554 => x"00",
          9555 => x"00",
          9556 => x"00",
          9557 => x"00",
          9558 => x"00",
          9559 => x"00",
          9560 => x"00",
          9561 => x"00",
          9562 => x"00",
          9563 => x"00",
          9564 => x"00",
          9565 => x"00",
          9566 => x"00",
          9567 => x"00",
          9568 => x"00",
          9569 => x"00",
          9570 => x"00",
          9571 => x"00",
          9572 => x"00",
          9573 => x"00",
          9574 => x"00",
          9575 => x"00",
          9576 => x"00",
          9577 => x"00",
          9578 => x"00",
          9579 => x"00",
          9580 => x"00",
          9581 => x"00",
          9582 => x"00",
          9583 => x"00",
          9584 => x"00",
          9585 => x"00",
          9586 => x"00",
          9587 => x"00",
          9588 => x"00",
          9589 => x"00",
          9590 => x"00",
          9591 => x"00",
          9592 => x"00",
          9593 => x"00",
          9594 => x"00",
          9595 => x"00",
          9596 => x"00",
          9597 => x"00",
          9598 => x"00",
          9599 => x"00",
          9600 => x"00",
          9601 => x"00",
          9602 => x"00",
          9603 => x"00",
          9604 => x"00",
          9605 => x"00",
          9606 => x"00",
          9607 => x"00",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"5b",
          9616 => x"5b",
          9617 => x"5b",
          9618 => x"5b",
          9619 => x"5b",
          9620 => x"5b",
          9621 => x"5b",
          9622 => x"30",
          9623 => x"5b",
          9624 => x"5b",
          9625 => x"5b",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"69",
          9638 => x"72",
          9639 => x"69",
          9640 => x"00",
          9641 => x"00",
          9642 => x"30",
          9643 => x"20",
          9644 => x"00",
          9645 => x"61",
          9646 => x"64",
          9647 => x"20",
          9648 => x"65",
          9649 => x"68",
          9650 => x"69",
          9651 => x"72",
          9652 => x"69",
          9653 => x"74",
          9654 => x"4f",
          9655 => x"00",
          9656 => x"61",
          9657 => x"74",
          9658 => x"65",
          9659 => x"72",
          9660 => x"65",
          9661 => x"73",
          9662 => x"79",
          9663 => x"6c",
          9664 => x"64",
          9665 => x"62",
          9666 => x"67",
          9667 => x"44",
          9668 => x"2a",
          9669 => x"3b",
          9670 => x"3f",
          9671 => x"7f",
          9672 => x"41",
          9673 => x"41",
          9674 => x"00",
          9675 => x"fe",
          9676 => x"44",
          9677 => x"2e",
          9678 => x"4f",
          9679 => x"4d",
          9680 => x"20",
          9681 => x"54",
          9682 => x"20",
          9683 => x"4f",
          9684 => x"4d",
          9685 => x"20",
          9686 => x"54",
          9687 => x"20",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"9a",
          9693 => x"41",
          9694 => x"45",
          9695 => x"49",
          9696 => x"92",
          9697 => x"4f",
          9698 => x"99",
          9699 => x"9d",
          9700 => x"49",
          9701 => x"a5",
          9702 => x"a9",
          9703 => x"ad",
          9704 => x"b1",
          9705 => x"b5",
          9706 => x"b9",
          9707 => x"bd",
          9708 => x"c1",
          9709 => x"c5",
          9710 => x"c9",
          9711 => x"cd",
          9712 => x"d1",
          9713 => x"d5",
          9714 => x"d9",
          9715 => x"dd",
          9716 => x"e1",
          9717 => x"e5",
          9718 => x"e9",
          9719 => x"ed",
          9720 => x"f1",
          9721 => x"f5",
          9722 => x"f9",
          9723 => x"fd",
          9724 => x"2e",
          9725 => x"5b",
          9726 => x"22",
          9727 => x"3e",
          9728 => x"00",
          9729 => x"01",
          9730 => x"10",
          9731 => x"00",
          9732 => x"00",
          9733 => x"01",
          9734 => x"04",
          9735 => x"10",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"02",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"04",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"14",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"2b",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"30",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"3c",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"3d",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"3f",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"40",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"41",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"42",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"43",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"50",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"51",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"54",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"55",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"79",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"78",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"82",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"83",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"85",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"87",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"8c",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"8d",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"8e",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"8f",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"00",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"01",
          9848 => x"00",
          9849 => x"01",
          9850 => x"81",
          9851 => x"00",
          9852 => x"7f",
          9853 => x"00",
          9854 => x"00",
          9855 => x"00",
          9856 => x"00",
          9857 => x"f5",
          9858 => x"f5",
          9859 => x"f5",
          9860 => x"00",
          9861 => x"01",
          9862 => x"01",
          9863 => x"01",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"00",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"00",
          9891 => x"00",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9b",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"b0",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"94",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"80",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"ef",
           278 => x"0b",
           279 => x"0b",
           280 => x"8d",
           281 => x"0b",
           282 => x"0b",
           283 => x"ab",
           284 => x"0b",
           285 => x"0b",
           286 => x"cb",
           287 => x"0b",
           288 => x"0b",
           289 => x"eb",
           290 => x"0b",
           291 => x"0b",
           292 => x"8b",
           293 => x"0b",
           294 => x"0b",
           295 => x"ab",
           296 => x"0b",
           297 => x"0b",
           298 => x"cb",
           299 => x"0b",
           300 => x"0b",
           301 => x"eb",
           302 => x"0b",
           303 => x"0b",
           304 => x"8b",
           305 => x"0b",
           306 => x"0b",
           307 => x"ab",
           308 => x"0b",
           309 => x"0b",
           310 => x"cb",
           311 => x"0b",
           312 => x"0b",
           313 => x"eb",
           314 => x"0b",
           315 => x"0b",
           316 => x"8b",
           317 => x"0b",
           318 => x"0b",
           319 => x"ab",
           320 => x"0b",
           321 => x"0b",
           322 => x"cb",
           323 => x"0b",
           324 => x"0b",
           325 => x"eb",
           326 => x"0b",
           327 => x"0b",
           328 => x"8b",
           329 => x"0b",
           330 => x"0b",
           331 => x"ab",
           332 => x"0b",
           333 => x"0b",
           334 => x"cb",
           335 => x"0b",
           336 => x"0b",
           337 => x"eb",
           338 => x"0b",
           339 => x"0b",
           340 => x"8b",
           341 => x"0b",
           342 => x"0b",
           343 => x"ab",
           344 => x"0b",
           345 => x"0b",
           346 => x"cb",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"bb",
           395 => x"b5",
           396 => x"d0",
           397 => x"b5",
           398 => x"fc",
           399 => x"b4",
           400 => x"90",
           401 => x"b4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"82",
           408 => x"82",
           409 => x"b5",
           410 => x"b5",
           411 => x"d0",
           412 => x"b5",
           413 => x"ab",
           414 => x"b4",
           415 => x"90",
           416 => x"b4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"82",
           423 => x"82",
           424 => x"97",
           425 => x"b5",
           426 => x"d0",
           427 => x"b5",
           428 => x"f7",
           429 => x"b5",
           430 => x"d0",
           431 => x"b5",
           432 => x"f8",
           433 => x"b5",
           434 => x"d0",
           435 => x"b5",
           436 => x"f0",
           437 => x"b5",
           438 => x"d0",
           439 => x"b5",
           440 => x"f2",
           441 => x"b5",
           442 => x"d0",
           443 => x"b5",
           444 => x"f3",
           445 => x"b5",
           446 => x"d0",
           447 => x"b5",
           448 => x"d7",
           449 => x"b5",
           450 => x"d0",
           451 => x"b5",
           452 => x"e4",
           453 => x"b5",
           454 => x"d0",
           455 => x"b5",
           456 => x"db",
           457 => x"b5",
           458 => x"d0",
           459 => x"b5",
           460 => x"de",
           461 => x"b5",
           462 => x"d0",
           463 => x"b5",
           464 => x"e9",
           465 => x"b5",
           466 => x"d0",
           467 => x"b5",
           468 => x"f1",
           469 => x"b5",
           470 => x"d0",
           471 => x"b5",
           472 => x"e2",
           473 => x"b5",
           474 => x"d0",
           475 => x"b5",
           476 => x"ec",
           477 => x"b5",
           478 => x"d0",
           479 => x"b5",
           480 => x"ed",
           481 => x"b5",
           482 => x"d0",
           483 => x"b5",
           484 => x"ed",
           485 => x"b5",
           486 => x"d0",
           487 => x"b5",
           488 => x"f5",
           489 => x"b5",
           490 => x"d0",
           491 => x"b5",
           492 => x"f3",
           493 => x"b5",
           494 => x"d0",
           495 => x"b5",
           496 => x"f8",
           497 => x"b5",
           498 => x"d0",
           499 => x"b5",
           500 => x"ee",
           501 => x"b5",
           502 => x"d0",
           503 => x"b5",
           504 => x"fb",
           505 => x"b5",
           506 => x"d0",
           507 => x"b5",
           508 => x"fc",
           509 => x"b5",
           510 => x"d0",
           511 => x"b5",
           512 => x"e4",
           513 => x"b5",
           514 => x"d0",
           515 => x"b5",
           516 => x"e4",
           517 => x"b5",
           518 => x"d0",
           519 => x"b5",
           520 => x"e5",
           521 => x"b5",
           522 => x"d0",
           523 => x"b5",
           524 => x"ef",
           525 => x"b5",
           526 => x"d0",
           527 => x"b5",
           528 => x"fd",
           529 => x"b5",
           530 => x"d0",
           531 => x"b5",
           532 => x"ff",
           533 => x"b5",
           534 => x"d0",
           535 => x"b5",
           536 => x"82",
           537 => x"b5",
           538 => x"d0",
           539 => x"b5",
           540 => x"d6",
           541 => x"b5",
           542 => x"d0",
           543 => x"b5",
           544 => x"85",
           545 => x"b5",
           546 => x"d0",
           547 => x"b5",
           548 => x"94",
           549 => x"b5",
           550 => x"d0",
           551 => x"b5",
           552 => x"91",
           553 => x"b5",
           554 => x"d0",
           555 => x"b5",
           556 => x"a7",
           557 => x"b5",
           558 => x"d0",
           559 => x"b5",
           560 => x"a9",
           561 => x"b5",
           562 => x"d0",
           563 => x"b5",
           564 => x"ab",
           565 => x"b5",
           566 => x"d0",
           567 => x"b5",
           568 => x"f0",
           569 => x"b5",
           570 => x"d0",
           571 => x"b5",
           572 => x"f1",
           573 => x"b5",
           574 => x"d0",
           575 => x"b5",
           576 => x"f5",
           577 => x"b5",
           578 => x"d0",
           579 => x"b5",
           580 => x"d6",
           581 => x"b5",
           582 => x"d0",
           583 => x"b5",
           584 => x"a1",
           585 => x"b5",
           586 => x"d0",
           587 => x"b5",
           588 => x"a2",
           589 => x"b5",
           590 => x"d0",
           591 => x"b5",
           592 => x"a6",
           593 => x"b5",
           594 => x"d0",
           595 => x"b5",
           596 => x"9e",
           597 => x"b5",
           598 => x"d0",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"b5",
           623 => x"cd",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"ba",
           628 => x"51",
           629 => x"04",
           630 => x"b4",
           631 => x"b5",
           632 => x"3d",
           633 => x"b4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"b4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"b4",
           651 => x"b5",
           652 => x"82",
           653 => x"fb",
           654 => x"b5",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"b4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"b4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"b5",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"ab",
           685 => x"b5",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"b4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"b4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"b4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"b5",
           712 => x"05",
           713 => x"b5",
           714 => x"05",
           715 => x"b5",
           716 => x"05",
           717 => x"a8",
           718 => x"0d",
           719 => x"0c",
           720 => x"b4",
           721 => x"b5",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"b5",
           726 => x"05",
           727 => x"b4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"b5",
           732 => x"05",
           733 => x"b4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"a8",
           743 => x"b5",
           744 => x"05",
           745 => x"b4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"b4",
           751 => x"08",
           752 => x"a8",
           753 => x"3d",
           754 => x"b4",
           755 => x"b5",
           756 => x"82",
           757 => x"fb",
           758 => x"b5",
           759 => x"05",
           760 => x"b4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"b4",
           778 => x"b5",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"b5",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"b5",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"b5",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"b5",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"b5",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"b4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"b4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"b4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"b5",
           848 => x"05",
           849 => x"b4",
           850 => x"33",
           851 => x"b4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"b5",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"b5",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"b4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"b5",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"b5",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"95",
           901 => x"08",
           902 => x"53",
           903 => x"b5",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"b5",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"b4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"b4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"b4",
           927 => x"22",
           928 => x"51",
           929 => x"b5",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"b4",
           935 => x"22",
           936 => x"51",
           937 => x"b5",
           938 => x"05",
           939 => x"39",
           940 => x"b5",
           941 => x"05",
           942 => x"b4",
           943 => x"22",
           944 => x"53",
           945 => x"b4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"b4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"b4",
           955 => x"0c",
           956 => x"53",
           957 => x"b4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"b5",
           965 => x"05",
           966 => x"b4",
           967 => x"08",
           968 => x"b5",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"b5",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"b4",
           987 => x"23",
           988 => x"b5",
           989 => x"05",
           990 => x"ac",
           991 => x"a8",
           992 => x"82",
           993 => x"f4",
           994 => x"b5",
           995 => x"05",
           996 => x"b5",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"b4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"b4",
          1007 => x"0c",
          1008 => x"b5",
          1009 => x"05",
          1010 => x"b4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"b5",
          1020 => x"05",
          1021 => x"ac",
          1022 => x"b5",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"b4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"b5",
          1031 => x"05",
          1032 => x"b4",
          1033 => x"22",
          1034 => x"b4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"b5",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"b4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"b4",
          1050 => x"0c",
          1051 => x"b5",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"b4",
          1061 => x"0c",
          1062 => x"b4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"b5",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"b5",
          1074 => x"05",
          1075 => x"b5",
          1076 => x"05",
          1077 => x"b4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"b5",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"b4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"b4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"b4",
          1106 => x"0c",
          1107 => x"b5",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"b4",
          1117 => x"0c",
          1118 => x"b4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"b5",
          1130 => x"05",
          1131 => x"b4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"95",
          1137 => x"a8",
          1138 => x"75",
          1139 => x"b4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"b5",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"b4",
          1154 => x"34",
          1155 => x"b5",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"b4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"b4",
          1166 => x"08",
          1167 => x"b5",
          1168 => x"05",
          1169 => x"b4",
          1170 => x"22",
          1171 => x"b5",
          1172 => x"05",
          1173 => x"ad",
          1174 => x"b5",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"b4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"b5",
          1187 => x"05",
          1188 => x"b4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"b5",
          1193 => x"05",
          1194 => x"51",
          1195 => x"b5",
          1196 => x"05",
          1197 => x"b4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"b4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"b4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"b4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"b4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"b5",
          1227 => x"05",
          1228 => x"b4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"b4",
          1245 => x"23",
          1246 => x"b5",
          1247 => x"05",
          1248 => x"b5",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"b5",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"b4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"b5",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"b4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"b5",
          1281 => x"05",
          1282 => x"b4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"b4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"b4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"b4",
          1295 => x"08",
          1296 => x"96",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"b4",
          1304 => x"08",
          1305 => x"95",
          1306 => x"c7",
          1307 => x"b4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"b5",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"b4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"b5",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"81",
          1333 => x"b4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"b4",
          1338 => x"08",
          1339 => x"b4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"b4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"b4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"b4",
          1356 => x"08",
          1357 => x"94",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"b4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"b4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"b4",
          1373 => x"08",
          1374 => x"93",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"b5",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"92",
          1401 => x"ee",
          1402 => x"b4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"b5",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"92",
          1424 => x"b7",
          1425 => x"b4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"91",
          1443 => x"b5",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"b4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"b5",
          1452 => x"05",
          1453 => x"b5",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"b5",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"b5",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"bd",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"90",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"b5",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"b4",
          1494 => x"23",
          1495 => x"b5",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"b4",
          1501 => x"08",
          1502 => x"b4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"b5",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"b5",
          1513 => x"3d",
          1514 => x"b4",
          1515 => x"b5",
          1516 => x"82",
          1517 => x"f7",
          1518 => x"0b",
          1519 => x"08",
          1520 => x"82",
          1521 => x"8c",
          1522 => x"80",
          1523 => x"b5",
          1524 => x"05",
          1525 => x"51",
          1526 => x"53",
          1527 => x"b4",
          1528 => x"34",
          1529 => x"06",
          1530 => x"2e",
          1531 => x"91",
          1532 => x"b4",
          1533 => x"08",
          1534 => x"05",
          1535 => x"ce",
          1536 => x"b4",
          1537 => x"33",
          1538 => x"2e",
          1539 => x"a4",
          1540 => x"82",
          1541 => x"f0",
          1542 => x"b5",
          1543 => x"05",
          1544 => x"81",
          1545 => x"70",
          1546 => x"72",
          1547 => x"b4",
          1548 => x"34",
          1549 => x"08",
          1550 => x"53",
          1551 => x"09",
          1552 => x"dc",
          1553 => x"b4",
          1554 => x"08",
          1555 => x"05",
          1556 => x"08",
          1557 => x"33",
          1558 => x"08",
          1559 => x"82",
          1560 => x"f8",
          1561 => x"b5",
          1562 => x"05",
          1563 => x"b4",
          1564 => x"08",
          1565 => x"b6",
          1566 => x"b4",
          1567 => x"08",
          1568 => x"84",
          1569 => x"39",
          1570 => x"b5",
          1571 => x"05",
          1572 => x"b4",
          1573 => x"08",
          1574 => x"05",
          1575 => x"08",
          1576 => x"33",
          1577 => x"08",
          1578 => x"81",
          1579 => x"0b",
          1580 => x"08",
          1581 => x"82",
          1582 => x"88",
          1583 => x"08",
          1584 => x"0c",
          1585 => x"53",
          1586 => x"b5",
          1587 => x"05",
          1588 => x"39",
          1589 => x"08",
          1590 => x"53",
          1591 => x"8d",
          1592 => x"82",
          1593 => x"ec",
          1594 => x"80",
          1595 => x"b4",
          1596 => x"33",
          1597 => x"27",
          1598 => x"b5",
          1599 => x"05",
          1600 => x"b9",
          1601 => x"8d",
          1602 => x"82",
          1603 => x"ec",
          1604 => x"d8",
          1605 => x"82",
          1606 => x"f4",
          1607 => x"39",
          1608 => x"08",
          1609 => x"53",
          1610 => x"90",
          1611 => x"b4",
          1612 => x"33",
          1613 => x"26",
          1614 => x"39",
          1615 => x"b5",
          1616 => x"05",
          1617 => x"39",
          1618 => x"b5",
          1619 => x"05",
          1620 => x"82",
          1621 => x"fc",
          1622 => x"b5",
          1623 => x"05",
          1624 => x"73",
          1625 => x"38",
          1626 => x"08",
          1627 => x"53",
          1628 => x"27",
          1629 => x"b5",
          1630 => x"05",
          1631 => x"51",
          1632 => x"b5",
          1633 => x"05",
          1634 => x"b4",
          1635 => x"33",
          1636 => x"53",
          1637 => x"b4",
          1638 => x"34",
          1639 => x"08",
          1640 => x"53",
          1641 => x"ad",
          1642 => x"b4",
          1643 => x"33",
          1644 => x"53",
          1645 => x"b4",
          1646 => x"34",
          1647 => x"08",
          1648 => x"53",
          1649 => x"8d",
          1650 => x"82",
          1651 => x"ec",
          1652 => x"98",
          1653 => x"b4",
          1654 => x"33",
          1655 => x"08",
          1656 => x"54",
          1657 => x"26",
          1658 => x"0b",
          1659 => x"08",
          1660 => x"80",
          1661 => x"b5",
          1662 => x"05",
          1663 => x"b5",
          1664 => x"05",
          1665 => x"b5",
          1666 => x"05",
          1667 => x"82",
          1668 => x"fc",
          1669 => x"b5",
          1670 => x"05",
          1671 => x"81",
          1672 => x"70",
          1673 => x"52",
          1674 => x"33",
          1675 => x"08",
          1676 => x"fe",
          1677 => x"b5",
          1678 => x"05",
          1679 => x"80",
          1680 => x"82",
          1681 => x"fc",
          1682 => x"82",
          1683 => x"fc",
          1684 => x"b5",
          1685 => x"05",
          1686 => x"b4",
          1687 => x"08",
          1688 => x"81",
          1689 => x"b4",
          1690 => x"0c",
          1691 => x"08",
          1692 => x"82",
          1693 => x"8b",
          1694 => x"b5",
          1695 => x"82",
          1696 => x"02",
          1697 => x"0c",
          1698 => x"82",
          1699 => x"53",
          1700 => x"08",
          1701 => x"52",
          1702 => x"08",
          1703 => x"51",
          1704 => x"82",
          1705 => x"70",
          1706 => x"0c",
          1707 => x"0d",
          1708 => x"0c",
          1709 => x"b4",
          1710 => x"b5",
          1711 => x"3d",
          1712 => x"82",
          1713 => x"f0",
          1714 => x"b5",
          1715 => x"05",
          1716 => x"73",
          1717 => x"b4",
          1718 => x"08",
          1719 => x"53",
          1720 => x"72",
          1721 => x"08",
          1722 => x"72",
          1723 => x"53",
          1724 => x"09",
          1725 => x"38",
          1726 => x"08",
          1727 => x"70",
          1728 => x"71",
          1729 => x"39",
          1730 => x"08",
          1731 => x"53",
          1732 => x"09",
          1733 => x"38",
          1734 => x"b5",
          1735 => x"05",
          1736 => x"b4",
          1737 => x"08",
          1738 => x"05",
          1739 => x"08",
          1740 => x"33",
          1741 => x"08",
          1742 => x"82",
          1743 => x"f8",
          1744 => x"72",
          1745 => x"81",
          1746 => x"38",
          1747 => x"08",
          1748 => x"70",
          1749 => x"71",
          1750 => x"51",
          1751 => x"82",
          1752 => x"f8",
          1753 => x"b5",
          1754 => x"05",
          1755 => x"b4",
          1756 => x"0c",
          1757 => x"08",
          1758 => x"80",
          1759 => x"38",
          1760 => x"08",
          1761 => x"80",
          1762 => x"38",
          1763 => x"90",
          1764 => x"b4",
          1765 => x"34",
          1766 => x"08",
          1767 => x"70",
          1768 => x"71",
          1769 => x"51",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"a4",
          1773 => x"82",
          1774 => x"f4",
          1775 => x"b5",
          1776 => x"05",
          1777 => x"81",
          1778 => x"70",
          1779 => x"72",
          1780 => x"b4",
          1781 => x"34",
          1782 => x"82",
          1783 => x"f8",
          1784 => x"72",
          1785 => x"38",
          1786 => x"b5",
          1787 => x"05",
          1788 => x"39",
          1789 => x"08",
          1790 => x"53",
          1791 => x"90",
          1792 => x"b4",
          1793 => x"33",
          1794 => x"26",
          1795 => x"39",
          1796 => x"b5",
          1797 => x"05",
          1798 => x"39",
          1799 => x"b5",
          1800 => x"05",
          1801 => x"82",
          1802 => x"f8",
          1803 => x"af",
          1804 => x"38",
          1805 => x"08",
          1806 => x"53",
          1807 => x"83",
          1808 => x"80",
          1809 => x"b4",
          1810 => x"0c",
          1811 => x"8a",
          1812 => x"b4",
          1813 => x"34",
          1814 => x"b5",
          1815 => x"05",
          1816 => x"b4",
          1817 => x"33",
          1818 => x"27",
          1819 => x"82",
          1820 => x"f8",
          1821 => x"80",
          1822 => x"94",
          1823 => x"b4",
          1824 => x"33",
          1825 => x"53",
          1826 => x"b4",
          1827 => x"34",
          1828 => x"08",
          1829 => x"d0",
          1830 => x"72",
          1831 => x"08",
          1832 => x"82",
          1833 => x"f8",
          1834 => x"90",
          1835 => x"38",
          1836 => x"08",
          1837 => x"f9",
          1838 => x"72",
          1839 => x"08",
          1840 => x"82",
          1841 => x"f8",
          1842 => x"72",
          1843 => x"38",
          1844 => x"b5",
          1845 => x"05",
          1846 => x"39",
          1847 => x"08",
          1848 => x"82",
          1849 => x"f4",
          1850 => x"54",
          1851 => x"8d",
          1852 => x"82",
          1853 => x"ec",
          1854 => x"f7",
          1855 => x"b4",
          1856 => x"33",
          1857 => x"b4",
          1858 => x"08",
          1859 => x"b4",
          1860 => x"33",
          1861 => x"b5",
          1862 => x"05",
          1863 => x"b4",
          1864 => x"08",
          1865 => x"05",
          1866 => x"08",
          1867 => x"55",
          1868 => x"82",
          1869 => x"f8",
          1870 => x"a5",
          1871 => x"b4",
          1872 => x"33",
          1873 => x"2e",
          1874 => x"b5",
          1875 => x"05",
          1876 => x"b5",
          1877 => x"05",
          1878 => x"b4",
          1879 => x"08",
          1880 => x"08",
          1881 => x"71",
          1882 => x"0b",
          1883 => x"08",
          1884 => x"82",
          1885 => x"ec",
          1886 => x"b5",
          1887 => x"3d",
          1888 => x"b4",
          1889 => x"b5",
          1890 => x"82",
          1891 => x"fb",
          1892 => x"0b",
          1893 => x"08",
          1894 => x"82",
          1895 => x"85",
          1896 => x"81",
          1897 => x"32",
          1898 => x"51",
          1899 => x"53",
          1900 => x"8d",
          1901 => x"82",
          1902 => x"f4",
          1903 => x"92",
          1904 => x"b4",
          1905 => x"08",
          1906 => x"82",
          1907 => x"88",
          1908 => x"05",
          1909 => x"08",
          1910 => x"53",
          1911 => x"b4",
          1912 => x"34",
          1913 => x"06",
          1914 => x"2e",
          1915 => x"cc",
          1916 => x"cc",
          1917 => x"82",
          1918 => x"fc",
          1919 => x"90",
          1920 => x"53",
          1921 => x"b5",
          1922 => x"72",
          1923 => x"b1",
          1924 => x"82",
          1925 => x"f8",
          1926 => x"a5",
          1927 => x"fc",
          1928 => x"fc",
          1929 => x"8a",
          1930 => x"08",
          1931 => x"82",
          1932 => x"53",
          1933 => x"8a",
          1934 => x"82",
          1935 => x"f8",
          1936 => x"b5",
          1937 => x"05",
          1938 => x"b5",
          1939 => x"05",
          1940 => x"b5",
          1941 => x"05",
          1942 => x"a8",
          1943 => x"0d",
          1944 => x"0c",
          1945 => x"b4",
          1946 => x"b5",
          1947 => x"3d",
          1948 => x"82",
          1949 => x"f8",
          1950 => x"b5",
          1951 => x"05",
          1952 => x"33",
          1953 => x"70",
          1954 => x"81",
          1955 => x"51",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"b4",
          1959 => x"0c",
          1960 => x"82",
          1961 => x"88",
          1962 => x"72",
          1963 => x"b4",
          1964 => x"08",
          1965 => x"b5",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"72",
          1971 => x"38",
          1972 => x"08",
          1973 => x"82",
          1974 => x"8c",
          1975 => x"82",
          1976 => x"fc",
          1977 => x"90",
          1978 => x"53",
          1979 => x"b5",
          1980 => x"72",
          1981 => x"ab",
          1982 => x"82",
          1983 => x"f8",
          1984 => x"9f",
          1985 => x"b4",
          1986 => x"08",
          1987 => x"b4",
          1988 => x"0c",
          1989 => x"b4",
          1990 => x"08",
          1991 => x"0c",
          1992 => x"82",
          1993 => x"04",
          1994 => x"08",
          1995 => x"b4",
          1996 => x"0d",
          1997 => x"08",
          1998 => x"b4",
          1999 => x"08",
          2000 => x"82",
          2001 => x"70",
          2002 => x"0c",
          2003 => x"0d",
          2004 => x"0c",
          2005 => x"b4",
          2006 => x"b5",
          2007 => x"3d",
          2008 => x"b4",
          2009 => x"08",
          2010 => x"70",
          2011 => x"81",
          2012 => x"06",
          2013 => x"51",
          2014 => x"2e",
          2015 => x"0b",
          2016 => x"08",
          2017 => x"81",
          2018 => x"b5",
          2019 => x"05",
          2020 => x"33",
          2021 => x"70",
          2022 => x"51",
          2023 => x"80",
          2024 => x"38",
          2025 => x"08",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"54",
          2029 => x"88",
          2030 => x"9f",
          2031 => x"b4",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"57",
          2036 => x"75",
          2037 => x"81",
          2038 => x"82",
          2039 => x"8c",
          2040 => x"11",
          2041 => x"8c",
          2042 => x"b5",
          2043 => x"05",
          2044 => x"b5",
          2045 => x"05",
          2046 => x"80",
          2047 => x"b5",
          2048 => x"05",
          2049 => x"b4",
          2050 => x"08",
          2051 => x"b4",
          2052 => x"08",
          2053 => x"06",
          2054 => x"08",
          2055 => x"72",
          2056 => x"a8",
          2057 => x"a3",
          2058 => x"b4",
          2059 => x"08",
          2060 => x"81",
          2061 => x"0c",
          2062 => x"08",
          2063 => x"70",
          2064 => x"08",
          2065 => x"51",
          2066 => x"ff",
          2067 => x"b4",
          2068 => x"0c",
          2069 => x"08",
          2070 => x"82",
          2071 => x"87",
          2072 => x"b5",
          2073 => x"82",
          2074 => x"02",
          2075 => x"0c",
          2076 => x"82",
          2077 => x"88",
          2078 => x"11",
          2079 => x"32",
          2080 => x"51",
          2081 => x"71",
          2082 => x"38",
          2083 => x"b5",
          2084 => x"05",
          2085 => x"39",
          2086 => x"08",
          2087 => x"85",
          2088 => x"86",
          2089 => x"06",
          2090 => x"52",
          2091 => x"80",
          2092 => x"b5",
          2093 => x"05",
          2094 => x"b4",
          2095 => x"08",
          2096 => x"12",
          2097 => x"bf",
          2098 => x"71",
          2099 => x"82",
          2100 => x"88",
          2101 => x"11",
          2102 => x"8c",
          2103 => x"b5",
          2104 => x"05",
          2105 => x"33",
          2106 => x"b4",
          2107 => x"0c",
          2108 => x"82",
          2109 => x"b5",
          2110 => x"05",
          2111 => x"33",
          2112 => x"70",
          2113 => x"51",
          2114 => x"80",
          2115 => x"38",
          2116 => x"08",
          2117 => x"70",
          2118 => x"82",
          2119 => x"fc",
          2120 => x"52",
          2121 => x"08",
          2122 => x"a9",
          2123 => x"b4",
          2124 => x"08",
          2125 => x"08",
          2126 => x"53",
          2127 => x"33",
          2128 => x"51",
          2129 => x"14",
          2130 => x"82",
          2131 => x"f8",
          2132 => x"d7",
          2133 => x"b4",
          2134 => x"08",
          2135 => x"05",
          2136 => x"81",
          2137 => x"b5",
          2138 => x"05",
          2139 => x"b4",
          2140 => x"08",
          2141 => x"08",
          2142 => x"2d",
          2143 => x"08",
          2144 => x"b4",
          2145 => x"0c",
          2146 => x"b4",
          2147 => x"08",
          2148 => x"f2",
          2149 => x"b4",
          2150 => x"08",
          2151 => x"08",
          2152 => x"82",
          2153 => x"88",
          2154 => x"11",
          2155 => x"b4",
          2156 => x"0c",
          2157 => x"b4",
          2158 => x"08",
          2159 => x"81",
          2160 => x"82",
          2161 => x"f0",
          2162 => x"07",
          2163 => x"b5",
          2164 => x"05",
          2165 => x"82",
          2166 => x"f0",
          2167 => x"07",
          2168 => x"b5",
          2169 => x"05",
          2170 => x"b4",
          2171 => x"08",
          2172 => x"b4",
          2173 => x"33",
          2174 => x"ff",
          2175 => x"b4",
          2176 => x"0c",
          2177 => x"b5",
          2178 => x"05",
          2179 => x"08",
          2180 => x"12",
          2181 => x"b4",
          2182 => x"08",
          2183 => x"06",
          2184 => x"b4",
          2185 => x"0c",
          2186 => x"82",
          2187 => x"f8",
          2188 => x"b5",
          2189 => x"3d",
          2190 => x"b4",
          2191 => x"b5",
          2192 => x"82",
          2193 => x"fd",
          2194 => x"b5",
          2195 => x"05",
          2196 => x"b4",
          2197 => x"0c",
          2198 => x"08",
          2199 => x"82",
          2200 => x"f8",
          2201 => x"b5",
          2202 => x"05",
          2203 => x"82",
          2204 => x"b5",
          2205 => x"05",
          2206 => x"b4",
          2207 => x"08",
          2208 => x"38",
          2209 => x"08",
          2210 => x"82",
          2211 => x"90",
          2212 => x"51",
          2213 => x"08",
          2214 => x"71",
          2215 => x"38",
          2216 => x"08",
          2217 => x"82",
          2218 => x"90",
          2219 => x"82",
          2220 => x"fc",
          2221 => x"b5",
          2222 => x"05",
          2223 => x"b4",
          2224 => x"08",
          2225 => x"b4",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"81",
          2229 => x"b4",
          2230 => x"0c",
          2231 => x"08",
          2232 => x"ff",
          2233 => x"b4",
          2234 => x"0c",
          2235 => x"08",
          2236 => x"80",
          2237 => x"38",
          2238 => x"08",
          2239 => x"ff",
          2240 => x"b4",
          2241 => x"0c",
          2242 => x"08",
          2243 => x"ff",
          2244 => x"b4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"82",
          2248 => x"f8",
          2249 => x"51",
          2250 => x"34",
          2251 => x"82",
          2252 => x"90",
          2253 => x"05",
          2254 => x"08",
          2255 => x"82",
          2256 => x"90",
          2257 => x"05",
          2258 => x"08",
          2259 => x"82",
          2260 => x"90",
          2261 => x"2e",
          2262 => x"b5",
          2263 => x"05",
          2264 => x"33",
          2265 => x"08",
          2266 => x"81",
          2267 => x"b4",
          2268 => x"0c",
          2269 => x"08",
          2270 => x"52",
          2271 => x"34",
          2272 => x"08",
          2273 => x"81",
          2274 => x"b4",
          2275 => x"0c",
          2276 => x"82",
          2277 => x"88",
          2278 => x"82",
          2279 => x"51",
          2280 => x"82",
          2281 => x"04",
          2282 => x"08",
          2283 => x"b4",
          2284 => x"0d",
          2285 => x"08",
          2286 => x"82",
          2287 => x"fc",
          2288 => x"b5",
          2289 => x"05",
          2290 => x"33",
          2291 => x"08",
          2292 => x"81",
          2293 => x"b4",
          2294 => x"0c",
          2295 => x"06",
          2296 => x"80",
          2297 => x"da",
          2298 => x"b4",
          2299 => x"08",
          2300 => x"b5",
          2301 => x"05",
          2302 => x"b4",
          2303 => x"08",
          2304 => x"08",
          2305 => x"31",
          2306 => x"a8",
          2307 => x"3d",
          2308 => x"b4",
          2309 => x"b5",
          2310 => x"82",
          2311 => x"fe",
          2312 => x"b5",
          2313 => x"05",
          2314 => x"b4",
          2315 => x"0c",
          2316 => x"08",
          2317 => x"52",
          2318 => x"b5",
          2319 => x"05",
          2320 => x"82",
          2321 => x"8c",
          2322 => x"b5",
          2323 => x"05",
          2324 => x"70",
          2325 => x"b5",
          2326 => x"05",
          2327 => x"82",
          2328 => x"fc",
          2329 => x"81",
          2330 => x"70",
          2331 => x"38",
          2332 => x"82",
          2333 => x"88",
          2334 => x"82",
          2335 => x"51",
          2336 => x"82",
          2337 => x"04",
          2338 => x"08",
          2339 => x"b4",
          2340 => x"0d",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"b5",
          2345 => x"05",
          2346 => x"b4",
          2347 => x"0c",
          2348 => x"08",
          2349 => x"80",
          2350 => x"38",
          2351 => x"08",
          2352 => x"81",
          2353 => x"b4",
          2354 => x"0c",
          2355 => x"08",
          2356 => x"ff",
          2357 => x"b4",
          2358 => x"0c",
          2359 => x"08",
          2360 => x"80",
          2361 => x"82",
          2362 => x"f8",
          2363 => x"70",
          2364 => x"b4",
          2365 => x"08",
          2366 => x"b5",
          2367 => x"05",
          2368 => x"b4",
          2369 => x"08",
          2370 => x"71",
          2371 => x"b4",
          2372 => x"08",
          2373 => x"b5",
          2374 => x"05",
          2375 => x"39",
          2376 => x"08",
          2377 => x"70",
          2378 => x"0c",
          2379 => x"0d",
          2380 => x"0c",
          2381 => x"b4",
          2382 => x"b5",
          2383 => x"3d",
          2384 => x"b4",
          2385 => x"08",
          2386 => x"f4",
          2387 => x"b4",
          2388 => x"08",
          2389 => x"82",
          2390 => x"8c",
          2391 => x"05",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"33",
          2396 => x"06",
          2397 => x"51",
          2398 => x"84",
          2399 => x"39",
          2400 => x"08",
          2401 => x"52",
          2402 => x"b5",
          2403 => x"05",
          2404 => x"82",
          2405 => x"88",
          2406 => x"81",
          2407 => x"51",
          2408 => x"80",
          2409 => x"b4",
          2410 => x"0c",
          2411 => x"82",
          2412 => x"90",
          2413 => x"05",
          2414 => x"08",
          2415 => x"82",
          2416 => x"90",
          2417 => x"2e",
          2418 => x"81",
          2419 => x"b4",
          2420 => x"08",
          2421 => x"e8",
          2422 => x"b4",
          2423 => x"08",
          2424 => x"53",
          2425 => x"ff",
          2426 => x"b4",
          2427 => x"0c",
          2428 => x"82",
          2429 => x"8c",
          2430 => x"05",
          2431 => x"08",
          2432 => x"82",
          2433 => x"8c",
          2434 => x"33",
          2435 => x"8c",
          2436 => x"82",
          2437 => x"fc",
          2438 => x"39",
          2439 => x"08",
          2440 => x"70",
          2441 => x"b4",
          2442 => x"08",
          2443 => x"71",
          2444 => x"b5",
          2445 => x"05",
          2446 => x"52",
          2447 => x"39",
          2448 => x"b5",
          2449 => x"05",
          2450 => x"b4",
          2451 => x"08",
          2452 => x"0c",
          2453 => x"82",
          2454 => x"04",
          2455 => x"08",
          2456 => x"b4",
          2457 => x"0d",
          2458 => x"08",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"b5",
          2462 => x"05",
          2463 => x"80",
          2464 => x"b4",
          2465 => x"0c",
          2466 => x"82",
          2467 => x"f8",
          2468 => x"71",
          2469 => x"b4",
          2470 => x"08",
          2471 => x"b5",
          2472 => x"05",
          2473 => x"ff",
          2474 => x"70",
          2475 => x"38",
          2476 => x"08",
          2477 => x"ff",
          2478 => x"b4",
          2479 => x"0c",
          2480 => x"08",
          2481 => x"ff",
          2482 => x"ff",
          2483 => x"b5",
          2484 => x"05",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"b5",
          2488 => x"05",
          2489 => x"b4",
          2490 => x"08",
          2491 => x"b5",
          2492 => x"05",
          2493 => x"b5",
          2494 => x"05",
          2495 => x"a8",
          2496 => x"0d",
          2497 => x"0c",
          2498 => x"b4",
          2499 => x"b5",
          2500 => x"3d",
          2501 => x"b4",
          2502 => x"08",
          2503 => x"08",
          2504 => x"82",
          2505 => x"90",
          2506 => x"2e",
          2507 => x"82",
          2508 => x"90",
          2509 => x"05",
          2510 => x"08",
          2511 => x"82",
          2512 => x"90",
          2513 => x"05",
          2514 => x"08",
          2515 => x"82",
          2516 => x"90",
          2517 => x"2e",
          2518 => x"b5",
          2519 => x"05",
          2520 => x"82",
          2521 => x"fc",
          2522 => x"52",
          2523 => x"82",
          2524 => x"fc",
          2525 => x"05",
          2526 => x"08",
          2527 => x"ff",
          2528 => x"b5",
          2529 => x"05",
          2530 => x"b5",
          2531 => x"84",
          2532 => x"b5",
          2533 => x"82",
          2534 => x"02",
          2535 => x"0c",
          2536 => x"80",
          2537 => x"b4",
          2538 => x"0c",
          2539 => x"08",
          2540 => x"80",
          2541 => x"82",
          2542 => x"88",
          2543 => x"82",
          2544 => x"88",
          2545 => x"0b",
          2546 => x"08",
          2547 => x"82",
          2548 => x"fc",
          2549 => x"38",
          2550 => x"b5",
          2551 => x"05",
          2552 => x"b4",
          2553 => x"08",
          2554 => x"08",
          2555 => x"82",
          2556 => x"8c",
          2557 => x"25",
          2558 => x"b5",
          2559 => x"05",
          2560 => x"b5",
          2561 => x"05",
          2562 => x"82",
          2563 => x"f0",
          2564 => x"b5",
          2565 => x"05",
          2566 => x"81",
          2567 => x"b4",
          2568 => x"0c",
          2569 => x"08",
          2570 => x"82",
          2571 => x"fc",
          2572 => x"53",
          2573 => x"08",
          2574 => x"52",
          2575 => x"08",
          2576 => x"51",
          2577 => x"82",
          2578 => x"70",
          2579 => x"08",
          2580 => x"54",
          2581 => x"08",
          2582 => x"80",
          2583 => x"82",
          2584 => x"f8",
          2585 => x"82",
          2586 => x"f8",
          2587 => x"b5",
          2588 => x"05",
          2589 => x"b5",
          2590 => x"89",
          2591 => x"b5",
          2592 => x"82",
          2593 => x"02",
          2594 => x"0c",
          2595 => x"80",
          2596 => x"b4",
          2597 => x"0c",
          2598 => x"08",
          2599 => x"80",
          2600 => x"82",
          2601 => x"88",
          2602 => x"82",
          2603 => x"88",
          2604 => x"0b",
          2605 => x"08",
          2606 => x"82",
          2607 => x"8c",
          2608 => x"25",
          2609 => x"b5",
          2610 => x"05",
          2611 => x"b5",
          2612 => x"05",
          2613 => x"82",
          2614 => x"8c",
          2615 => x"82",
          2616 => x"88",
          2617 => x"81",
          2618 => x"b5",
          2619 => x"82",
          2620 => x"f8",
          2621 => x"82",
          2622 => x"fc",
          2623 => x"2e",
          2624 => x"b5",
          2625 => x"05",
          2626 => x"b5",
          2627 => x"05",
          2628 => x"b4",
          2629 => x"08",
          2630 => x"a8",
          2631 => x"3d",
          2632 => x"b4",
          2633 => x"b5",
          2634 => x"82",
          2635 => x"fd",
          2636 => x"53",
          2637 => x"08",
          2638 => x"52",
          2639 => x"08",
          2640 => x"51",
          2641 => x"82",
          2642 => x"70",
          2643 => x"0c",
          2644 => x"0d",
          2645 => x"0c",
          2646 => x"b4",
          2647 => x"b5",
          2648 => x"3d",
          2649 => x"82",
          2650 => x"8c",
          2651 => x"82",
          2652 => x"88",
          2653 => x"93",
          2654 => x"a8",
          2655 => x"b5",
          2656 => x"85",
          2657 => x"b5",
          2658 => x"82",
          2659 => x"02",
          2660 => x"0c",
          2661 => x"81",
          2662 => x"b4",
          2663 => x"0c",
          2664 => x"b5",
          2665 => x"05",
          2666 => x"b4",
          2667 => x"08",
          2668 => x"08",
          2669 => x"27",
          2670 => x"b5",
          2671 => x"05",
          2672 => x"ae",
          2673 => x"82",
          2674 => x"8c",
          2675 => x"a2",
          2676 => x"b4",
          2677 => x"08",
          2678 => x"b4",
          2679 => x"0c",
          2680 => x"08",
          2681 => x"10",
          2682 => x"08",
          2683 => x"ff",
          2684 => x"b5",
          2685 => x"05",
          2686 => x"80",
          2687 => x"b5",
          2688 => x"05",
          2689 => x"b4",
          2690 => x"08",
          2691 => x"82",
          2692 => x"88",
          2693 => x"b5",
          2694 => x"05",
          2695 => x"b5",
          2696 => x"05",
          2697 => x"b4",
          2698 => x"08",
          2699 => x"08",
          2700 => x"07",
          2701 => x"08",
          2702 => x"82",
          2703 => x"fc",
          2704 => x"2a",
          2705 => x"08",
          2706 => x"82",
          2707 => x"8c",
          2708 => x"2a",
          2709 => x"08",
          2710 => x"ff",
          2711 => x"b5",
          2712 => x"05",
          2713 => x"93",
          2714 => x"b4",
          2715 => x"08",
          2716 => x"b4",
          2717 => x"0c",
          2718 => x"82",
          2719 => x"f8",
          2720 => x"82",
          2721 => x"f4",
          2722 => x"82",
          2723 => x"f4",
          2724 => x"b5",
          2725 => x"3d",
          2726 => x"b4",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"f1",
          2733 => x"b5",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"a8",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"c5",
          2748 => x"a8",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"a8",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"9a",
          2766 => x"f9",
          2767 => x"ac",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"9a",
          2773 => x"dd",
          2774 => x"f4",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"9b",
          2780 => x"c1",
          2781 => x"cc",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"fc",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"bc",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"f0",
          2791 => x"82",
          2792 => x"91",
          2793 => x"a0",
          2794 => x"82",
          2795 => x"85",
          2796 => x"c4",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"fa",
          2806 => x"b5",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"d4",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"dc",
          2830 => x"a8",
          2831 => x"b5",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"a8",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"83",
          2840 => x"b5",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"81",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"b5",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"58",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"a8",
          2868 => x"76",
          2869 => x"38",
          2870 => x"9a",
          2871 => x"62",
          2872 => x"60",
          2873 => x"a8",
          2874 => x"7e",
          2875 => x"82",
          2876 => x"58",
          2877 => x"04",
          2878 => x"a8",
          2879 => x"0d",
          2880 => x"0d",
          2881 => x"02",
          2882 => x"cf",
          2883 => x"73",
          2884 => x"5f",
          2885 => x"5e",
          2886 => x"82",
          2887 => x"ff",
          2888 => x"82",
          2889 => x"e0",
          2890 => x"55",
          2891 => x"80",
          2892 => x"90",
          2893 => x"7b",
          2894 => x"38",
          2895 => x"74",
          2896 => x"7a",
          2897 => x"72",
          2898 => x"9e",
          2899 => x"b9",
          2900 => x"39",
          2901 => x"51",
          2902 => x"82",
          2903 => x"c1",
          2904 => x"53",
          2905 => x"8e",
          2906 => x"52",
          2907 => x"51",
          2908 => x"3f",
          2909 => x"9e",
          2910 => x"8a",
          2911 => x"55",
          2912 => x"18",
          2913 => x"27",
          2914 => x"33",
          2915 => x"a0",
          2916 => x"c5",
          2917 => x"82",
          2918 => x"df",
          2919 => x"15",
          2920 => x"fc",
          2921 => x"51",
          2922 => x"fe",
          2923 => x"9e",
          2924 => x"d2",
          2925 => x"74",
          2926 => x"c6",
          2927 => x"70",
          2928 => x"80",
          2929 => x"27",
          2930 => x"56",
          2931 => x"74",
          2932 => x"81",
          2933 => x"06",
          2934 => x"06",
          2935 => x"80",
          2936 => x"73",
          2937 => x"8a",
          2938 => x"fc",
          2939 => x"51",
          2940 => x"cc",
          2941 => x"a0",
          2942 => x"3f",
          2943 => x"ff",
          2944 => x"9e",
          2945 => x"fe",
          2946 => x"79",
          2947 => x"9c",
          2948 => x"b5",
          2949 => x"2b",
          2950 => x"51",
          2951 => x"2e",
          2952 => x"aa",
          2953 => x"3f",
          2954 => x"08",
          2955 => x"98",
          2956 => x"32",
          2957 => x"9b",
          2958 => x"70",
          2959 => x"75",
          2960 => x"58",
          2961 => x"51",
          2962 => x"24",
          2963 => x"9b",
          2964 => x"06",
          2965 => x"53",
          2966 => x"1e",
          2967 => x"26",
          2968 => x"ff",
          2969 => x"b5",
          2970 => x"3d",
          2971 => x"3d",
          2972 => x"05",
          2973 => x"b4",
          2974 => x"b8",
          2975 => x"b6",
          2976 => x"b4",
          2977 => x"a5",
          2978 => x"9e",
          2979 => x"9e",
          2980 => x"b4",
          2981 => x"82",
          2982 => x"ff",
          2983 => x"74",
          2984 => x"38",
          2985 => x"86",
          2986 => x"fe",
          2987 => x"c0",
          2988 => x"53",
          2989 => x"81",
          2990 => x"3f",
          2991 => x"51",
          2992 => x"80",
          2993 => x"3f",
          2994 => x"70",
          2995 => x"52",
          2996 => x"92",
          2997 => x"97",
          2998 => x"9f",
          2999 => x"fa",
          3000 => x"97",
          3001 => x"82",
          3002 => x"06",
          3003 => x"80",
          3004 => x"81",
          3005 => x"3f",
          3006 => x"51",
          3007 => x"80",
          3008 => x"3f",
          3009 => x"70",
          3010 => x"52",
          3011 => x"92",
          3012 => x"97",
          3013 => x"9f",
          3014 => x"be",
          3015 => x"97",
          3016 => x"84",
          3017 => x"06",
          3018 => x"80",
          3019 => x"81",
          3020 => x"3f",
          3021 => x"51",
          3022 => x"80",
          3023 => x"3f",
          3024 => x"70",
          3025 => x"52",
          3026 => x"92",
          3027 => x"96",
          3028 => x"9f",
          3029 => x"82",
          3030 => x"96",
          3031 => x"86",
          3032 => x"06",
          3033 => x"80",
          3034 => x"81",
          3035 => x"3f",
          3036 => x"51",
          3037 => x"80",
          3038 => x"3f",
          3039 => x"70",
          3040 => x"52",
          3041 => x"92",
          3042 => x"96",
          3043 => x"a0",
          3044 => x"c6",
          3045 => x"96",
          3046 => x"88",
          3047 => x"06",
          3048 => x"80",
          3049 => x"81",
          3050 => x"3f",
          3051 => x"51",
          3052 => x"80",
          3053 => x"3f",
          3054 => x"84",
          3055 => x"fb",
          3056 => x"02",
          3057 => x"05",
          3058 => x"56",
          3059 => x"75",
          3060 => x"3f",
          3061 => x"b0",
          3062 => x"73",
          3063 => x"53",
          3064 => x"52",
          3065 => x"51",
          3066 => x"3f",
          3067 => x"08",
          3068 => x"b5",
          3069 => x"80",
          3070 => x"31",
          3071 => x"73",
          3072 => x"b0",
          3073 => x"0b",
          3074 => x"33",
          3075 => x"2e",
          3076 => x"af",
          3077 => x"a8",
          3078 => x"75",
          3079 => x"da",
          3080 => x"a8",
          3081 => x"8b",
          3082 => x"a8",
          3083 => x"d6",
          3084 => x"82",
          3085 => x"81",
          3086 => x"82",
          3087 => x"82",
          3088 => x"0b",
          3089 => x"a4",
          3090 => x"82",
          3091 => x"06",
          3092 => x"a0",
          3093 => x"52",
          3094 => x"a2",
          3095 => x"82",
          3096 => x"87",
          3097 => x"cd",
          3098 => x"70",
          3099 => x"a4",
          3100 => x"81",
          3101 => x"80",
          3102 => x"82",
          3103 => x"81",
          3104 => x"79",
          3105 => x"81",
          3106 => x"97",
          3107 => x"53",
          3108 => x"52",
          3109 => x"f0",
          3110 => x"79",
          3111 => x"d4",
          3112 => x"8f",
          3113 => x"a8",
          3114 => x"88",
          3115 => x"f0",
          3116 => x"39",
          3117 => x"5e",
          3118 => x"51",
          3119 => x"97",
          3120 => x"5b",
          3121 => x"7a",
          3122 => x"3f",
          3123 => x"84",
          3124 => x"ca",
          3125 => x"a8",
          3126 => x"70",
          3127 => x"5a",
          3128 => x"2e",
          3129 => x"79",
          3130 => x"b2",
          3131 => x"2e",
          3132 => x"79",
          3133 => x"38",
          3134 => x"ff",
          3135 => x"bc",
          3136 => x"38",
          3137 => x"79",
          3138 => x"83",
          3139 => x"80",
          3140 => x"c9",
          3141 => x"2e",
          3142 => x"8a",
          3143 => x"80",
          3144 => x"c5",
          3145 => x"f9",
          3146 => x"79",
          3147 => x"87",
          3148 => x"80",
          3149 => x"8d",
          3150 => x"39",
          3151 => x"2e",
          3152 => x"79",
          3153 => x"8b",
          3154 => x"82",
          3155 => x"38",
          3156 => x"79",
          3157 => x"89",
          3158 => x"ea",
          3159 => x"ff",
          3160 => x"ff",
          3161 => x"d2",
          3162 => x"b5",
          3163 => x"2e",
          3164 => x"b5",
          3165 => x"11",
          3166 => x"05",
          3167 => x"3f",
          3168 => x"08",
          3169 => x"b0",
          3170 => x"fe",
          3171 => x"ff",
          3172 => x"d2",
          3173 => x"b5",
          3174 => x"38",
          3175 => x"08",
          3176 => x"ac",
          3177 => x"3f",
          3178 => x"5b",
          3179 => x"81",
          3180 => x"5a",
          3181 => x"84",
          3182 => x"7b",
          3183 => x"38",
          3184 => x"b5",
          3185 => x"11",
          3186 => x"05",
          3187 => x"3f",
          3188 => x"08",
          3189 => x"e0",
          3190 => x"fe",
          3191 => x"ff",
          3192 => x"d1",
          3193 => x"b5",
          3194 => x"2e",
          3195 => x"b5",
          3196 => x"11",
          3197 => x"05",
          3198 => x"3f",
          3199 => x"08",
          3200 => x"b4",
          3201 => x"bc",
          3202 => x"3f",
          3203 => x"64",
          3204 => x"38",
          3205 => x"70",
          3206 => x"33",
          3207 => x"81",
          3208 => x"39",
          3209 => x"80",
          3210 => x"84",
          3211 => x"85",
          3212 => x"a8",
          3213 => x"fc",
          3214 => x"3d",
          3215 => x"53",
          3216 => x"51",
          3217 => x"82",
          3218 => x"80",
          3219 => x"38",
          3220 => x"f8",
          3221 => x"84",
          3222 => x"d9",
          3223 => x"a8",
          3224 => x"fc",
          3225 => x"a1",
          3226 => x"9a",
          3227 => x"7a",
          3228 => x"38",
          3229 => x"7c",
          3230 => x"5c",
          3231 => x"92",
          3232 => x"7b",
          3233 => x"53",
          3234 => x"a1",
          3235 => x"ae",
          3236 => x"1b",
          3237 => x"44",
          3238 => x"82",
          3239 => x"89",
          3240 => x"3d",
          3241 => x"53",
          3242 => x"51",
          3243 => x"82",
          3244 => x"80",
          3245 => x"b4",
          3246 => x"79",
          3247 => x"38",
          3248 => x"08",
          3249 => x"39",
          3250 => x"33",
          3251 => x"2e",
          3252 => x"b3",
          3253 => x"bc",
          3254 => x"96",
          3255 => x"80",
          3256 => x"82",
          3257 => x"45",
          3258 => x"b4",
          3259 => x"79",
          3260 => x"38",
          3261 => x"08",
          3262 => x"82",
          3263 => x"5a",
          3264 => x"88",
          3265 => x"ec",
          3266 => x"39",
          3267 => x"08",
          3268 => x"45",
          3269 => x"fc",
          3270 => x"84",
          3271 => x"95",
          3272 => x"a8",
          3273 => x"38",
          3274 => x"33",
          3275 => x"2e",
          3276 => x"b3",
          3277 => x"80",
          3278 => x"b4",
          3279 => x"79",
          3280 => x"38",
          3281 => x"08",
          3282 => x"82",
          3283 => x"5a",
          3284 => x"88",
          3285 => x"e0",
          3286 => x"39",
          3287 => x"33",
          3288 => x"2e",
          3289 => x"b3",
          3290 => x"99",
          3291 => x"92",
          3292 => x"80",
          3293 => x"82",
          3294 => x"44",
          3295 => x"b3",
          3296 => x"05",
          3297 => x"fe",
          3298 => x"ff",
          3299 => x"ce",
          3300 => x"b5",
          3301 => x"2e",
          3302 => x"63",
          3303 => x"88",
          3304 => x"81",
          3305 => x"32",
          3306 => x"72",
          3307 => x"70",
          3308 => x"51",
          3309 => x"80",
          3310 => x"7b",
          3311 => x"38",
          3312 => x"a1",
          3313 => x"be",
          3314 => x"64",
          3315 => x"63",
          3316 => x"f2",
          3317 => x"a2",
          3318 => x"ec",
          3319 => x"ff",
          3320 => x"ff",
          3321 => x"cd",
          3322 => x"b5",
          3323 => x"2e",
          3324 => x"b5",
          3325 => x"11",
          3326 => x"05",
          3327 => x"3f",
          3328 => x"08",
          3329 => x"38",
          3330 => x"80",
          3331 => x"7a",
          3332 => x"05",
          3333 => x"fe",
          3334 => x"ff",
          3335 => x"cd",
          3336 => x"b5",
          3337 => x"38",
          3338 => x"64",
          3339 => x"52",
          3340 => x"51",
          3341 => x"3f",
          3342 => x"7a",
          3343 => x"3f",
          3344 => x"33",
          3345 => x"2e",
          3346 => x"9f",
          3347 => x"38",
          3348 => x"fc",
          3349 => x"84",
          3350 => x"d9",
          3351 => x"a8",
          3352 => x"91",
          3353 => x"02",
          3354 => x"33",
          3355 => x"81",
          3356 => x"b7",
          3357 => x"9c",
          3358 => x"3f",
          3359 => x"b5",
          3360 => x"11",
          3361 => x"05",
          3362 => x"3f",
          3363 => x"08",
          3364 => x"a4",
          3365 => x"fe",
          3366 => x"ff",
          3367 => x"c6",
          3368 => x"b5",
          3369 => x"2e",
          3370 => x"5a",
          3371 => x"05",
          3372 => x"82",
          3373 => x"79",
          3374 => x"fe",
          3375 => x"ff",
          3376 => x"c5",
          3377 => x"b5",
          3378 => x"38",
          3379 => x"61",
          3380 => x"52",
          3381 => x"51",
          3382 => x"3f",
          3383 => x"7a",
          3384 => x"3f",
          3385 => x"33",
          3386 => x"2e",
          3387 => x"79",
          3388 => x"38",
          3389 => x"42",
          3390 => x"3d",
          3391 => x"53",
          3392 => x"51",
          3393 => x"82",
          3394 => x"80",
          3395 => x"61",
          3396 => x"c2",
          3397 => x"70",
          3398 => x"23",
          3399 => x"af",
          3400 => x"9c",
          3401 => x"3f",
          3402 => x"b5",
          3403 => x"11",
          3404 => x"05",
          3405 => x"3f",
          3406 => x"08",
          3407 => x"f8",
          3408 => x"fe",
          3409 => x"ff",
          3410 => x"c4",
          3411 => x"b5",
          3412 => x"2e",
          3413 => x"61",
          3414 => x"61",
          3415 => x"b5",
          3416 => x"11",
          3417 => x"05",
          3418 => x"3f",
          3419 => x"08",
          3420 => x"c4",
          3421 => x"08",
          3422 => x"a2",
          3423 => x"a8",
          3424 => x"f8",
          3425 => x"c9",
          3426 => x"46",
          3427 => x"79",
          3428 => x"a4",
          3429 => x"27",
          3430 => x"3d",
          3431 => x"53",
          3432 => x"51",
          3433 => x"82",
          3434 => x"80",
          3435 => x"61",
          3436 => x"5a",
          3437 => x"42",
          3438 => x"82",
          3439 => x"cf",
          3440 => x"b1",
          3441 => x"ff",
          3442 => x"ff",
          3443 => x"c9",
          3444 => x"b5",
          3445 => x"2e",
          3446 => x"64",
          3447 => x"bc",
          3448 => x"f5",
          3449 => x"79",
          3450 => x"ff",
          3451 => x"ff",
          3452 => x"c9",
          3453 => x"b5",
          3454 => x"2e",
          3455 => x"64",
          3456 => x"d8",
          3457 => x"d1",
          3458 => x"79",
          3459 => x"a8",
          3460 => x"f5",
          3461 => x"b5",
          3462 => x"82",
          3463 => x"ff",
          3464 => x"f5",
          3465 => x"a3",
          3466 => x"da",
          3467 => x"8a",
          3468 => x"39",
          3469 => x"51",
          3470 => x"80",
          3471 => x"39",
          3472 => x"f4",
          3473 => x"46",
          3474 => x"79",
          3475 => x"e8",
          3476 => x"06",
          3477 => x"2e",
          3478 => x"b5",
          3479 => x"05",
          3480 => x"3f",
          3481 => x"08",
          3482 => x"7b",
          3483 => x"38",
          3484 => x"89",
          3485 => x"2e",
          3486 => x"cd",
          3487 => x"2e",
          3488 => x"c5",
          3489 => x"c0",
          3490 => x"82",
          3491 => x"80",
          3492 => x"c8",
          3493 => x"ff",
          3494 => x"ff",
          3495 => x"bb",
          3496 => x"e8",
          3497 => x"ff",
          3498 => x"ff",
          3499 => x"ab",
          3500 => x"82",
          3501 => x"80",
          3502 => x"d8",
          3503 => x"ff",
          3504 => x"ff",
          3505 => x"93",
          3506 => x"80",
          3507 => x"e4",
          3508 => x"ff",
          3509 => x"ff",
          3510 => x"82",
          3511 => x"82",
          3512 => x"82",
          3513 => x"80",
          3514 => x"80",
          3515 => x"80",
          3516 => x"80",
          3517 => x"ff",
          3518 => x"eb",
          3519 => x"b5",
          3520 => x"b5",
          3521 => x"70",
          3522 => x"07",
          3523 => x"5c",
          3524 => x"5b",
          3525 => x"83",
          3526 => x"79",
          3527 => x"79",
          3528 => x"38",
          3529 => x"81",
          3530 => x"5a",
          3531 => x"38",
          3532 => x"7e",
          3533 => x"5a",
          3534 => x"7f",
          3535 => x"81",
          3536 => x"38",
          3537 => x"51",
          3538 => x"f2",
          3539 => x"3d",
          3540 => x"82",
          3541 => x"87",
          3542 => x"70",
          3543 => x"87",
          3544 => x"72",
          3545 => x"3f",
          3546 => x"08",
          3547 => x"08",
          3548 => x"84",
          3549 => x"51",
          3550 => x"72",
          3551 => x"08",
          3552 => x"87",
          3553 => x"70",
          3554 => x"87",
          3555 => x"72",
          3556 => x"3f",
          3557 => x"08",
          3558 => x"08",
          3559 => x"84",
          3560 => x"51",
          3561 => x"72",
          3562 => x"08",
          3563 => x"8c",
          3564 => x"87",
          3565 => x"0c",
          3566 => x"0b",
          3567 => x"94",
          3568 => x"fc",
          3569 => x"3f",
          3570 => x"5a",
          3571 => x"5b",
          3572 => x"05",
          3573 => x"80",
          3574 => x"e4",
          3575 => x"fc",
          3576 => x"3f",
          3577 => x"82",
          3578 => x"cb",
          3579 => x"a4",
          3580 => x"92",
          3581 => x"b0",
          3582 => x"3f",
          3583 => x"51",
          3584 => x"81",
          3585 => x"3f",
          3586 => x"80",
          3587 => x"0d",
          3588 => x"53",
          3589 => x"52",
          3590 => x"82",
          3591 => x"81",
          3592 => x"07",
          3593 => x"52",
          3594 => x"e8",
          3595 => x"b5",
          3596 => x"3d",
          3597 => x"3d",
          3598 => x"08",
          3599 => x"73",
          3600 => x"74",
          3601 => x"38",
          3602 => x"70",
          3603 => x"81",
          3604 => x"81",
          3605 => x"39",
          3606 => x"70",
          3607 => x"81",
          3608 => x"81",
          3609 => x"54",
          3610 => x"81",
          3611 => x"06",
          3612 => x"39",
          3613 => x"80",
          3614 => x"54",
          3615 => x"83",
          3616 => x"70",
          3617 => x"38",
          3618 => x"98",
          3619 => x"52",
          3620 => x"52",
          3621 => x"2e",
          3622 => x"54",
          3623 => x"84",
          3624 => x"38",
          3625 => x"52",
          3626 => x"2e",
          3627 => x"83",
          3628 => x"70",
          3629 => x"30",
          3630 => x"76",
          3631 => x"51",
          3632 => x"88",
          3633 => x"70",
          3634 => x"34",
          3635 => x"72",
          3636 => x"b5",
          3637 => x"3d",
          3638 => x"3d",
          3639 => x"72",
          3640 => x"92",
          3641 => x"fc",
          3642 => x"51",
          3643 => x"3f",
          3644 => x"08",
          3645 => x"53",
          3646 => x"53",
          3647 => x"a8",
          3648 => x"0d",
          3649 => x"0d",
          3650 => x"33",
          3651 => x"53",
          3652 => x"8b",
          3653 => x"38",
          3654 => x"ff",
          3655 => x"52",
          3656 => x"81",
          3657 => x"13",
          3658 => x"52",
          3659 => x"80",
          3660 => x"13",
          3661 => x"52",
          3662 => x"80",
          3663 => x"13",
          3664 => x"52",
          3665 => x"80",
          3666 => x"13",
          3667 => x"52",
          3668 => x"26",
          3669 => x"8a",
          3670 => x"87",
          3671 => x"e7",
          3672 => x"38",
          3673 => x"c0",
          3674 => x"72",
          3675 => x"98",
          3676 => x"13",
          3677 => x"98",
          3678 => x"13",
          3679 => x"98",
          3680 => x"13",
          3681 => x"98",
          3682 => x"13",
          3683 => x"98",
          3684 => x"13",
          3685 => x"98",
          3686 => x"87",
          3687 => x"0c",
          3688 => x"98",
          3689 => x"0b",
          3690 => x"9c",
          3691 => x"71",
          3692 => x"0c",
          3693 => x"04",
          3694 => x"7f",
          3695 => x"98",
          3696 => x"7d",
          3697 => x"98",
          3698 => x"7d",
          3699 => x"c0",
          3700 => x"5a",
          3701 => x"34",
          3702 => x"b4",
          3703 => x"83",
          3704 => x"c0",
          3705 => x"5a",
          3706 => x"34",
          3707 => x"ac",
          3708 => x"85",
          3709 => x"c0",
          3710 => x"5a",
          3711 => x"34",
          3712 => x"a4",
          3713 => x"88",
          3714 => x"c0",
          3715 => x"5a",
          3716 => x"23",
          3717 => x"79",
          3718 => x"06",
          3719 => x"ff",
          3720 => x"86",
          3721 => x"85",
          3722 => x"84",
          3723 => x"83",
          3724 => x"82",
          3725 => x"7d",
          3726 => x"06",
          3727 => x"c8",
          3728 => x"95",
          3729 => x"0d",
          3730 => x"0d",
          3731 => x"33",
          3732 => x"33",
          3733 => x"06",
          3734 => x"87",
          3735 => x"51",
          3736 => x"86",
          3737 => x"94",
          3738 => x"08",
          3739 => x"70",
          3740 => x"54",
          3741 => x"2e",
          3742 => x"91",
          3743 => x"06",
          3744 => x"d7",
          3745 => x"32",
          3746 => x"51",
          3747 => x"2e",
          3748 => x"93",
          3749 => x"06",
          3750 => x"ff",
          3751 => x"81",
          3752 => x"87",
          3753 => x"52",
          3754 => x"86",
          3755 => x"94",
          3756 => x"72",
          3757 => x"b5",
          3758 => x"3d",
          3759 => x"3d",
          3760 => x"05",
          3761 => x"70",
          3762 => x"52",
          3763 => x"b3",
          3764 => x"3d",
          3765 => x"3d",
          3766 => x"05",
          3767 => x"8a",
          3768 => x"06",
          3769 => x"52",
          3770 => x"3f",
          3771 => x"33",
          3772 => x"06",
          3773 => x"c0",
          3774 => x"76",
          3775 => x"38",
          3776 => x"94",
          3777 => x"70",
          3778 => x"81",
          3779 => x"54",
          3780 => x"8c",
          3781 => x"2a",
          3782 => x"51",
          3783 => x"38",
          3784 => x"70",
          3785 => x"53",
          3786 => x"8d",
          3787 => x"2a",
          3788 => x"51",
          3789 => x"be",
          3790 => x"ff",
          3791 => x"c0",
          3792 => x"72",
          3793 => x"38",
          3794 => x"90",
          3795 => x"0c",
          3796 => x"b5",
          3797 => x"3d",
          3798 => x"3d",
          3799 => x"80",
          3800 => x"81",
          3801 => x"53",
          3802 => x"2e",
          3803 => x"71",
          3804 => x"81",
          3805 => x"c8",
          3806 => x"ff",
          3807 => x"55",
          3808 => x"94",
          3809 => x"80",
          3810 => x"87",
          3811 => x"51",
          3812 => x"96",
          3813 => x"06",
          3814 => x"70",
          3815 => x"38",
          3816 => x"70",
          3817 => x"51",
          3818 => x"72",
          3819 => x"81",
          3820 => x"70",
          3821 => x"38",
          3822 => x"70",
          3823 => x"51",
          3824 => x"38",
          3825 => x"06",
          3826 => x"94",
          3827 => x"80",
          3828 => x"87",
          3829 => x"52",
          3830 => x"81",
          3831 => x"70",
          3832 => x"53",
          3833 => x"ff",
          3834 => x"82",
          3835 => x"89",
          3836 => x"fe",
          3837 => x"b3",
          3838 => x"81",
          3839 => x"52",
          3840 => x"84",
          3841 => x"2e",
          3842 => x"c0",
          3843 => x"70",
          3844 => x"2a",
          3845 => x"51",
          3846 => x"80",
          3847 => x"71",
          3848 => x"51",
          3849 => x"80",
          3850 => x"2e",
          3851 => x"c0",
          3852 => x"71",
          3853 => x"ff",
          3854 => x"a8",
          3855 => x"3d",
          3856 => x"af",
          3857 => x"a8",
          3858 => x"06",
          3859 => x"0c",
          3860 => x"0d",
          3861 => x"33",
          3862 => x"06",
          3863 => x"c0",
          3864 => x"70",
          3865 => x"38",
          3866 => x"94",
          3867 => x"70",
          3868 => x"81",
          3869 => x"51",
          3870 => x"80",
          3871 => x"72",
          3872 => x"51",
          3873 => x"80",
          3874 => x"2e",
          3875 => x"c0",
          3876 => x"71",
          3877 => x"2b",
          3878 => x"51",
          3879 => x"82",
          3880 => x"84",
          3881 => x"ff",
          3882 => x"c0",
          3883 => x"70",
          3884 => x"06",
          3885 => x"80",
          3886 => x"38",
          3887 => x"a4",
          3888 => x"cc",
          3889 => x"9e",
          3890 => x"b3",
          3891 => x"c0",
          3892 => x"82",
          3893 => x"87",
          3894 => x"08",
          3895 => x"0c",
          3896 => x"9c",
          3897 => x"dc",
          3898 => x"9e",
          3899 => x"b3",
          3900 => x"c0",
          3901 => x"82",
          3902 => x"87",
          3903 => x"08",
          3904 => x"0c",
          3905 => x"b4",
          3906 => x"ec",
          3907 => x"9e",
          3908 => x"b3",
          3909 => x"c0",
          3910 => x"82",
          3911 => x"87",
          3912 => x"08",
          3913 => x"0c",
          3914 => x"c4",
          3915 => x"fc",
          3916 => x"9e",
          3917 => x"70",
          3918 => x"23",
          3919 => x"84",
          3920 => x"84",
          3921 => x"9e",
          3922 => x"b4",
          3923 => x"c0",
          3924 => x"82",
          3925 => x"81",
          3926 => x"90",
          3927 => x"87",
          3928 => x"08",
          3929 => x"0a",
          3930 => x"52",
          3931 => x"83",
          3932 => x"71",
          3933 => x"34",
          3934 => x"c0",
          3935 => x"70",
          3936 => x"06",
          3937 => x"70",
          3938 => x"38",
          3939 => x"82",
          3940 => x"80",
          3941 => x"9e",
          3942 => x"90",
          3943 => x"51",
          3944 => x"80",
          3945 => x"81",
          3946 => x"b4",
          3947 => x"0b",
          3948 => x"90",
          3949 => x"80",
          3950 => x"52",
          3951 => x"2e",
          3952 => x"52",
          3953 => x"94",
          3954 => x"87",
          3955 => x"08",
          3956 => x"80",
          3957 => x"52",
          3958 => x"83",
          3959 => x"71",
          3960 => x"34",
          3961 => x"c0",
          3962 => x"70",
          3963 => x"06",
          3964 => x"70",
          3965 => x"38",
          3966 => x"82",
          3967 => x"80",
          3968 => x"9e",
          3969 => x"84",
          3970 => x"51",
          3971 => x"80",
          3972 => x"81",
          3973 => x"b4",
          3974 => x"0b",
          3975 => x"90",
          3976 => x"80",
          3977 => x"52",
          3978 => x"2e",
          3979 => x"52",
          3980 => x"98",
          3981 => x"87",
          3982 => x"08",
          3983 => x"80",
          3984 => x"52",
          3985 => x"83",
          3986 => x"71",
          3987 => x"34",
          3988 => x"c0",
          3989 => x"70",
          3990 => x"06",
          3991 => x"70",
          3992 => x"38",
          3993 => x"82",
          3994 => x"80",
          3995 => x"9e",
          3996 => x"a0",
          3997 => x"52",
          3998 => x"2e",
          3999 => x"52",
          4000 => x"9b",
          4001 => x"9e",
          4002 => x"98",
          4003 => x"8a",
          4004 => x"51",
          4005 => x"9c",
          4006 => x"87",
          4007 => x"08",
          4008 => x"06",
          4009 => x"70",
          4010 => x"38",
          4011 => x"82",
          4012 => x"87",
          4013 => x"08",
          4014 => x"06",
          4015 => x"51",
          4016 => x"82",
          4017 => x"80",
          4018 => x"9e",
          4019 => x"88",
          4020 => x"52",
          4021 => x"83",
          4022 => x"71",
          4023 => x"34",
          4024 => x"90",
          4025 => x"06",
          4026 => x"82",
          4027 => x"83",
          4028 => x"fb",
          4029 => x"a4",
          4030 => x"bd",
          4031 => x"b4",
          4032 => x"73",
          4033 => x"38",
          4034 => x"51",
          4035 => x"3f",
          4036 => x"51",
          4037 => x"3f",
          4038 => x"33",
          4039 => x"2e",
          4040 => x"b3",
          4041 => x"b3",
          4042 => x"54",
          4043 => x"a0",
          4044 => x"a5",
          4045 => x"97",
          4046 => x"80",
          4047 => x"82",
          4048 => x"82",
          4049 => x"11",
          4050 => x"a5",
          4051 => x"95",
          4052 => x"b4",
          4053 => x"73",
          4054 => x"38",
          4055 => x"08",
          4056 => x"08",
          4057 => x"82",
          4058 => x"ff",
          4059 => x"82",
          4060 => x"54",
          4061 => x"94",
          4062 => x"d4",
          4063 => x"d8",
          4064 => x"52",
          4065 => x"51",
          4066 => x"3f",
          4067 => x"33",
          4068 => x"2e",
          4069 => x"b3",
          4070 => x"b3",
          4071 => x"54",
          4072 => x"90",
          4073 => x"b1",
          4074 => x"9b",
          4075 => x"80",
          4076 => x"82",
          4077 => x"52",
          4078 => x"51",
          4079 => x"3f",
          4080 => x"33",
          4081 => x"2e",
          4082 => x"b4",
          4083 => x"82",
          4084 => x"ff",
          4085 => x"82",
          4086 => x"54",
          4087 => x"8e",
          4088 => x"9e",
          4089 => x"a6",
          4090 => x"93",
          4091 => x"b4",
          4092 => x"73",
          4093 => x"38",
          4094 => x"51",
          4095 => x"3f",
          4096 => x"33",
          4097 => x"2e",
          4098 => x"a7",
          4099 => x"ba",
          4100 => x"b4",
          4101 => x"73",
          4102 => x"38",
          4103 => x"51",
          4104 => x"3f",
          4105 => x"33",
          4106 => x"2e",
          4107 => x"a7",
          4108 => x"ba",
          4109 => x"b4",
          4110 => x"73",
          4111 => x"38",
          4112 => x"51",
          4113 => x"3f",
          4114 => x"51",
          4115 => x"3f",
          4116 => x"08",
          4117 => x"dc",
          4118 => x"fd",
          4119 => x"f8",
          4120 => x"a8",
          4121 => x"92",
          4122 => x"b3",
          4123 => x"82",
          4124 => x"ff",
          4125 => x"82",
          4126 => x"ff",
          4127 => x"82",
          4128 => x"52",
          4129 => x"51",
          4130 => x"3f",
          4131 => x"08",
          4132 => x"c0",
          4133 => x"d1",
          4134 => x"b5",
          4135 => x"84",
          4136 => x"71",
          4137 => x"82",
          4138 => x"52",
          4139 => x"51",
          4140 => x"3f",
          4141 => x"33",
          4142 => x"2e",
          4143 => x"b4",
          4144 => x"bd",
          4145 => x"75",
          4146 => x"3f",
          4147 => x"08",
          4148 => x"29",
          4149 => x"54",
          4150 => x"a8",
          4151 => x"a9",
          4152 => x"91",
          4153 => x"b4",
          4154 => x"73",
          4155 => x"38",
          4156 => x"08",
          4157 => x"c0",
          4158 => x"d0",
          4159 => x"b5",
          4160 => x"84",
          4161 => x"71",
          4162 => x"82",
          4163 => x"52",
          4164 => x"51",
          4165 => x"3f",
          4166 => x"51",
          4167 => x"3f",
          4168 => x"04",
          4169 => x"02",
          4170 => x"ff",
          4171 => x"84",
          4172 => x"71",
          4173 => x"95",
          4174 => x"71",
          4175 => x"aa",
          4176 => x"39",
          4177 => x"51",
          4178 => x"aa",
          4179 => x"39",
          4180 => x"51",
          4181 => x"aa",
          4182 => x"39",
          4183 => x"51",
          4184 => x"3f",
          4185 => x"04",
          4186 => x"0c",
          4187 => x"87",
          4188 => x"0c",
          4189 => x"a4",
          4190 => x"96",
          4191 => x"fd",
          4192 => x"98",
          4193 => x"2c",
          4194 => x"70",
          4195 => x"10",
          4196 => x"2b",
          4197 => x"54",
          4198 => x"0b",
          4199 => x"12",
          4200 => x"71",
          4201 => x"38",
          4202 => x"11",
          4203 => x"84",
          4204 => x"33",
          4205 => x"52",
          4206 => x"2e",
          4207 => x"83",
          4208 => x"72",
          4209 => x"0c",
          4210 => x"04",
          4211 => x"78",
          4212 => x"9f",
          4213 => x"33",
          4214 => x"71",
          4215 => x"38",
          4216 => x"ba",
          4217 => x"51",
          4218 => x"3f",
          4219 => x"ba",
          4220 => x"33",
          4221 => x"71",
          4222 => x"81",
          4223 => x"db",
          4224 => x"ff",
          4225 => x"73",
          4226 => x"3d",
          4227 => x"3d",
          4228 => x"84",
          4229 => x"33",
          4230 => x"bb",
          4231 => x"b5",
          4232 => x"84",
          4233 => x"a8",
          4234 => x"51",
          4235 => x"58",
          4236 => x"2e",
          4237 => x"51",
          4238 => x"82",
          4239 => x"70",
          4240 => x"b4",
          4241 => x"19",
          4242 => x"56",
          4243 => x"3f",
          4244 => x"08",
          4245 => x"b5",
          4246 => x"84",
          4247 => x"a8",
          4248 => x"51",
          4249 => x"80",
          4250 => x"75",
          4251 => x"74",
          4252 => x"3f",
          4253 => x"33",
          4254 => x"74",
          4255 => x"34",
          4256 => x"06",
          4257 => x"27",
          4258 => x"0b",
          4259 => x"34",
          4260 => x"b6",
          4261 => x"fc",
          4262 => x"80",
          4263 => x"82",
          4264 => x"55",
          4265 => x"8c",
          4266 => x"54",
          4267 => x"52",
          4268 => x"d9",
          4269 => x"b4",
          4270 => x"8a",
          4271 => x"ce",
          4272 => x"fc",
          4273 => x"dd",
          4274 => x"3d",
          4275 => x"3d",
          4276 => x"a8",
          4277 => x"72",
          4278 => x"80",
          4279 => x"71",
          4280 => x"3f",
          4281 => x"ff",
          4282 => x"54",
          4283 => x"25",
          4284 => x"0b",
          4285 => x"34",
          4286 => x"08",
          4287 => x"2e",
          4288 => x"51",
          4289 => x"3f",
          4290 => x"08",
          4291 => x"3f",
          4292 => x"b4",
          4293 => x"3d",
          4294 => x"3d",
          4295 => x"80",
          4296 => x"fc",
          4297 => x"e2",
          4298 => x"b5",
          4299 => x"d2",
          4300 => x"fc",
          4301 => x"f8",
          4302 => x"70",
          4303 => x"8b",
          4304 => x"b5",
          4305 => x"2e",
          4306 => x"51",
          4307 => x"82",
          4308 => x"55",
          4309 => x"b5",
          4310 => x"9d",
          4311 => x"a8",
          4312 => x"70",
          4313 => x"80",
          4314 => x"53",
          4315 => x"17",
          4316 => x"52",
          4317 => x"e1",
          4318 => x"2e",
          4319 => x"ff",
          4320 => x"3d",
          4321 => x"3d",
          4322 => x"08",
          4323 => x"5a",
          4324 => x"58",
          4325 => x"82",
          4326 => x"51",
          4327 => x"3f",
          4328 => x"08",
          4329 => x"ff",
          4330 => x"fc",
          4331 => x"80",
          4332 => x"3d",
          4333 => x"81",
          4334 => x"82",
          4335 => x"80",
          4336 => x"75",
          4337 => x"e0",
          4338 => x"a8",
          4339 => x"58",
          4340 => x"82",
          4341 => x"25",
          4342 => x"b5",
          4343 => x"05",
          4344 => x"55",
          4345 => x"74",
          4346 => x"70",
          4347 => x"2a",
          4348 => x"78",
          4349 => x"38",
          4350 => x"38",
          4351 => x"08",
          4352 => x"53",
          4353 => x"8c",
          4354 => x"a8",
          4355 => x"89",
          4356 => x"b4",
          4357 => x"ee",
          4358 => x"2e",
          4359 => x"9b",
          4360 => x"79",
          4361 => x"ee",
          4362 => x"ff",
          4363 => x"ab",
          4364 => x"82",
          4365 => x"74",
          4366 => x"77",
          4367 => x"0c",
          4368 => x"04",
          4369 => x"7c",
          4370 => x"71",
          4371 => x"59",
          4372 => x"a0",
          4373 => x"06",
          4374 => x"33",
          4375 => x"77",
          4376 => x"38",
          4377 => x"5b",
          4378 => x"56",
          4379 => x"a0",
          4380 => x"06",
          4381 => x"75",
          4382 => x"80",
          4383 => x"29",
          4384 => x"05",
          4385 => x"55",
          4386 => x"3f",
          4387 => x"08",
          4388 => x"74",
          4389 => x"9d",
          4390 => x"a8",
          4391 => x"38",
          4392 => x"55",
          4393 => x"88",
          4394 => x"2e",
          4395 => x"39",
          4396 => x"ad",
          4397 => x"5a",
          4398 => x"11",
          4399 => x"51",
          4400 => x"3f",
          4401 => x"08",
          4402 => x"38",
          4403 => x"78",
          4404 => x"fd",
          4405 => x"b5",
          4406 => x"ff",
          4407 => x"85",
          4408 => x"91",
          4409 => x"70",
          4410 => x"51",
          4411 => x"27",
          4412 => x"80",
          4413 => x"b5",
          4414 => x"3d",
          4415 => x"3d",
          4416 => x"08",
          4417 => x"b4",
          4418 => x"5f",
          4419 => x"af",
          4420 => x"b5",
          4421 => x"b4",
          4422 => x"5b",
          4423 => x"38",
          4424 => x"f8",
          4425 => x"73",
          4426 => x"55",
          4427 => x"81",
          4428 => x"70",
          4429 => x"56",
          4430 => x"81",
          4431 => x"51",
          4432 => x"82",
          4433 => x"82",
          4434 => x"82",
          4435 => x"80",
          4436 => x"38",
          4437 => x"52",
          4438 => x"08",
          4439 => x"b4",
          4440 => x"a8",
          4441 => x"8c",
          4442 => x"e0",
          4443 => x"96",
          4444 => x"39",
          4445 => x"08",
          4446 => x"fc",
          4447 => x"f8",
          4448 => x"70",
          4449 => x"86",
          4450 => x"b5",
          4451 => x"82",
          4452 => x"74",
          4453 => x"06",
          4454 => x"82",
          4455 => x"51",
          4456 => x"3f",
          4457 => x"08",
          4458 => x"82",
          4459 => x"25",
          4460 => x"b5",
          4461 => x"05",
          4462 => x"55",
          4463 => x"80",
          4464 => x"ff",
          4465 => x"51",
          4466 => x"81",
          4467 => x"ff",
          4468 => x"93",
          4469 => x"38",
          4470 => x"ff",
          4471 => x"06",
          4472 => x"86",
          4473 => x"b4",
          4474 => x"8c",
          4475 => x"fc",
          4476 => x"84",
          4477 => x"3f",
          4478 => x"ec",
          4479 => x"b5",
          4480 => x"2b",
          4481 => x"51",
          4482 => x"2e",
          4483 => x"81",
          4484 => x"cc",
          4485 => x"98",
          4486 => x"2c",
          4487 => x"33",
          4488 => x"70",
          4489 => x"98",
          4490 => x"84",
          4491 => x"b4",
          4492 => x"15",
          4493 => x"51",
          4494 => x"59",
          4495 => x"58",
          4496 => x"78",
          4497 => x"38",
          4498 => x"b4",
          4499 => x"80",
          4500 => x"ff",
          4501 => x"98",
          4502 => x"80",
          4503 => x"ce",
          4504 => x"74",
          4505 => x"f6",
          4506 => x"b5",
          4507 => x"ff",
          4508 => x"80",
          4509 => x"74",
          4510 => x"34",
          4511 => x"39",
          4512 => x"0a",
          4513 => x"0a",
          4514 => x"2c",
          4515 => x"06",
          4516 => x"73",
          4517 => x"38",
          4518 => x"52",
          4519 => x"df",
          4520 => x"a8",
          4521 => x"06",
          4522 => x"38",
          4523 => x"56",
          4524 => x"80",
          4525 => x"1c",
          4526 => x"cc",
          4527 => x"98",
          4528 => x"2c",
          4529 => x"33",
          4530 => x"70",
          4531 => x"10",
          4532 => x"2b",
          4533 => x"11",
          4534 => x"51",
          4535 => x"51",
          4536 => x"2e",
          4537 => x"fe",
          4538 => x"aa",
          4539 => x"7d",
          4540 => x"82",
          4541 => x"80",
          4542 => x"d0",
          4543 => x"75",
          4544 => x"34",
          4545 => x"d0",
          4546 => x"3d",
          4547 => x"0c",
          4548 => x"95",
          4549 => x"38",
          4550 => x"82",
          4551 => x"54",
          4552 => x"82",
          4553 => x"54",
          4554 => x"fd",
          4555 => x"cc",
          4556 => x"73",
          4557 => x"38",
          4558 => x"70",
          4559 => x"55",
          4560 => x"9e",
          4561 => x"54",
          4562 => x"15",
          4563 => x"80",
          4564 => x"ff",
          4565 => x"98",
          4566 => x"dc",
          4567 => x"55",
          4568 => x"cc",
          4569 => x"11",
          4570 => x"82",
          4571 => x"73",
          4572 => x"3d",
          4573 => x"82",
          4574 => x"54",
          4575 => x"89",
          4576 => x"54",
          4577 => x"d8",
          4578 => x"dc",
          4579 => x"80",
          4580 => x"ff",
          4581 => x"98",
          4582 => x"d8",
          4583 => x"56",
          4584 => x"25",
          4585 => x"1a",
          4586 => x"54",
          4587 => x"3f",
          4588 => x"0a",
          4589 => x"0a",
          4590 => x"2c",
          4591 => x"33",
          4592 => x"73",
          4593 => x"38",
          4594 => x"33",
          4595 => x"70",
          4596 => x"cc",
          4597 => x"51",
          4598 => x"77",
          4599 => x"38",
          4600 => x"ae",
          4601 => x"81",
          4602 => x"81",
          4603 => x"70",
          4604 => x"cc",
          4605 => x"51",
          4606 => x"24",
          4607 => x"f8",
          4608 => x"34",
          4609 => x"1b",
          4610 => x"dc",
          4611 => x"82",
          4612 => x"f3",
          4613 => x"e4",
          4614 => x"dc",
          4615 => x"ff",
          4616 => x"73",
          4617 => x"d0",
          4618 => x"d8",
          4619 => x"54",
          4620 => x"d8",
          4621 => x"54",
          4622 => x"dc",
          4623 => x"ff",
          4624 => x"82",
          4625 => x"70",
          4626 => x"98",
          4627 => x"d8",
          4628 => x"56",
          4629 => x"25",
          4630 => x"1a",
          4631 => x"33",
          4632 => x"33",
          4633 => x"c0",
          4634 => x"80",
          4635 => x"80",
          4636 => x"98",
          4637 => x"d8",
          4638 => x"55",
          4639 => x"da",
          4640 => x"ff",
          4641 => x"82",
          4642 => x"70",
          4643 => x"98",
          4644 => x"d8",
          4645 => x"56",
          4646 => x"24",
          4647 => x"88",
          4648 => x"84",
          4649 => x"80",
          4650 => x"80",
          4651 => x"98",
          4652 => x"d8",
          4653 => x"55",
          4654 => x"e3",
          4655 => x"39",
          4656 => x"33",
          4657 => x"80",
          4658 => x"51",
          4659 => x"3f",
          4660 => x"52",
          4661 => x"ec",
          4662 => x"a8",
          4663 => x"06",
          4664 => x"38",
          4665 => x"33",
          4666 => x"2e",
          4667 => x"53",
          4668 => x"51",
          4669 => x"84",
          4670 => x"34",
          4671 => x"cc",
          4672 => x"0b",
          4673 => x"34",
          4674 => x"a8",
          4675 => x"0d",
          4676 => x"dc",
          4677 => x"80",
          4678 => x"38",
          4679 => x"ac",
          4680 => x"cc",
          4681 => x"05",
          4682 => x"cc",
          4683 => x"81",
          4684 => x"e2",
          4685 => x"dc",
          4686 => x"d8",
          4687 => x"73",
          4688 => x"b4",
          4689 => x"54",
          4690 => x"d8",
          4691 => x"2b",
          4692 => x"75",
          4693 => x"56",
          4694 => x"74",
          4695 => x"74",
          4696 => x"14",
          4697 => x"73",
          4698 => x"ab",
          4699 => x"81",
          4700 => x"81",
          4701 => x"70",
          4702 => x"cc",
          4703 => x"51",
          4704 => x"24",
          4705 => x"51",
          4706 => x"3f",
          4707 => x"33",
          4708 => x"70",
          4709 => x"cc",
          4710 => x"51",
          4711 => x"74",
          4712 => x"38",
          4713 => x"aa",
          4714 => x"81",
          4715 => x"81",
          4716 => x"70",
          4717 => x"cc",
          4718 => x"51",
          4719 => x"25",
          4720 => x"b4",
          4721 => x"dc",
          4722 => x"ff",
          4723 => x"d8",
          4724 => x"54",
          4725 => x"f8",
          4726 => x"14",
          4727 => x"cc",
          4728 => x"1a",
          4729 => x"54",
          4730 => x"3f",
          4731 => x"33",
          4732 => x"06",
          4733 => x"33",
          4734 => x"75",
          4735 => x"38",
          4736 => x"82",
          4737 => x"80",
          4738 => x"f0",
          4739 => x"3f",
          4740 => x"cc",
          4741 => x"0b",
          4742 => x"34",
          4743 => x"7a",
          4744 => x"b4",
          4745 => x"74",
          4746 => x"38",
          4747 => x"b2",
          4748 => x"b5",
          4749 => x"cc",
          4750 => x"b5",
          4751 => x"ff",
          4752 => x"53",
          4753 => x"51",
          4754 => x"3f",
          4755 => x"c0",
          4756 => x"29",
          4757 => x"05",
          4758 => x"56",
          4759 => x"2e",
          4760 => x"51",
          4761 => x"3f",
          4762 => x"08",
          4763 => x"34",
          4764 => x"08",
          4765 => x"81",
          4766 => x"52",
          4767 => x"b4",
          4768 => x"1b",
          4769 => x"39",
          4770 => x"74",
          4771 => x"e8",
          4772 => x"ff",
          4773 => x"99",
          4774 => x"2e",
          4775 => x"ae",
          4776 => x"a8",
          4777 => x"80",
          4778 => x"74",
          4779 => x"f8",
          4780 => x"a8",
          4781 => x"d8",
          4782 => x"a8",
          4783 => x"06",
          4784 => x"74",
          4785 => x"ff",
          4786 => x"80",
          4787 => x"84",
          4788 => x"ac",
          4789 => x"56",
          4790 => x"2e",
          4791 => x"51",
          4792 => x"3f",
          4793 => x"08",
          4794 => x"34",
          4795 => x"08",
          4796 => x"81",
          4797 => x"52",
          4798 => x"b3",
          4799 => x"1b",
          4800 => x"ff",
          4801 => x"39",
          4802 => x"d8",
          4803 => x"34",
          4804 => x"53",
          4805 => x"33",
          4806 => x"ed",
          4807 => x"d8",
          4808 => x"dc",
          4809 => x"ff",
          4810 => x"d8",
          4811 => x"54",
          4812 => x"f5",
          4813 => x"14",
          4814 => x"cc",
          4815 => x"1a",
          4816 => x"54",
          4817 => x"3f",
          4818 => x"82",
          4819 => x"54",
          4820 => x"f5",
          4821 => x"51",
          4822 => x"3f",
          4823 => x"33",
          4824 => x"73",
          4825 => x"34",
          4826 => x"f9",
          4827 => x"df",
          4828 => x"b5",
          4829 => x"80",
          4830 => x"9c",
          4831 => x"53",
          4832 => x"df",
          4833 => x"b7",
          4834 => x"b5",
          4835 => x"80",
          4836 => x"34",
          4837 => x"81",
          4838 => x"b5",
          4839 => x"77",
          4840 => x"76",
          4841 => x"82",
          4842 => x"54",
          4843 => x"34",
          4844 => x"34",
          4845 => x"08",
          4846 => x"22",
          4847 => x"80",
          4848 => x"83",
          4849 => x"70",
          4850 => x"51",
          4851 => x"88",
          4852 => x"89",
          4853 => x"b5",
          4854 => x"88",
          4855 => x"a0",
          4856 => x"11",
          4857 => x"77",
          4858 => x"76",
          4859 => x"89",
          4860 => x"ff",
          4861 => x"52",
          4862 => x"72",
          4863 => x"fb",
          4864 => x"82",
          4865 => x"ff",
          4866 => x"51",
          4867 => x"b5",
          4868 => x"3d",
          4869 => x"3d",
          4870 => x"05",
          4871 => x"05",
          4872 => x"71",
          4873 => x"a0",
          4874 => x"2b",
          4875 => x"83",
          4876 => x"70",
          4877 => x"33",
          4878 => x"07",
          4879 => x"ae",
          4880 => x"81",
          4881 => x"07",
          4882 => x"53",
          4883 => x"54",
          4884 => x"53",
          4885 => x"77",
          4886 => x"18",
          4887 => x"a0",
          4888 => x"88",
          4889 => x"70",
          4890 => x"74",
          4891 => x"82",
          4892 => x"70",
          4893 => x"81",
          4894 => x"88",
          4895 => x"83",
          4896 => x"f8",
          4897 => x"56",
          4898 => x"73",
          4899 => x"06",
          4900 => x"54",
          4901 => x"82",
          4902 => x"81",
          4903 => x"72",
          4904 => x"82",
          4905 => x"16",
          4906 => x"34",
          4907 => x"34",
          4908 => x"04",
          4909 => x"82",
          4910 => x"02",
          4911 => x"05",
          4912 => x"2b",
          4913 => x"11",
          4914 => x"33",
          4915 => x"71",
          4916 => x"58",
          4917 => x"55",
          4918 => x"84",
          4919 => x"13",
          4920 => x"2b",
          4921 => x"2a",
          4922 => x"52",
          4923 => x"34",
          4924 => x"34",
          4925 => x"08",
          4926 => x"11",
          4927 => x"33",
          4928 => x"71",
          4929 => x"56",
          4930 => x"72",
          4931 => x"33",
          4932 => x"71",
          4933 => x"70",
          4934 => x"56",
          4935 => x"86",
          4936 => x"87",
          4937 => x"b5",
          4938 => x"70",
          4939 => x"33",
          4940 => x"07",
          4941 => x"ff",
          4942 => x"2a",
          4943 => x"53",
          4944 => x"34",
          4945 => x"34",
          4946 => x"04",
          4947 => x"02",
          4948 => x"82",
          4949 => x"71",
          4950 => x"11",
          4951 => x"12",
          4952 => x"2b",
          4953 => x"29",
          4954 => x"81",
          4955 => x"98",
          4956 => x"2b",
          4957 => x"53",
          4958 => x"56",
          4959 => x"71",
          4960 => x"f6",
          4961 => x"fe",
          4962 => x"b5",
          4963 => x"16",
          4964 => x"12",
          4965 => x"2b",
          4966 => x"07",
          4967 => x"33",
          4968 => x"71",
          4969 => x"70",
          4970 => x"ff",
          4971 => x"52",
          4972 => x"5a",
          4973 => x"05",
          4974 => x"54",
          4975 => x"13",
          4976 => x"13",
          4977 => x"a0",
          4978 => x"70",
          4979 => x"33",
          4980 => x"71",
          4981 => x"56",
          4982 => x"72",
          4983 => x"81",
          4984 => x"88",
          4985 => x"81",
          4986 => x"70",
          4987 => x"51",
          4988 => x"72",
          4989 => x"81",
          4990 => x"3d",
          4991 => x"3d",
          4992 => x"a0",
          4993 => x"05",
          4994 => x"70",
          4995 => x"11",
          4996 => x"83",
          4997 => x"8b",
          4998 => x"2b",
          4999 => x"59",
          5000 => x"73",
          5001 => x"81",
          5002 => x"88",
          5003 => x"8c",
          5004 => x"22",
          5005 => x"88",
          5006 => x"53",
          5007 => x"73",
          5008 => x"14",
          5009 => x"a0",
          5010 => x"70",
          5011 => x"33",
          5012 => x"71",
          5013 => x"56",
          5014 => x"72",
          5015 => x"33",
          5016 => x"71",
          5017 => x"70",
          5018 => x"55",
          5019 => x"82",
          5020 => x"83",
          5021 => x"b5",
          5022 => x"82",
          5023 => x"12",
          5024 => x"2b",
          5025 => x"a8",
          5026 => x"87",
          5027 => x"f7",
          5028 => x"82",
          5029 => x"31",
          5030 => x"83",
          5031 => x"70",
          5032 => x"fd",
          5033 => x"b5",
          5034 => x"83",
          5035 => x"82",
          5036 => x"12",
          5037 => x"2b",
          5038 => x"07",
          5039 => x"33",
          5040 => x"71",
          5041 => x"90",
          5042 => x"42",
          5043 => x"5b",
          5044 => x"54",
          5045 => x"8d",
          5046 => x"80",
          5047 => x"fe",
          5048 => x"84",
          5049 => x"33",
          5050 => x"71",
          5051 => x"83",
          5052 => x"11",
          5053 => x"53",
          5054 => x"55",
          5055 => x"34",
          5056 => x"06",
          5057 => x"14",
          5058 => x"a0",
          5059 => x"84",
          5060 => x"13",
          5061 => x"2b",
          5062 => x"2a",
          5063 => x"56",
          5064 => x"16",
          5065 => x"16",
          5066 => x"a0",
          5067 => x"80",
          5068 => x"34",
          5069 => x"14",
          5070 => x"a0",
          5071 => x"84",
          5072 => x"85",
          5073 => x"b5",
          5074 => x"70",
          5075 => x"33",
          5076 => x"07",
          5077 => x"80",
          5078 => x"2a",
          5079 => x"56",
          5080 => x"34",
          5081 => x"34",
          5082 => x"04",
          5083 => x"73",
          5084 => x"a0",
          5085 => x"f7",
          5086 => x"80",
          5087 => x"71",
          5088 => x"3f",
          5089 => x"04",
          5090 => x"80",
          5091 => x"f8",
          5092 => x"b5",
          5093 => x"ff",
          5094 => x"b5",
          5095 => x"11",
          5096 => x"33",
          5097 => x"07",
          5098 => x"56",
          5099 => x"ff",
          5100 => x"78",
          5101 => x"38",
          5102 => x"17",
          5103 => x"12",
          5104 => x"2b",
          5105 => x"ff",
          5106 => x"31",
          5107 => x"ff",
          5108 => x"27",
          5109 => x"56",
          5110 => x"79",
          5111 => x"73",
          5112 => x"38",
          5113 => x"5b",
          5114 => x"85",
          5115 => x"88",
          5116 => x"54",
          5117 => x"78",
          5118 => x"2e",
          5119 => x"79",
          5120 => x"76",
          5121 => x"b5",
          5122 => x"70",
          5123 => x"33",
          5124 => x"07",
          5125 => x"ff",
          5126 => x"5a",
          5127 => x"73",
          5128 => x"38",
          5129 => x"54",
          5130 => x"81",
          5131 => x"54",
          5132 => x"81",
          5133 => x"7a",
          5134 => x"06",
          5135 => x"51",
          5136 => x"81",
          5137 => x"80",
          5138 => x"52",
          5139 => x"c6",
          5140 => x"a0",
          5141 => x"86",
          5142 => x"12",
          5143 => x"2b",
          5144 => x"07",
          5145 => x"55",
          5146 => x"17",
          5147 => x"ff",
          5148 => x"2a",
          5149 => x"54",
          5150 => x"34",
          5151 => x"06",
          5152 => x"15",
          5153 => x"a0",
          5154 => x"2b",
          5155 => x"1e",
          5156 => x"87",
          5157 => x"88",
          5158 => x"88",
          5159 => x"5e",
          5160 => x"54",
          5161 => x"34",
          5162 => x"34",
          5163 => x"08",
          5164 => x"11",
          5165 => x"33",
          5166 => x"71",
          5167 => x"53",
          5168 => x"74",
          5169 => x"86",
          5170 => x"87",
          5171 => x"b5",
          5172 => x"16",
          5173 => x"11",
          5174 => x"33",
          5175 => x"07",
          5176 => x"53",
          5177 => x"56",
          5178 => x"16",
          5179 => x"16",
          5180 => x"a0",
          5181 => x"05",
          5182 => x"b5",
          5183 => x"3d",
          5184 => x"3d",
          5185 => x"82",
          5186 => x"84",
          5187 => x"3f",
          5188 => x"80",
          5189 => x"71",
          5190 => x"3f",
          5191 => x"08",
          5192 => x"b5",
          5193 => x"3d",
          5194 => x"3d",
          5195 => x"40",
          5196 => x"42",
          5197 => x"a0",
          5198 => x"09",
          5199 => x"38",
          5200 => x"7b",
          5201 => x"51",
          5202 => x"82",
          5203 => x"54",
          5204 => x"7e",
          5205 => x"51",
          5206 => x"7e",
          5207 => x"39",
          5208 => x"8f",
          5209 => x"a8",
          5210 => x"ff",
          5211 => x"a0",
          5212 => x"31",
          5213 => x"83",
          5214 => x"70",
          5215 => x"11",
          5216 => x"12",
          5217 => x"2b",
          5218 => x"31",
          5219 => x"ff",
          5220 => x"29",
          5221 => x"88",
          5222 => x"33",
          5223 => x"71",
          5224 => x"70",
          5225 => x"44",
          5226 => x"41",
          5227 => x"5b",
          5228 => x"5b",
          5229 => x"25",
          5230 => x"81",
          5231 => x"75",
          5232 => x"ff",
          5233 => x"54",
          5234 => x"83",
          5235 => x"88",
          5236 => x"88",
          5237 => x"33",
          5238 => x"71",
          5239 => x"90",
          5240 => x"47",
          5241 => x"54",
          5242 => x"8b",
          5243 => x"31",
          5244 => x"ff",
          5245 => x"77",
          5246 => x"fe",
          5247 => x"54",
          5248 => x"09",
          5249 => x"38",
          5250 => x"c0",
          5251 => x"ff",
          5252 => x"81",
          5253 => x"8e",
          5254 => x"24",
          5255 => x"51",
          5256 => x"81",
          5257 => x"18",
          5258 => x"24",
          5259 => x"79",
          5260 => x"33",
          5261 => x"71",
          5262 => x"53",
          5263 => x"f4",
          5264 => x"78",
          5265 => x"3f",
          5266 => x"08",
          5267 => x"06",
          5268 => x"53",
          5269 => x"82",
          5270 => x"11",
          5271 => x"55",
          5272 => x"da",
          5273 => x"a0",
          5274 => x"05",
          5275 => x"ff",
          5276 => x"81",
          5277 => x"15",
          5278 => x"24",
          5279 => x"78",
          5280 => x"3f",
          5281 => x"08",
          5282 => x"33",
          5283 => x"71",
          5284 => x"53",
          5285 => x"9c",
          5286 => x"78",
          5287 => x"3f",
          5288 => x"08",
          5289 => x"06",
          5290 => x"53",
          5291 => x"82",
          5292 => x"11",
          5293 => x"55",
          5294 => x"82",
          5295 => x"a0",
          5296 => x"05",
          5297 => x"19",
          5298 => x"83",
          5299 => x"58",
          5300 => x"7f",
          5301 => x"b0",
          5302 => x"a8",
          5303 => x"b5",
          5304 => x"2e",
          5305 => x"53",
          5306 => x"b5",
          5307 => x"ff",
          5308 => x"73",
          5309 => x"3f",
          5310 => x"78",
          5311 => x"80",
          5312 => x"78",
          5313 => x"3f",
          5314 => x"2b",
          5315 => x"08",
          5316 => x"51",
          5317 => x"7b",
          5318 => x"b5",
          5319 => x"3d",
          5320 => x"3d",
          5321 => x"29",
          5322 => x"fb",
          5323 => x"b5",
          5324 => x"82",
          5325 => x"80",
          5326 => x"73",
          5327 => x"82",
          5328 => x"51",
          5329 => x"3f",
          5330 => x"a8",
          5331 => x"0d",
          5332 => x"0d",
          5333 => x"33",
          5334 => x"70",
          5335 => x"38",
          5336 => x"11",
          5337 => x"82",
          5338 => x"83",
          5339 => x"fc",
          5340 => x"9b",
          5341 => x"84",
          5342 => x"33",
          5343 => x"51",
          5344 => x"80",
          5345 => x"84",
          5346 => x"92",
          5347 => x"51",
          5348 => x"80",
          5349 => x"81",
          5350 => x"72",
          5351 => x"92",
          5352 => x"81",
          5353 => x"0b",
          5354 => x"8c",
          5355 => x"71",
          5356 => x"06",
          5357 => x"80",
          5358 => x"87",
          5359 => x"08",
          5360 => x"38",
          5361 => x"80",
          5362 => x"71",
          5363 => x"c0",
          5364 => x"51",
          5365 => x"87",
          5366 => x"b5",
          5367 => x"82",
          5368 => x"33",
          5369 => x"b5",
          5370 => x"3d",
          5371 => x"3d",
          5372 => x"64",
          5373 => x"bf",
          5374 => x"40",
          5375 => x"74",
          5376 => x"cd",
          5377 => x"a8",
          5378 => x"7a",
          5379 => x"81",
          5380 => x"72",
          5381 => x"87",
          5382 => x"11",
          5383 => x"8c",
          5384 => x"92",
          5385 => x"5a",
          5386 => x"58",
          5387 => x"c0",
          5388 => x"76",
          5389 => x"76",
          5390 => x"70",
          5391 => x"81",
          5392 => x"54",
          5393 => x"8e",
          5394 => x"52",
          5395 => x"81",
          5396 => x"81",
          5397 => x"74",
          5398 => x"53",
          5399 => x"83",
          5400 => x"78",
          5401 => x"8f",
          5402 => x"2e",
          5403 => x"c0",
          5404 => x"52",
          5405 => x"87",
          5406 => x"08",
          5407 => x"2e",
          5408 => x"84",
          5409 => x"38",
          5410 => x"87",
          5411 => x"15",
          5412 => x"70",
          5413 => x"52",
          5414 => x"ff",
          5415 => x"39",
          5416 => x"81",
          5417 => x"ff",
          5418 => x"57",
          5419 => x"90",
          5420 => x"80",
          5421 => x"71",
          5422 => x"78",
          5423 => x"38",
          5424 => x"80",
          5425 => x"80",
          5426 => x"81",
          5427 => x"72",
          5428 => x"0c",
          5429 => x"04",
          5430 => x"60",
          5431 => x"8c",
          5432 => x"33",
          5433 => x"5b",
          5434 => x"74",
          5435 => x"e1",
          5436 => x"a8",
          5437 => x"79",
          5438 => x"78",
          5439 => x"06",
          5440 => x"77",
          5441 => x"87",
          5442 => x"11",
          5443 => x"8c",
          5444 => x"92",
          5445 => x"59",
          5446 => x"85",
          5447 => x"98",
          5448 => x"7d",
          5449 => x"0c",
          5450 => x"08",
          5451 => x"70",
          5452 => x"53",
          5453 => x"2e",
          5454 => x"70",
          5455 => x"33",
          5456 => x"18",
          5457 => x"2a",
          5458 => x"51",
          5459 => x"2e",
          5460 => x"c0",
          5461 => x"52",
          5462 => x"87",
          5463 => x"08",
          5464 => x"2e",
          5465 => x"84",
          5466 => x"38",
          5467 => x"87",
          5468 => x"15",
          5469 => x"70",
          5470 => x"52",
          5471 => x"ff",
          5472 => x"39",
          5473 => x"81",
          5474 => x"80",
          5475 => x"52",
          5476 => x"90",
          5477 => x"80",
          5478 => x"71",
          5479 => x"7a",
          5480 => x"38",
          5481 => x"80",
          5482 => x"80",
          5483 => x"81",
          5484 => x"72",
          5485 => x"0c",
          5486 => x"04",
          5487 => x"7a",
          5488 => x"a3",
          5489 => x"88",
          5490 => x"33",
          5491 => x"56",
          5492 => x"3f",
          5493 => x"08",
          5494 => x"83",
          5495 => x"fe",
          5496 => x"87",
          5497 => x"0c",
          5498 => x"76",
          5499 => x"38",
          5500 => x"93",
          5501 => x"2b",
          5502 => x"8c",
          5503 => x"71",
          5504 => x"38",
          5505 => x"71",
          5506 => x"c6",
          5507 => x"39",
          5508 => x"81",
          5509 => x"06",
          5510 => x"71",
          5511 => x"38",
          5512 => x"8c",
          5513 => x"e8",
          5514 => x"98",
          5515 => x"71",
          5516 => x"73",
          5517 => x"92",
          5518 => x"72",
          5519 => x"06",
          5520 => x"f7",
          5521 => x"80",
          5522 => x"88",
          5523 => x"0c",
          5524 => x"80",
          5525 => x"56",
          5526 => x"56",
          5527 => x"82",
          5528 => x"88",
          5529 => x"fe",
          5530 => x"81",
          5531 => x"33",
          5532 => x"07",
          5533 => x"0c",
          5534 => x"3d",
          5535 => x"3d",
          5536 => x"11",
          5537 => x"33",
          5538 => x"71",
          5539 => x"81",
          5540 => x"72",
          5541 => x"75",
          5542 => x"82",
          5543 => x"52",
          5544 => x"54",
          5545 => x"0d",
          5546 => x"0d",
          5547 => x"05",
          5548 => x"52",
          5549 => x"70",
          5550 => x"34",
          5551 => x"51",
          5552 => x"83",
          5553 => x"ff",
          5554 => x"75",
          5555 => x"72",
          5556 => x"54",
          5557 => x"2a",
          5558 => x"70",
          5559 => x"34",
          5560 => x"51",
          5561 => x"81",
          5562 => x"70",
          5563 => x"70",
          5564 => x"3d",
          5565 => x"3d",
          5566 => x"77",
          5567 => x"70",
          5568 => x"38",
          5569 => x"05",
          5570 => x"70",
          5571 => x"34",
          5572 => x"eb",
          5573 => x"0d",
          5574 => x"0d",
          5575 => x"54",
          5576 => x"72",
          5577 => x"54",
          5578 => x"51",
          5579 => x"84",
          5580 => x"fc",
          5581 => x"77",
          5582 => x"53",
          5583 => x"05",
          5584 => x"70",
          5585 => x"33",
          5586 => x"ff",
          5587 => x"52",
          5588 => x"2e",
          5589 => x"80",
          5590 => x"71",
          5591 => x"0c",
          5592 => x"04",
          5593 => x"74",
          5594 => x"89",
          5595 => x"2e",
          5596 => x"11",
          5597 => x"52",
          5598 => x"70",
          5599 => x"a8",
          5600 => x"0d",
          5601 => x"82",
          5602 => x"04",
          5603 => x"b5",
          5604 => x"f7",
          5605 => x"56",
          5606 => x"17",
          5607 => x"74",
          5608 => x"d6",
          5609 => x"b0",
          5610 => x"b4",
          5611 => x"81",
          5612 => x"59",
          5613 => x"82",
          5614 => x"7a",
          5615 => x"06",
          5616 => x"b5",
          5617 => x"17",
          5618 => x"08",
          5619 => x"08",
          5620 => x"08",
          5621 => x"74",
          5622 => x"38",
          5623 => x"55",
          5624 => x"09",
          5625 => x"38",
          5626 => x"18",
          5627 => x"81",
          5628 => x"f9",
          5629 => x"39",
          5630 => x"82",
          5631 => x"8b",
          5632 => x"fa",
          5633 => x"7a",
          5634 => x"57",
          5635 => x"08",
          5636 => x"75",
          5637 => x"3f",
          5638 => x"08",
          5639 => x"a8",
          5640 => x"81",
          5641 => x"b4",
          5642 => x"16",
          5643 => x"be",
          5644 => x"a8",
          5645 => x"85",
          5646 => x"81",
          5647 => x"17",
          5648 => x"b5",
          5649 => x"3d",
          5650 => x"3d",
          5651 => x"52",
          5652 => x"3f",
          5653 => x"08",
          5654 => x"a8",
          5655 => x"38",
          5656 => x"74",
          5657 => x"81",
          5658 => x"38",
          5659 => x"59",
          5660 => x"09",
          5661 => x"e3",
          5662 => x"53",
          5663 => x"08",
          5664 => x"70",
          5665 => x"91",
          5666 => x"d5",
          5667 => x"17",
          5668 => x"3f",
          5669 => x"a4",
          5670 => x"51",
          5671 => x"86",
          5672 => x"f2",
          5673 => x"17",
          5674 => x"3f",
          5675 => x"52",
          5676 => x"51",
          5677 => x"8c",
          5678 => x"84",
          5679 => x"fc",
          5680 => x"17",
          5681 => x"70",
          5682 => x"79",
          5683 => x"52",
          5684 => x"51",
          5685 => x"77",
          5686 => x"80",
          5687 => x"81",
          5688 => x"f9",
          5689 => x"b5",
          5690 => x"2e",
          5691 => x"58",
          5692 => x"a8",
          5693 => x"0d",
          5694 => x"0d",
          5695 => x"98",
          5696 => x"05",
          5697 => x"80",
          5698 => x"27",
          5699 => x"14",
          5700 => x"29",
          5701 => x"05",
          5702 => x"82",
          5703 => x"87",
          5704 => x"f9",
          5705 => x"7a",
          5706 => x"54",
          5707 => x"27",
          5708 => x"76",
          5709 => x"27",
          5710 => x"ff",
          5711 => x"58",
          5712 => x"80",
          5713 => x"82",
          5714 => x"72",
          5715 => x"38",
          5716 => x"72",
          5717 => x"8e",
          5718 => x"39",
          5719 => x"17",
          5720 => x"a4",
          5721 => x"53",
          5722 => x"fd",
          5723 => x"b5",
          5724 => x"9f",
          5725 => x"ff",
          5726 => x"11",
          5727 => x"70",
          5728 => x"18",
          5729 => x"76",
          5730 => x"53",
          5731 => x"82",
          5732 => x"80",
          5733 => x"83",
          5734 => x"b4",
          5735 => x"88",
          5736 => x"79",
          5737 => x"84",
          5738 => x"58",
          5739 => x"80",
          5740 => x"9f",
          5741 => x"80",
          5742 => x"88",
          5743 => x"08",
          5744 => x"51",
          5745 => x"82",
          5746 => x"80",
          5747 => x"10",
          5748 => x"74",
          5749 => x"51",
          5750 => x"82",
          5751 => x"83",
          5752 => x"58",
          5753 => x"87",
          5754 => x"08",
          5755 => x"51",
          5756 => x"82",
          5757 => x"9b",
          5758 => x"2b",
          5759 => x"74",
          5760 => x"51",
          5761 => x"82",
          5762 => x"f0",
          5763 => x"83",
          5764 => x"77",
          5765 => x"0c",
          5766 => x"04",
          5767 => x"7a",
          5768 => x"58",
          5769 => x"81",
          5770 => x"9e",
          5771 => x"17",
          5772 => x"96",
          5773 => x"53",
          5774 => x"81",
          5775 => x"79",
          5776 => x"72",
          5777 => x"38",
          5778 => x"72",
          5779 => x"b8",
          5780 => x"39",
          5781 => x"17",
          5782 => x"a4",
          5783 => x"53",
          5784 => x"fb",
          5785 => x"b5",
          5786 => x"82",
          5787 => x"81",
          5788 => x"83",
          5789 => x"b4",
          5790 => x"78",
          5791 => x"56",
          5792 => x"76",
          5793 => x"38",
          5794 => x"9f",
          5795 => x"33",
          5796 => x"07",
          5797 => x"74",
          5798 => x"83",
          5799 => x"89",
          5800 => x"08",
          5801 => x"51",
          5802 => x"82",
          5803 => x"59",
          5804 => x"08",
          5805 => x"74",
          5806 => x"16",
          5807 => x"84",
          5808 => x"76",
          5809 => x"88",
          5810 => x"81",
          5811 => x"8f",
          5812 => x"53",
          5813 => x"80",
          5814 => x"88",
          5815 => x"08",
          5816 => x"51",
          5817 => x"82",
          5818 => x"59",
          5819 => x"08",
          5820 => x"77",
          5821 => x"06",
          5822 => x"83",
          5823 => x"05",
          5824 => x"f7",
          5825 => x"39",
          5826 => x"a4",
          5827 => x"52",
          5828 => x"ef",
          5829 => x"a8",
          5830 => x"b5",
          5831 => x"38",
          5832 => x"06",
          5833 => x"83",
          5834 => x"18",
          5835 => x"54",
          5836 => x"f6",
          5837 => x"b5",
          5838 => x"0a",
          5839 => x"52",
          5840 => x"83",
          5841 => x"83",
          5842 => x"82",
          5843 => x"8a",
          5844 => x"f8",
          5845 => x"7c",
          5846 => x"59",
          5847 => x"81",
          5848 => x"38",
          5849 => x"08",
          5850 => x"73",
          5851 => x"38",
          5852 => x"52",
          5853 => x"a4",
          5854 => x"a8",
          5855 => x"b5",
          5856 => x"f2",
          5857 => x"82",
          5858 => x"39",
          5859 => x"e6",
          5860 => x"a8",
          5861 => x"de",
          5862 => x"78",
          5863 => x"3f",
          5864 => x"08",
          5865 => x"a8",
          5866 => x"80",
          5867 => x"b5",
          5868 => x"2e",
          5869 => x"b5",
          5870 => x"2e",
          5871 => x"53",
          5872 => x"51",
          5873 => x"82",
          5874 => x"c5",
          5875 => x"08",
          5876 => x"18",
          5877 => x"57",
          5878 => x"90",
          5879 => x"90",
          5880 => x"16",
          5881 => x"54",
          5882 => x"34",
          5883 => x"78",
          5884 => x"38",
          5885 => x"82",
          5886 => x"8a",
          5887 => x"f6",
          5888 => x"7e",
          5889 => x"5b",
          5890 => x"38",
          5891 => x"58",
          5892 => x"88",
          5893 => x"08",
          5894 => x"38",
          5895 => x"39",
          5896 => x"51",
          5897 => x"81",
          5898 => x"b5",
          5899 => x"82",
          5900 => x"b5",
          5901 => x"82",
          5902 => x"ff",
          5903 => x"38",
          5904 => x"82",
          5905 => x"26",
          5906 => x"79",
          5907 => x"08",
          5908 => x"73",
          5909 => x"b9",
          5910 => x"2e",
          5911 => x"80",
          5912 => x"1a",
          5913 => x"08",
          5914 => x"38",
          5915 => x"52",
          5916 => x"af",
          5917 => x"82",
          5918 => x"81",
          5919 => x"06",
          5920 => x"b5",
          5921 => x"82",
          5922 => x"09",
          5923 => x"72",
          5924 => x"70",
          5925 => x"b5",
          5926 => x"51",
          5927 => x"73",
          5928 => x"82",
          5929 => x"80",
          5930 => x"8c",
          5931 => x"81",
          5932 => x"38",
          5933 => x"08",
          5934 => x"73",
          5935 => x"75",
          5936 => x"77",
          5937 => x"56",
          5938 => x"76",
          5939 => x"82",
          5940 => x"26",
          5941 => x"75",
          5942 => x"f8",
          5943 => x"b5",
          5944 => x"2e",
          5945 => x"59",
          5946 => x"08",
          5947 => x"81",
          5948 => x"82",
          5949 => x"59",
          5950 => x"08",
          5951 => x"70",
          5952 => x"25",
          5953 => x"51",
          5954 => x"73",
          5955 => x"75",
          5956 => x"81",
          5957 => x"38",
          5958 => x"f5",
          5959 => x"75",
          5960 => x"f9",
          5961 => x"b5",
          5962 => x"b5",
          5963 => x"70",
          5964 => x"08",
          5965 => x"51",
          5966 => x"80",
          5967 => x"73",
          5968 => x"38",
          5969 => x"52",
          5970 => x"d0",
          5971 => x"a8",
          5972 => x"a5",
          5973 => x"18",
          5974 => x"08",
          5975 => x"18",
          5976 => x"74",
          5977 => x"38",
          5978 => x"18",
          5979 => x"33",
          5980 => x"73",
          5981 => x"97",
          5982 => x"74",
          5983 => x"38",
          5984 => x"55",
          5985 => x"b5",
          5986 => x"85",
          5987 => x"75",
          5988 => x"b5",
          5989 => x"3d",
          5990 => x"3d",
          5991 => x"52",
          5992 => x"3f",
          5993 => x"08",
          5994 => x"82",
          5995 => x"80",
          5996 => x"52",
          5997 => x"c1",
          5998 => x"a8",
          5999 => x"a8",
          6000 => x"0c",
          6001 => x"53",
          6002 => x"15",
          6003 => x"f2",
          6004 => x"56",
          6005 => x"16",
          6006 => x"22",
          6007 => x"27",
          6008 => x"54",
          6009 => x"76",
          6010 => x"33",
          6011 => x"3f",
          6012 => x"08",
          6013 => x"38",
          6014 => x"76",
          6015 => x"70",
          6016 => x"9f",
          6017 => x"56",
          6018 => x"b5",
          6019 => x"3d",
          6020 => x"3d",
          6021 => x"71",
          6022 => x"57",
          6023 => x"0a",
          6024 => x"38",
          6025 => x"53",
          6026 => x"38",
          6027 => x"0c",
          6028 => x"54",
          6029 => x"75",
          6030 => x"73",
          6031 => x"a8",
          6032 => x"73",
          6033 => x"85",
          6034 => x"0b",
          6035 => x"5a",
          6036 => x"27",
          6037 => x"a8",
          6038 => x"18",
          6039 => x"39",
          6040 => x"70",
          6041 => x"58",
          6042 => x"b2",
          6043 => x"76",
          6044 => x"3f",
          6045 => x"08",
          6046 => x"a8",
          6047 => x"bd",
          6048 => x"82",
          6049 => x"27",
          6050 => x"16",
          6051 => x"a8",
          6052 => x"38",
          6053 => x"39",
          6054 => x"55",
          6055 => x"52",
          6056 => x"d5",
          6057 => x"a8",
          6058 => x"0c",
          6059 => x"0c",
          6060 => x"53",
          6061 => x"80",
          6062 => x"85",
          6063 => x"94",
          6064 => x"2a",
          6065 => x"0c",
          6066 => x"06",
          6067 => x"9c",
          6068 => x"58",
          6069 => x"a8",
          6070 => x"0d",
          6071 => x"0d",
          6072 => x"90",
          6073 => x"05",
          6074 => x"f0",
          6075 => x"27",
          6076 => x"0b",
          6077 => x"98",
          6078 => x"84",
          6079 => x"2e",
          6080 => x"76",
          6081 => x"58",
          6082 => x"38",
          6083 => x"15",
          6084 => x"08",
          6085 => x"38",
          6086 => x"88",
          6087 => x"53",
          6088 => x"81",
          6089 => x"c0",
          6090 => x"22",
          6091 => x"89",
          6092 => x"72",
          6093 => x"74",
          6094 => x"f3",
          6095 => x"b5",
          6096 => x"82",
          6097 => x"82",
          6098 => x"27",
          6099 => x"81",
          6100 => x"a8",
          6101 => x"80",
          6102 => x"16",
          6103 => x"a8",
          6104 => x"ca",
          6105 => x"38",
          6106 => x"0c",
          6107 => x"dd",
          6108 => x"08",
          6109 => x"f9",
          6110 => x"b5",
          6111 => x"87",
          6112 => x"a8",
          6113 => x"80",
          6114 => x"55",
          6115 => x"08",
          6116 => x"38",
          6117 => x"b5",
          6118 => x"2e",
          6119 => x"b5",
          6120 => x"75",
          6121 => x"3f",
          6122 => x"08",
          6123 => x"94",
          6124 => x"52",
          6125 => x"c1",
          6126 => x"a8",
          6127 => x"0c",
          6128 => x"0c",
          6129 => x"05",
          6130 => x"80",
          6131 => x"b5",
          6132 => x"3d",
          6133 => x"3d",
          6134 => x"71",
          6135 => x"57",
          6136 => x"51",
          6137 => x"82",
          6138 => x"54",
          6139 => x"08",
          6140 => x"82",
          6141 => x"56",
          6142 => x"52",
          6143 => x"83",
          6144 => x"a8",
          6145 => x"b5",
          6146 => x"d2",
          6147 => x"a8",
          6148 => x"08",
          6149 => x"54",
          6150 => x"e5",
          6151 => x"06",
          6152 => x"58",
          6153 => x"08",
          6154 => x"38",
          6155 => x"75",
          6156 => x"80",
          6157 => x"81",
          6158 => x"7a",
          6159 => x"06",
          6160 => x"39",
          6161 => x"08",
          6162 => x"76",
          6163 => x"3f",
          6164 => x"08",
          6165 => x"a8",
          6166 => x"ff",
          6167 => x"84",
          6168 => x"06",
          6169 => x"54",
          6170 => x"a8",
          6171 => x"0d",
          6172 => x"0d",
          6173 => x"52",
          6174 => x"3f",
          6175 => x"08",
          6176 => x"06",
          6177 => x"51",
          6178 => x"83",
          6179 => x"06",
          6180 => x"14",
          6181 => x"3f",
          6182 => x"08",
          6183 => x"07",
          6184 => x"b5",
          6185 => x"3d",
          6186 => x"3d",
          6187 => x"70",
          6188 => x"06",
          6189 => x"53",
          6190 => x"ed",
          6191 => x"33",
          6192 => x"83",
          6193 => x"06",
          6194 => x"90",
          6195 => x"15",
          6196 => x"3f",
          6197 => x"04",
          6198 => x"7b",
          6199 => x"84",
          6200 => x"58",
          6201 => x"80",
          6202 => x"38",
          6203 => x"52",
          6204 => x"8f",
          6205 => x"a8",
          6206 => x"b5",
          6207 => x"f5",
          6208 => x"08",
          6209 => x"53",
          6210 => x"84",
          6211 => x"39",
          6212 => x"70",
          6213 => x"81",
          6214 => x"51",
          6215 => x"16",
          6216 => x"a8",
          6217 => x"81",
          6218 => x"38",
          6219 => x"ae",
          6220 => x"81",
          6221 => x"54",
          6222 => x"2e",
          6223 => x"8f",
          6224 => x"82",
          6225 => x"76",
          6226 => x"54",
          6227 => x"09",
          6228 => x"38",
          6229 => x"7a",
          6230 => x"80",
          6231 => x"fa",
          6232 => x"b5",
          6233 => x"82",
          6234 => x"89",
          6235 => x"08",
          6236 => x"86",
          6237 => x"98",
          6238 => x"82",
          6239 => x"8b",
          6240 => x"fb",
          6241 => x"70",
          6242 => x"81",
          6243 => x"fc",
          6244 => x"b5",
          6245 => x"82",
          6246 => x"b4",
          6247 => x"08",
          6248 => x"ec",
          6249 => x"b5",
          6250 => x"82",
          6251 => x"a0",
          6252 => x"82",
          6253 => x"52",
          6254 => x"51",
          6255 => x"8b",
          6256 => x"52",
          6257 => x"51",
          6258 => x"81",
          6259 => x"34",
          6260 => x"a8",
          6261 => x"0d",
          6262 => x"0d",
          6263 => x"98",
          6264 => x"70",
          6265 => x"ec",
          6266 => x"b5",
          6267 => x"38",
          6268 => x"53",
          6269 => x"81",
          6270 => x"34",
          6271 => x"04",
          6272 => x"78",
          6273 => x"80",
          6274 => x"34",
          6275 => x"80",
          6276 => x"38",
          6277 => x"18",
          6278 => x"9c",
          6279 => x"70",
          6280 => x"56",
          6281 => x"a0",
          6282 => x"71",
          6283 => x"81",
          6284 => x"81",
          6285 => x"89",
          6286 => x"06",
          6287 => x"73",
          6288 => x"55",
          6289 => x"55",
          6290 => x"81",
          6291 => x"81",
          6292 => x"74",
          6293 => x"75",
          6294 => x"52",
          6295 => x"13",
          6296 => x"08",
          6297 => x"33",
          6298 => x"9c",
          6299 => x"11",
          6300 => x"8a",
          6301 => x"a8",
          6302 => x"96",
          6303 => x"e7",
          6304 => x"a8",
          6305 => x"23",
          6306 => x"e7",
          6307 => x"b5",
          6308 => x"17",
          6309 => x"0d",
          6310 => x"0d",
          6311 => x"5e",
          6312 => x"70",
          6313 => x"55",
          6314 => x"83",
          6315 => x"73",
          6316 => x"91",
          6317 => x"2e",
          6318 => x"1d",
          6319 => x"0c",
          6320 => x"15",
          6321 => x"70",
          6322 => x"56",
          6323 => x"09",
          6324 => x"38",
          6325 => x"80",
          6326 => x"30",
          6327 => x"78",
          6328 => x"54",
          6329 => x"73",
          6330 => x"60",
          6331 => x"54",
          6332 => x"96",
          6333 => x"0b",
          6334 => x"80",
          6335 => x"f6",
          6336 => x"b5",
          6337 => x"85",
          6338 => x"3d",
          6339 => x"5c",
          6340 => x"53",
          6341 => x"51",
          6342 => x"80",
          6343 => x"88",
          6344 => x"5c",
          6345 => x"09",
          6346 => x"d4",
          6347 => x"70",
          6348 => x"71",
          6349 => x"30",
          6350 => x"73",
          6351 => x"51",
          6352 => x"57",
          6353 => x"38",
          6354 => x"75",
          6355 => x"17",
          6356 => x"75",
          6357 => x"30",
          6358 => x"51",
          6359 => x"80",
          6360 => x"38",
          6361 => x"87",
          6362 => x"26",
          6363 => x"77",
          6364 => x"a4",
          6365 => x"27",
          6366 => x"a0",
          6367 => x"39",
          6368 => x"33",
          6369 => x"57",
          6370 => x"27",
          6371 => x"75",
          6372 => x"30",
          6373 => x"32",
          6374 => x"80",
          6375 => x"25",
          6376 => x"56",
          6377 => x"80",
          6378 => x"84",
          6379 => x"58",
          6380 => x"70",
          6381 => x"55",
          6382 => x"09",
          6383 => x"38",
          6384 => x"80",
          6385 => x"30",
          6386 => x"77",
          6387 => x"54",
          6388 => x"81",
          6389 => x"ae",
          6390 => x"06",
          6391 => x"54",
          6392 => x"74",
          6393 => x"80",
          6394 => x"7b",
          6395 => x"30",
          6396 => x"70",
          6397 => x"25",
          6398 => x"07",
          6399 => x"51",
          6400 => x"a7",
          6401 => x"8b",
          6402 => x"39",
          6403 => x"54",
          6404 => x"8c",
          6405 => x"ff",
          6406 => x"f0",
          6407 => x"54",
          6408 => x"e1",
          6409 => x"a8",
          6410 => x"b2",
          6411 => x"70",
          6412 => x"71",
          6413 => x"54",
          6414 => x"82",
          6415 => x"80",
          6416 => x"38",
          6417 => x"76",
          6418 => x"df",
          6419 => x"54",
          6420 => x"81",
          6421 => x"55",
          6422 => x"34",
          6423 => x"52",
          6424 => x"51",
          6425 => x"82",
          6426 => x"bf",
          6427 => x"16",
          6428 => x"26",
          6429 => x"16",
          6430 => x"06",
          6431 => x"17",
          6432 => x"34",
          6433 => x"fd",
          6434 => x"19",
          6435 => x"80",
          6436 => x"79",
          6437 => x"81",
          6438 => x"81",
          6439 => x"85",
          6440 => x"54",
          6441 => x"8f",
          6442 => x"86",
          6443 => x"39",
          6444 => x"f3",
          6445 => x"73",
          6446 => x"80",
          6447 => x"52",
          6448 => x"ce",
          6449 => x"a8",
          6450 => x"b5",
          6451 => x"d7",
          6452 => x"08",
          6453 => x"e6",
          6454 => x"b5",
          6455 => x"82",
          6456 => x"80",
          6457 => x"1b",
          6458 => x"55",
          6459 => x"2e",
          6460 => x"8b",
          6461 => x"06",
          6462 => x"1c",
          6463 => x"33",
          6464 => x"70",
          6465 => x"55",
          6466 => x"38",
          6467 => x"52",
          6468 => x"9f",
          6469 => x"a8",
          6470 => x"8b",
          6471 => x"7a",
          6472 => x"3f",
          6473 => x"75",
          6474 => x"57",
          6475 => x"2e",
          6476 => x"84",
          6477 => x"06",
          6478 => x"75",
          6479 => x"81",
          6480 => x"2a",
          6481 => x"73",
          6482 => x"38",
          6483 => x"54",
          6484 => x"fb",
          6485 => x"80",
          6486 => x"34",
          6487 => x"c1",
          6488 => x"06",
          6489 => x"38",
          6490 => x"39",
          6491 => x"70",
          6492 => x"54",
          6493 => x"86",
          6494 => x"84",
          6495 => x"06",
          6496 => x"73",
          6497 => x"38",
          6498 => x"83",
          6499 => x"b4",
          6500 => x"51",
          6501 => x"82",
          6502 => x"88",
          6503 => x"ea",
          6504 => x"b5",
          6505 => x"3d",
          6506 => x"3d",
          6507 => x"ff",
          6508 => x"71",
          6509 => x"5c",
          6510 => x"80",
          6511 => x"38",
          6512 => x"05",
          6513 => x"a0",
          6514 => x"71",
          6515 => x"38",
          6516 => x"71",
          6517 => x"81",
          6518 => x"38",
          6519 => x"11",
          6520 => x"06",
          6521 => x"70",
          6522 => x"38",
          6523 => x"81",
          6524 => x"05",
          6525 => x"76",
          6526 => x"38",
          6527 => x"ae",
          6528 => x"77",
          6529 => x"57",
          6530 => x"05",
          6531 => x"70",
          6532 => x"33",
          6533 => x"53",
          6534 => x"99",
          6535 => x"e0",
          6536 => x"ff",
          6537 => x"ff",
          6538 => x"70",
          6539 => x"38",
          6540 => x"81",
          6541 => x"51",
          6542 => x"9f",
          6543 => x"72",
          6544 => x"81",
          6545 => x"70",
          6546 => x"72",
          6547 => x"32",
          6548 => x"72",
          6549 => x"73",
          6550 => x"53",
          6551 => x"70",
          6552 => x"38",
          6553 => x"19",
          6554 => x"75",
          6555 => x"38",
          6556 => x"83",
          6557 => x"74",
          6558 => x"59",
          6559 => x"39",
          6560 => x"33",
          6561 => x"b5",
          6562 => x"3d",
          6563 => x"3d",
          6564 => x"80",
          6565 => x"34",
          6566 => x"17",
          6567 => x"75",
          6568 => x"3f",
          6569 => x"b5",
          6570 => x"80",
          6571 => x"16",
          6572 => x"3f",
          6573 => x"08",
          6574 => x"06",
          6575 => x"73",
          6576 => x"2e",
          6577 => x"80",
          6578 => x"0b",
          6579 => x"56",
          6580 => x"e9",
          6581 => x"06",
          6582 => x"57",
          6583 => x"32",
          6584 => x"80",
          6585 => x"51",
          6586 => x"8a",
          6587 => x"e8",
          6588 => x"06",
          6589 => x"53",
          6590 => x"52",
          6591 => x"51",
          6592 => x"82",
          6593 => x"55",
          6594 => x"08",
          6595 => x"38",
          6596 => x"ae",
          6597 => x"86",
          6598 => x"97",
          6599 => x"a8",
          6600 => x"b5",
          6601 => x"2e",
          6602 => x"55",
          6603 => x"a8",
          6604 => x"0d",
          6605 => x"0d",
          6606 => x"05",
          6607 => x"33",
          6608 => x"75",
          6609 => x"fc",
          6610 => x"b5",
          6611 => x"8b",
          6612 => x"82",
          6613 => x"24",
          6614 => x"82",
          6615 => x"84",
          6616 => x"e0",
          6617 => x"55",
          6618 => x"73",
          6619 => x"e6",
          6620 => x"0c",
          6621 => x"06",
          6622 => x"57",
          6623 => x"ae",
          6624 => x"33",
          6625 => x"3f",
          6626 => x"08",
          6627 => x"70",
          6628 => x"55",
          6629 => x"76",
          6630 => x"b8",
          6631 => x"2a",
          6632 => x"51",
          6633 => x"72",
          6634 => x"86",
          6635 => x"74",
          6636 => x"15",
          6637 => x"81",
          6638 => x"d7",
          6639 => x"b5",
          6640 => x"ff",
          6641 => x"06",
          6642 => x"56",
          6643 => x"38",
          6644 => x"8f",
          6645 => x"2a",
          6646 => x"51",
          6647 => x"72",
          6648 => x"80",
          6649 => x"52",
          6650 => x"3f",
          6651 => x"08",
          6652 => x"57",
          6653 => x"09",
          6654 => x"e2",
          6655 => x"74",
          6656 => x"56",
          6657 => x"33",
          6658 => x"72",
          6659 => x"38",
          6660 => x"51",
          6661 => x"82",
          6662 => x"57",
          6663 => x"84",
          6664 => x"ff",
          6665 => x"56",
          6666 => x"25",
          6667 => x"0b",
          6668 => x"56",
          6669 => x"05",
          6670 => x"83",
          6671 => x"2e",
          6672 => x"52",
          6673 => x"c6",
          6674 => x"a8",
          6675 => x"06",
          6676 => x"27",
          6677 => x"16",
          6678 => x"27",
          6679 => x"56",
          6680 => x"84",
          6681 => x"56",
          6682 => x"84",
          6683 => x"14",
          6684 => x"3f",
          6685 => x"08",
          6686 => x"06",
          6687 => x"80",
          6688 => x"06",
          6689 => x"80",
          6690 => x"db",
          6691 => x"b5",
          6692 => x"ff",
          6693 => x"77",
          6694 => x"d8",
          6695 => x"de",
          6696 => x"a8",
          6697 => x"9c",
          6698 => x"c4",
          6699 => x"15",
          6700 => x"14",
          6701 => x"70",
          6702 => x"51",
          6703 => x"56",
          6704 => x"84",
          6705 => x"81",
          6706 => x"71",
          6707 => x"16",
          6708 => x"53",
          6709 => x"23",
          6710 => x"8b",
          6711 => x"73",
          6712 => x"80",
          6713 => x"8d",
          6714 => x"39",
          6715 => x"51",
          6716 => x"82",
          6717 => x"53",
          6718 => x"08",
          6719 => x"72",
          6720 => x"8d",
          6721 => x"ce",
          6722 => x"14",
          6723 => x"3f",
          6724 => x"08",
          6725 => x"06",
          6726 => x"38",
          6727 => x"51",
          6728 => x"82",
          6729 => x"55",
          6730 => x"51",
          6731 => x"82",
          6732 => x"83",
          6733 => x"53",
          6734 => x"80",
          6735 => x"38",
          6736 => x"78",
          6737 => x"2a",
          6738 => x"78",
          6739 => x"86",
          6740 => x"22",
          6741 => x"31",
          6742 => x"ca",
          6743 => x"a8",
          6744 => x"b5",
          6745 => x"2e",
          6746 => x"82",
          6747 => x"80",
          6748 => x"f5",
          6749 => x"83",
          6750 => x"ff",
          6751 => x"38",
          6752 => x"9f",
          6753 => x"38",
          6754 => x"39",
          6755 => x"80",
          6756 => x"38",
          6757 => x"98",
          6758 => x"a0",
          6759 => x"1c",
          6760 => x"0c",
          6761 => x"17",
          6762 => x"76",
          6763 => x"81",
          6764 => x"80",
          6765 => x"d9",
          6766 => x"b5",
          6767 => x"ff",
          6768 => x"8d",
          6769 => x"8e",
          6770 => x"8a",
          6771 => x"14",
          6772 => x"3f",
          6773 => x"08",
          6774 => x"74",
          6775 => x"a2",
          6776 => x"79",
          6777 => x"ee",
          6778 => x"a8",
          6779 => x"15",
          6780 => x"2e",
          6781 => x"10",
          6782 => x"2a",
          6783 => x"05",
          6784 => x"ff",
          6785 => x"53",
          6786 => x"9c",
          6787 => x"81",
          6788 => x"0b",
          6789 => x"ff",
          6790 => x"0c",
          6791 => x"84",
          6792 => x"83",
          6793 => x"06",
          6794 => x"80",
          6795 => x"d8",
          6796 => x"b5",
          6797 => x"ff",
          6798 => x"72",
          6799 => x"81",
          6800 => x"38",
          6801 => x"73",
          6802 => x"3f",
          6803 => x"08",
          6804 => x"82",
          6805 => x"84",
          6806 => x"b2",
          6807 => x"87",
          6808 => x"a8",
          6809 => x"ff",
          6810 => x"82",
          6811 => x"09",
          6812 => x"c8",
          6813 => x"51",
          6814 => x"82",
          6815 => x"84",
          6816 => x"d2",
          6817 => x"06",
          6818 => x"98",
          6819 => x"ee",
          6820 => x"a8",
          6821 => x"85",
          6822 => x"09",
          6823 => x"38",
          6824 => x"51",
          6825 => x"82",
          6826 => x"90",
          6827 => x"a0",
          6828 => x"ca",
          6829 => x"a8",
          6830 => x"0c",
          6831 => x"82",
          6832 => x"81",
          6833 => x"82",
          6834 => x"72",
          6835 => x"80",
          6836 => x"0c",
          6837 => x"82",
          6838 => x"90",
          6839 => x"fb",
          6840 => x"54",
          6841 => x"80",
          6842 => x"73",
          6843 => x"80",
          6844 => x"72",
          6845 => x"80",
          6846 => x"86",
          6847 => x"15",
          6848 => x"71",
          6849 => x"81",
          6850 => x"81",
          6851 => x"d0",
          6852 => x"b5",
          6853 => x"06",
          6854 => x"38",
          6855 => x"54",
          6856 => x"80",
          6857 => x"71",
          6858 => x"82",
          6859 => x"87",
          6860 => x"fa",
          6861 => x"ab",
          6862 => x"58",
          6863 => x"05",
          6864 => x"e6",
          6865 => x"80",
          6866 => x"a8",
          6867 => x"38",
          6868 => x"08",
          6869 => x"cc",
          6870 => x"08",
          6871 => x"80",
          6872 => x"80",
          6873 => x"54",
          6874 => x"84",
          6875 => x"34",
          6876 => x"75",
          6877 => x"2e",
          6878 => x"53",
          6879 => x"53",
          6880 => x"f7",
          6881 => x"b5",
          6882 => x"73",
          6883 => x"0c",
          6884 => x"04",
          6885 => x"67",
          6886 => x"80",
          6887 => x"59",
          6888 => x"78",
          6889 => x"c8",
          6890 => x"06",
          6891 => x"3d",
          6892 => x"99",
          6893 => x"52",
          6894 => x"3f",
          6895 => x"08",
          6896 => x"a8",
          6897 => x"38",
          6898 => x"52",
          6899 => x"52",
          6900 => x"3f",
          6901 => x"08",
          6902 => x"a8",
          6903 => x"02",
          6904 => x"33",
          6905 => x"55",
          6906 => x"25",
          6907 => x"55",
          6908 => x"54",
          6909 => x"81",
          6910 => x"80",
          6911 => x"74",
          6912 => x"81",
          6913 => x"75",
          6914 => x"3f",
          6915 => x"08",
          6916 => x"02",
          6917 => x"91",
          6918 => x"81",
          6919 => x"82",
          6920 => x"06",
          6921 => x"80",
          6922 => x"88",
          6923 => x"39",
          6924 => x"58",
          6925 => x"38",
          6926 => x"70",
          6927 => x"54",
          6928 => x"81",
          6929 => x"52",
          6930 => x"a5",
          6931 => x"a8",
          6932 => x"88",
          6933 => x"62",
          6934 => x"d4",
          6935 => x"54",
          6936 => x"15",
          6937 => x"62",
          6938 => x"e8",
          6939 => x"52",
          6940 => x"51",
          6941 => x"7a",
          6942 => x"83",
          6943 => x"80",
          6944 => x"38",
          6945 => x"08",
          6946 => x"53",
          6947 => x"3d",
          6948 => x"dd",
          6949 => x"b5",
          6950 => x"82",
          6951 => x"82",
          6952 => x"39",
          6953 => x"38",
          6954 => x"33",
          6955 => x"70",
          6956 => x"55",
          6957 => x"2e",
          6958 => x"55",
          6959 => x"77",
          6960 => x"81",
          6961 => x"73",
          6962 => x"38",
          6963 => x"54",
          6964 => x"a0",
          6965 => x"82",
          6966 => x"52",
          6967 => x"a3",
          6968 => x"a8",
          6969 => x"18",
          6970 => x"55",
          6971 => x"a8",
          6972 => x"38",
          6973 => x"70",
          6974 => x"54",
          6975 => x"86",
          6976 => x"c0",
          6977 => x"b0",
          6978 => x"1b",
          6979 => x"1b",
          6980 => x"70",
          6981 => x"d9",
          6982 => x"a8",
          6983 => x"a8",
          6984 => x"0c",
          6985 => x"52",
          6986 => x"3f",
          6987 => x"08",
          6988 => x"08",
          6989 => x"77",
          6990 => x"86",
          6991 => x"1a",
          6992 => x"1a",
          6993 => x"91",
          6994 => x"0b",
          6995 => x"80",
          6996 => x"0c",
          6997 => x"70",
          6998 => x"54",
          6999 => x"81",
          7000 => x"b5",
          7001 => x"2e",
          7002 => x"82",
          7003 => x"94",
          7004 => x"17",
          7005 => x"2b",
          7006 => x"57",
          7007 => x"52",
          7008 => x"9f",
          7009 => x"a8",
          7010 => x"b5",
          7011 => x"26",
          7012 => x"55",
          7013 => x"08",
          7014 => x"81",
          7015 => x"79",
          7016 => x"31",
          7017 => x"70",
          7018 => x"25",
          7019 => x"76",
          7020 => x"81",
          7021 => x"55",
          7022 => x"38",
          7023 => x"0c",
          7024 => x"75",
          7025 => x"54",
          7026 => x"a2",
          7027 => x"7a",
          7028 => x"3f",
          7029 => x"08",
          7030 => x"55",
          7031 => x"89",
          7032 => x"a8",
          7033 => x"1a",
          7034 => x"80",
          7035 => x"54",
          7036 => x"a8",
          7037 => x"0d",
          7038 => x"0d",
          7039 => x"64",
          7040 => x"59",
          7041 => x"90",
          7042 => x"52",
          7043 => x"cf",
          7044 => x"a8",
          7045 => x"b5",
          7046 => x"38",
          7047 => x"55",
          7048 => x"86",
          7049 => x"82",
          7050 => x"19",
          7051 => x"55",
          7052 => x"80",
          7053 => x"38",
          7054 => x"0b",
          7055 => x"82",
          7056 => x"39",
          7057 => x"1a",
          7058 => x"82",
          7059 => x"19",
          7060 => x"08",
          7061 => x"7c",
          7062 => x"74",
          7063 => x"2e",
          7064 => x"94",
          7065 => x"83",
          7066 => x"56",
          7067 => x"38",
          7068 => x"22",
          7069 => x"89",
          7070 => x"55",
          7071 => x"75",
          7072 => x"19",
          7073 => x"39",
          7074 => x"52",
          7075 => x"93",
          7076 => x"a8",
          7077 => x"75",
          7078 => x"38",
          7079 => x"ff",
          7080 => x"98",
          7081 => x"19",
          7082 => x"51",
          7083 => x"82",
          7084 => x"80",
          7085 => x"38",
          7086 => x"08",
          7087 => x"2a",
          7088 => x"80",
          7089 => x"38",
          7090 => x"8a",
          7091 => x"5c",
          7092 => x"27",
          7093 => x"7a",
          7094 => x"54",
          7095 => x"52",
          7096 => x"51",
          7097 => x"82",
          7098 => x"fe",
          7099 => x"83",
          7100 => x"56",
          7101 => x"9f",
          7102 => x"08",
          7103 => x"74",
          7104 => x"38",
          7105 => x"b4",
          7106 => x"16",
          7107 => x"89",
          7108 => x"51",
          7109 => x"77",
          7110 => x"b9",
          7111 => x"1a",
          7112 => x"08",
          7113 => x"84",
          7114 => x"57",
          7115 => x"27",
          7116 => x"56",
          7117 => x"52",
          7118 => x"c7",
          7119 => x"a8",
          7120 => x"38",
          7121 => x"19",
          7122 => x"06",
          7123 => x"52",
          7124 => x"a2",
          7125 => x"31",
          7126 => x"7f",
          7127 => x"94",
          7128 => x"94",
          7129 => x"5c",
          7130 => x"80",
          7131 => x"b5",
          7132 => x"3d",
          7133 => x"3d",
          7134 => x"65",
          7135 => x"5d",
          7136 => x"0c",
          7137 => x"05",
          7138 => x"f6",
          7139 => x"b5",
          7140 => x"82",
          7141 => x"8a",
          7142 => x"33",
          7143 => x"2e",
          7144 => x"56",
          7145 => x"90",
          7146 => x"81",
          7147 => x"06",
          7148 => x"87",
          7149 => x"2e",
          7150 => x"95",
          7151 => x"91",
          7152 => x"56",
          7153 => x"81",
          7154 => x"34",
          7155 => x"8e",
          7156 => x"08",
          7157 => x"56",
          7158 => x"84",
          7159 => x"5c",
          7160 => x"82",
          7161 => x"18",
          7162 => x"ff",
          7163 => x"74",
          7164 => x"7e",
          7165 => x"ff",
          7166 => x"2a",
          7167 => x"7a",
          7168 => x"8c",
          7169 => x"08",
          7170 => x"38",
          7171 => x"39",
          7172 => x"52",
          7173 => x"e7",
          7174 => x"a8",
          7175 => x"b5",
          7176 => x"2e",
          7177 => x"74",
          7178 => x"91",
          7179 => x"2e",
          7180 => x"74",
          7181 => x"88",
          7182 => x"38",
          7183 => x"0c",
          7184 => x"15",
          7185 => x"08",
          7186 => x"06",
          7187 => x"51",
          7188 => x"82",
          7189 => x"fe",
          7190 => x"18",
          7191 => x"51",
          7192 => x"82",
          7193 => x"80",
          7194 => x"38",
          7195 => x"08",
          7196 => x"2a",
          7197 => x"80",
          7198 => x"38",
          7199 => x"8a",
          7200 => x"5b",
          7201 => x"27",
          7202 => x"7b",
          7203 => x"54",
          7204 => x"52",
          7205 => x"51",
          7206 => x"82",
          7207 => x"fe",
          7208 => x"b0",
          7209 => x"31",
          7210 => x"79",
          7211 => x"84",
          7212 => x"16",
          7213 => x"89",
          7214 => x"52",
          7215 => x"cc",
          7216 => x"55",
          7217 => x"16",
          7218 => x"2b",
          7219 => x"39",
          7220 => x"94",
          7221 => x"93",
          7222 => x"cd",
          7223 => x"b5",
          7224 => x"e3",
          7225 => x"b0",
          7226 => x"76",
          7227 => x"94",
          7228 => x"ff",
          7229 => x"71",
          7230 => x"7b",
          7231 => x"38",
          7232 => x"18",
          7233 => x"51",
          7234 => x"82",
          7235 => x"fd",
          7236 => x"53",
          7237 => x"18",
          7238 => x"06",
          7239 => x"51",
          7240 => x"7e",
          7241 => x"83",
          7242 => x"76",
          7243 => x"17",
          7244 => x"1e",
          7245 => x"18",
          7246 => x"0c",
          7247 => x"58",
          7248 => x"74",
          7249 => x"38",
          7250 => x"8c",
          7251 => x"90",
          7252 => x"33",
          7253 => x"55",
          7254 => x"34",
          7255 => x"82",
          7256 => x"90",
          7257 => x"f8",
          7258 => x"8b",
          7259 => x"53",
          7260 => x"f2",
          7261 => x"b5",
          7262 => x"82",
          7263 => x"80",
          7264 => x"16",
          7265 => x"2a",
          7266 => x"51",
          7267 => x"80",
          7268 => x"38",
          7269 => x"52",
          7270 => x"e7",
          7271 => x"a8",
          7272 => x"b5",
          7273 => x"d4",
          7274 => x"08",
          7275 => x"a0",
          7276 => x"73",
          7277 => x"88",
          7278 => x"74",
          7279 => x"51",
          7280 => x"8c",
          7281 => x"9c",
          7282 => x"fb",
          7283 => x"b2",
          7284 => x"15",
          7285 => x"3f",
          7286 => x"15",
          7287 => x"3f",
          7288 => x"0b",
          7289 => x"78",
          7290 => x"3f",
          7291 => x"08",
          7292 => x"81",
          7293 => x"57",
          7294 => x"34",
          7295 => x"a8",
          7296 => x"0d",
          7297 => x"0d",
          7298 => x"54",
          7299 => x"82",
          7300 => x"53",
          7301 => x"08",
          7302 => x"3d",
          7303 => x"73",
          7304 => x"3f",
          7305 => x"08",
          7306 => x"a8",
          7307 => x"82",
          7308 => x"74",
          7309 => x"b5",
          7310 => x"3d",
          7311 => x"3d",
          7312 => x"51",
          7313 => x"8b",
          7314 => x"82",
          7315 => x"24",
          7316 => x"b5",
          7317 => x"cc",
          7318 => x"52",
          7319 => x"a8",
          7320 => x"0d",
          7321 => x"0d",
          7322 => x"3d",
          7323 => x"94",
          7324 => x"c1",
          7325 => x"a8",
          7326 => x"b5",
          7327 => x"e0",
          7328 => x"63",
          7329 => x"d4",
          7330 => x"8d",
          7331 => x"a8",
          7332 => x"b5",
          7333 => x"38",
          7334 => x"05",
          7335 => x"2b",
          7336 => x"80",
          7337 => x"76",
          7338 => x"0c",
          7339 => x"02",
          7340 => x"70",
          7341 => x"81",
          7342 => x"56",
          7343 => x"9e",
          7344 => x"53",
          7345 => x"db",
          7346 => x"b5",
          7347 => x"15",
          7348 => x"82",
          7349 => x"84",
          7350 => x"06",
          7351 => x"55",
          7352 => x"a8",
          7353 => x"0d",
          7354 => x"0d",
          7355 => x"5b",
          7356 => x"80",
          7357 => x"ff",
          7358 => x"9f",
          7359 => x"b5",
          7360 => x"a8",
          7361 => x"b5",
          7362 => x"fc",
          7363 => x"7a",
          7364 => x"08",
          7365 => x"64",
          7366 => x"2e",
          7367 => x"a0",
          7368 => x"70",
          7369 => x"ea",
          7370 => x"a8",
          7371 => x"b5",
          7372 => x"d4",
          7373 => x"7b",
          7374 => x"3f",
          7375 => x"08",
          7376 => x"a8",
          7377 => x"38",
          7378 => x"51",
          7379 => x"82",
          7380 => x"45",
          7381 => x"51",
          7382 => x"82",
          7383 => x"57",
          7384 => x"08",
          7385 => x"80",
          7386 => x"da",
          7387 => x"b5",
          7388 => x"82",
          7389 => x"a4",
          7390 => x"7b",
          7391 => x"3f",
          7392 => x"a8",
          7393 => x"38",
          7394 => x"51",
          7395 => x"82",
          7396 => x"57",
          7397 => x"08",
          7398 => x"38",
          7399 => x"09",
          7400 => x"38",
          7401 => x"e0",
          7402 => x"dc",
          7403 => x"ff",
          7404 => x"74",
          7405 => x"3f",
          7406 => x"78",
          7407 => x"33",
          7408 => x"56",
          7409 => x"91",
          7410 => x"05",
          7411 => x"81",
          7412 => x"56",
          7413 => x"f5",
          7414 => x"54",
          7415 => x"81",
          7416 => x"80",
          7417 => x"78",
          7418 => x"55",
          7419 => x"11",
          7420 => x"18",
          7421 => x"58",
          7422 => x"34",
          7423 => x"ff",
          7424 => x"55",
          7425 => x"34",
          7426 => x"77",
          7427 => x"81",
          7428 => x"ff",
          7429 => x"55",
          7430 => x"34",
          7431 => x"cc",
          7432 => x"84",
          7433 => x"e0",
          7434 => x"70",
          7435 => x"56",
          7436 => x"76",
          7437 => x"81",
          7438 => x"70",
          7439 => x"56",
          7440 => x"82",
          7441 => x"78",
          7442 => x"80",
          7443 => x"27",
          7444 => x"19",
          7445 => x"7a",
          7446 => x"5c",
          7447 => x"55",
          7448 => x"7a",
          7449 => x"5c",
          7450 => x"2e",
          7451 => x"85",
          7452 => x"94",
          7453 => x"81",
          7454 => x"73",
          7455 => x"81",
          7456 => x"7a",
          7457 => x"38",
          7458 => x"76",
          7459 => x"0c",
          7460 => x"04",
          7461 => x"7b",
          7462 => x"fc",
          7463 => x"53",
          7464 => x"bb",
          7465 => x"a8",
          7466 => x"b5",
          7467 => x"fa",
          7468 => x"33",
          7469 => x"f2",
          7470 => x"08",
          7471 => x"27",
          7472 => x"15",
          7473 => x"2a",
          7474 => x"51",
          7475 => x"83",
          7476 => x"94",
          7477 => x"80",
          7478 => x"0c",
          7479 => x"2e",
          7480 => x"79",
          7481 => x"70",
          7482 => x"51",
          7483 => x"2e",
          7484 => x"52",
          7485 => x"fe",
          7486 => x"82",
          7487 => x"ff",
          7488 => x"70",
          7489 => x"fe",
          7490 => x"82",
          7491 => x"73",
          7492 => x"76",
          7493 => x"06",
          7494 => x"0c",
          7495 => x"98",
          7496 => x"58",
          7497 => x"39",
          7498 => x"54",
          7499 => x"73",
          7500 => x"cd",
          7501 => x"b5",
          7502 => x"82",
          7503 => x"81",
          7504 => x"38",
          7505 => x"08",
          7506 => x"9b",
          7507 => x"a8",
          7508 => x"0c",
          7509 => x"0c",
          7510 => x"81",
          7511 => x"76",
          7512 => x"38",
          7513 => x"94",
          7514 => x"94",
          7515 => x"16",
          7516 => x"2a",
          7517 => x"51",
          7518 => x"72",
          7519 => x"38",
          7520 => x"51",
          7521 => x"82",
          7522 => x"54",
          7523 => x"08",
          7524 => x"b5",
          7525 => x"a7",
          7526 => x"74",
          7527 => x"3f",
          7528 => x"08",
          7529 => x"2e",
          7530 => x"74",
          7531 => x"79",
          7532 => x"14",
          7533 => x"38",
          7534 => x"0c",
          7535 => x"94",
          7536 => x"94",
          7537 => x"83",
          7538 => x"72",
          7539 => x"38",
          7540 => x"51",
          7541 => x"82",
          7542 => x"94",
          7543 => x"91",
          7544 => x"53",
          7545 => x"81",
          7546 => x"34",
          7547 => x"39",
          7548 => x"82",
          7549 => x"05",
          7550 => x"08",
          7551 => x"08",
          7552 => x"38",
          7553 => x"0c",
          7554 => x"80",
          7555 => x"72",
          7556 => x"73",
          7557 => x"53",
          7558 => x"8c",
          7559 => x"16",
          7560 => x"38",
          7561 => x"0c",
          7562 => x"82",
          7563 => x"8b",
          7564 => x"f9",
          7565 => x"56",
          7566 => x"80",
          7567 => x"38",
          7568 => x"3d",
          7569 => x"8a",
          7570 => x"51",
          7571 => x"82",
          7572 => x"55",
          7573 => x"08",
          7574 => x"77",
          7575 => x"52",
          7576 => x"b5",
          7577 => x"a8",
          7578 => x"b5",
          7579 => x"c3",
          7580 => x"33",
          7581 => x"55",
          7582 => x"24",
          7583 => x"16",
          7584 => x"2a",
          7585 => x"51",
          7586 => x"80",
          7587 => x"9c",
          7588 => x"77",
          7589 => x"3f",
          7590 => x"08",
          7591 => x"77",
          7592 => x"22",
          7593 => x"74",
          7594 => x"ce",
          7595 => x"b5",
          7596 => x"74",
          7597 => x"81",
          7598 => x"85",
          7599 => x"74",
          7600 => x"38",
          7601 => x"74",
          7602 => x"b5",
          7603 => x"3d",
          7604 => x"3d",
          7605 => x"3d",
          7606 => x"70",
          7607 => x"ff",
          7608 => x"a8",
          7609 => x"82",
          7610 => x"73",
          7611 => x"0d",
          7612 => x"0d",
          7613 => x"3d",
          7614 => x"71",
          7615 => x"e7",
          7616 => x"b5",
          7617 => x"82",
          7618 => x"80",
          7619 => x"93",
          7620 => x"a8",
          7621 => x"51",
          7622 => x"82",
          7623 => x"53",
          7624 => x"82",
          7625 => x"52",
          7626 => x"ac",
          7627 => x"a8",
          7628 => x"b5",
          7629 => x"2e",
          7630 => x"85",
          7631 => x"87",
          7632 => x"a8",
          7633 => x"74",
          7634 => x"d5",
          7635 => x"52",
          7636 => x"89",
          7637 => x"a8",
          7638 => x"70",
          7639 => x"07",
          7640 => x"82",
          7641 => x"06",
          7642 => x"54",
          7643 => x"a8",
          7644 => x"0d",
          7645 => x"0d",
          7646 => x"53",
          7647 => x"53",
          7648 => x"56",
          7649 => x"82",
          7650 => x"55",
          7651 => x"08",
          7652 => x"52",
          7653 => x"81",
          7654 => x"a8",
          7655 => x"b5",
          7656 => x"38",
          7657 => x"05",
          7658 => x"2b",
          7659 => x"80",
          7660 => x"86",
          7661 => x"76",
          7662 => x"38",
          7663 => x"51",
          7664 => x"74",
          7665 => x"0c",
          7666 => x"04",
          7667 => x"63",
          7668 => x"80",
          7669 => x"ec",
          7670 => x"3d",
          7671 => x"3f",
          7672 => x"08",
          7673 => x"a8",
          7674 => x"38",
          7675 => x"73",
          7676 => x"08",
          7677 => x"13",
          7678 => x"58",
          7679 => x"26",
          7680 => x"7c",
          7681 => x"39",
          7682 => x"cc",
          7683 => x"81",
          7684 => x"b5",
          7685 => x"33",
          7686 => x"81",
          7687 => x"06",
          7688 => x"75",
          7689 => x"52",
          7690 => x"05",
          7691 => x"3f",
          7692 => x"08",
          7693 => x"38",
          7694 => x"08",
          7695 => x"38",
          7696 => x"08",
          7697 => x"b5",
          7698 => x"80",
          7699 => x"81",
          7700 => x"59",
          7701 => x"14",
          7702 => x"ca",
          7703 => x"39",
          7704 => x"82",
          7705 => x"57",
          7706 => x"38",
          7707 => x"18",
          7708 => x"ff",
          7709 => x"82",
          7710 => x"5b",
          7711 => x"08",
          7712 => x"7c",
          7713 => x"12",
          7714 => x"52",
          7715 => x"82",
          7716 => x"06",
          7717 => x"14",
          7718 => x"cb",
          7719 => x"a8",
          7720 => x"ff",
          7721 => x"70",
          7722 => x"82",
          7723 => x"51",
          7724 => x"b4",
          7725 => x"bb",
          7726 => x"b5",
          7727 => x"0a",
          7728 => x"70",
          7729 => x"84",
          7730 => x"51",
          7731 => x"ff",
          7732 => x"56",
          7733 => x"38",
          7734 => x"7c",
          7735 => x"0c",
          7736 => x"81",
          7737 => x"74",
          7738 => x"7a",
          7739 => x"0c",
          7740 => x"04",
          7741 => x"79",
          7742 => x"05",
          7743 => x"57",
          7744 => x"82",
          7745 => x"56",
          7746 => x"08",
          7747 => x"91",
          7748 => x"75",
          7749 => x"90",
          7750 => x"81",
          7751 => x"06",
          7752 => x"87",
          7753 => x"2e",
          7754 => x"94",
          7755 => x"73",
          7756 => x"27",
          7757 => x"73",
          7758 => x"b5",
          7759 => x"88",
          7760 => x"76",
          7761 => x"3f",
          7762 => x"08",
          7763 => x"0c",
          7764 => x"39",
          7765 => x"52",
          7766 => x"bf",
          7767 => x"b5",
          7768 => x"2e",
          7769 => x"83",
          7770 => x"82",
          7771 => x"81",
          7772 => x"06",
          7773 => x"56",
          7774 => x"a0",
          7775 => x"82",
          7776 => x"98",
          7777 => x"94",
          7778 => x"08",
          7779 => x"a8",
          7780 => x"51",
          7781 => x"82",
          7782 => x"56",
          7783 => x"8c",
          7784 => x"17",
          7785 => x"07",
          7786 => x"18",
          7787 => x"2e",
          7788 => x"91",
          7789 => x"55",
          7790 => x"a8",
          7791 => x"0d",
          7792 => x"0d",
          7793 => x"3d",
          7794 => x"52",
          7795 => x"da",
          7796 => x"b5",
          7797 => x"82",
          7798 => x"81",
          7799 => x"45",
          7800 => x"52",
          7801 => x"52",
          7802 => x"3f",
          7803 => x"08",
          7804 => x"a8",
          7805 => x"38",
          7806 => x"05",
          7807 => x"2a",
          7808 => x"51",
          7809 => x"55",
          7810 => x"38",
          7811 => x"54",
          7812 => x"81",
          7813 => x"80",
          7814 => x"70",
          7815 => x"54",
          7816 => x"81",
          7817 => x"52",
          7818 => x"c5",
          7819 => x"a8",
          7820 => x"2a",
          7821 => x"51",
          7822 => x"80",
          7823 => x"38",
          7824 => x"b5",
          7825 => x"15",
          7826 => x"86",
          7827 => x"82",
          7828 => x"5c",
          7829 => x"3d",
          7830 => x"c7",
          7831 => x"b5",
          7832 => x"82",
          7833 => x"80",
          7834 => x"b5",
          7835 => x"73",
          7836 => x"3f",
          7837 => x"08",
          7838 => x"a8",
          7839 => x"87",
          7840 => x"39",
          7841 => x"08",
          7842 => x"38",
          7843 => x"08",
          7844 => x"77",
          7845 => x"3f",
          7846 => x"08",
          7847 => x"08",
          7848 => x"b5",
          7849 => x"80",
          7850 => x"55",
          7851 => x"94",
          7852 => x"2e",
          7853 => x"53",
          7854 => x"51",
          7855 => x"82",
          7856 => x"55",
          7857 => x"78",
          7858 => x"fe",
          7859 => x"a8",
          7860 => x"82",
          7861 => x"a0",
          7862 => x"e9",
          7863 => x"53",
          7864 => x"05",
          7865 => x"51",
          7866 => x"82",
          7867 => x"54",
          7868 => x"08",
          7869 => x"78",
          7870 => x"8e",
          7871 => x"58",
          7872 => x"82",
          7873 => x"54",
          7874 => x"08",
          7875 => x"54",
          7876 => x"82",
          7877 => x"84",
          7878 => x"06",
          7879 => x"02",
          7880 => x"33",
          7881 => x"81",
          7882 => x"86",
          7883 => x"f6",
          7884 => x"74",
          7885 => x"70",
          7886 => x"c3",
          7887 => x"a8",
          7888 => x"56",
          7889 => x"08",
          7890 => x"54",
          7891 => x"08",
          7892 => x"81",
          7893 => x"82",
          7894 => x"a8",
          7895 => x"09",
          7896 => x"38",
          7897 => x"b4",
          7898 => x"b0",
          7899 => x"a8",
          7900 => x"51",
          7901 => x"82",
          7902 => x"54",
          7903 => x"08",
          7904 => x"8b",
          7905 => x"b4",
          7906 => x"b7",
          7907 => x"54",
          7908 => x"15",
          7909 => x"90",
          7910 => x"34",
          7911 => x"0a",
          7912 => x"19",
          7913 => x"9f",
          7914 => x"78",
          7915 => x"51",
          7916 => x"a0",
          7917 => x"11",
          7918 => x"05",
          7919 => x"b6",
          7920 => x"ae",
          7921 => x"15",
          7922 => x"78",
          7923 => x"53",
          7924 => x"3f",
          7925 => x"0b",
          7926 => x"77",
          7927 => x"3f",
          7928 => x"08",
          7929 => x"a8",
          7930 => x"82",
          7931 => x"52",
          7932 => x"51",
          7933 => x"3f",
          7934 => x"52",
          7935 => x"aa",
          7936 => x"90",
          7937 => x"34",
          7938 => x"0b",
          7939 => x"78",
          7940 => x"b6",
          7941 => x"a8",
          7942 => x"39",
          7943 => x"52",
          7944 => x"be",
          7945 => x"82",
          7946 => x"99",
          7947 => x"da",
          7948 => x"3d",
          7949 => x"d2",
          7950 => x"53",
          7951 => x"84",
          7952 => x"3d",
          7953 => x"3f",
          7954 => x"08",
          7955 => x"a8",
          7956 => x"38",
          7957 => x"3d",
          7958 => x"3d",
          7959 => x"cc",
          7960 => x"b5",
          7961 => x"82",
          7962 => x"82",
          7963 => x"81",
          7964 => x"81",
          7965 => x"86",
          7966 => x"aa",
          7967 => x"a4",
          7968 => x"a8",
          7969 => x"05",
          7970 => x"ea",
          7971 => x"77",
          7972 => x"70",
          7973 => x"b4",
          7974 => x"3d",
          7975 => x"51",
          7976 => x"82",
          7977 => x"55",
          7978 => x"08",
          7979 => x"6f",
          7980 => x"06",
          7981 => x"a2",
          7982 => x"92",
          7983 => x"81",
          7984 => x"b5",
          7985 => x"2e",
          7986 => x"81",
          7987 => x"51",
          7988 => x"82",
          7989 => x"55",
          7990 => x"08",
          7991 => x"68",
          7992 => x"a8",
          7993 => x"05",
          7994 => x"51",
          7995 => x"3f",
          7996 => x"33",
          7997 => x"8b",
          7998 => x"84",
          7999 => x"06",
          8000 => x"73",
          8001 => x"a0",
          8002 => x"8b",
          8003 => x"54",
          8004 => x"15",
          8005 => x"33",
          8006 => x"70",
          8007 => x"55",
          8008 => x"2e",
          8009 => x"6e",
          8010 => x"df",
          8011 => x"78",
          8012 => x"3f",
          8013 => x"08",
          8014 => x"ff",
          8015 => x"82",
          8016 => x"a8",
          8017 => x"80",
          8018 => x"b5",
          8019 => x"78",
          8020 => x"af",
          8021 => x"a8",
          8022 => x"d4",
          8023 => x"55",
          8024 => x"08",
          8025 => x"81",
          8026 => x"73",
          8027 => x"81",
          8028 => x"63",
          8029 => x"76",
          8030 => x"3f",
          8031 => x"0b",
          8032 => x"87",
          8033 => x"a8",
          8034 => x"77",
          8035 => x"3f",
          8036 => x"08",
          8037 => x"a8",
          8038 => x"78",
          8039 => x"aa",
          8040 => x"a8",
          8041 => x"82",
          8042 => x"a8",
          8043 => x"ed",
          8044 => x"80",
          8045 => x"02",
          8046 => x"df",
          8047 => x"57",
          8048 => x"3d",
          8049 => x"96",
          8050 => x"e9",
          8051 => x"a8",
          8052 => x"b5",
          8053 => x"cf",
          8054 => x"65",
          8055 => x"d4",
          8056 => x"b5",
          8057 => x"a8",
          8058 => x"b5",
          8059 => x"38",
          8060 => x"05",
          8061 => x"06",
          8062 => x"73",
          8063 => x"a7",
          8064 => x"09",
          8065 => x"71",
          8066 => x"06",
          8067 => x"55",
          8068 => x"15",
          8069 => x"81",
          8070 => x"34",
          8071 => x"b4",
          8072 => x"b5",
          8073 => x"74",
          8074 => x"0c",
          8075 => x"04",
          8076 => x"64",
          8077 => x"93",
          8078 => x"52",
          8079 => x"d1",
          8080 => x"b5",
          8081 => x"82",
          8082 => x"80",
          8083 => x"58",
          8084 => x"3d",
          8085 => x"c8",
          8086 => x"b5",
          8087 => x"82",
          8088 => x"b4",
          8089 => x"c7",
          8090 => x"a0",
          8091 => x"55",
          8092 => x"84",
          8093 => x"17",
          8094 => x"2b",
          8095 => x"96",
          8096 => x"b0",
          8097 => x"54",
          8098 => x"15",
          8099 => x"ff",
          8100 => x"82",
          8101 => x"55",
          8102 => x"a8",
          8103 => x"0d",
          8104 => x"0d",
          8105 => x"5a",
          8106 => x"3d",
          8107 => x"99",
          8108 => x"81",
          8109 => x"a8",
          8110 => x"a8",
          8111 => x"82",
          8112 => x"07",
          8113 => x"55",
          8114 => x"2e",
          8115 => x"81",
          8116 => x"55",
          8117 => x"2e",
          8118 => x"7b",
          8119 => x"80",
          8120 => x"70",
          8121 => x"be",
          8122 => x"b5",
          8123 => x"82",
          8124 => x"80",
          8125 => x"52",
          8126 => x"dc",
          8127 => x"a8",
          8128 => x"b5",
          8129 => x"38",
          8130 => x"08",
          8131 => x"08",
          8132 => x"56",
          8133 => x"19",
          8134 => x"59",
          8135 => x"74",
          8136 => x"56",
          8137 => x"ec",
          8138 => x"75",
          8139 => x"74",
          8140 => x"2e",
          8141 => x"16",
          8142 => x"33",
          8143 => x"73",
          8144 => x"38",
          8145 => x"84",
          8146 => x"06",
          8147 => x"7a",
          8148 => x"76",
          8149 => x"07",
          8150 => x"54",
          8151 => x"80",
          8152 => x"80",
          8153 => x"7b",
          8154 => x"53",
          8155 => x"93",
          8156 => x"a8",
          8157 => x"b5",
          8158 => x"38",
          8159 => x"55",
          8160 => x"56",
          8161 => x"8b",
          8162 => x"56",
          8163 => x"83",
          8164 => x"75",
          8165 => x"51",
          8166 => x"3f",
          8167 => x"08",
          8168 => x"82",
          8169 => x"98",
          8170 => x"e6",
          8171 => x"53",
          8172 => x"b8",
          8173 => x"3d",
          8174 => x"3f",
          8175 => x"08",
          8176 => x"08",
          8177 => x"b5",
          8178 => x"98",
          8179 => x"a0",
          8180 => x"70",
          8181 => x"ae",
          8182 => x"6d",
          8183 => x"81",
          8184 => x"57",
          8185 => x"74",
          8186 => x"38",
          8187 => x"81",
          8188 => x"81",
          8189 => x"52",
          8190 => x"89",
          8191 => x"a8",
          8192 => x"a5",
          8193 => x"33",
          8194 => x"54",
          8195 => x"3f",
          8196 => x"08",
          8197 => x"38",
          8198 => x"76",
          8199 => x"05",
          8200 => x"39",
          8201 => x"08",
          8202 => x"15",
          8203 => x"ff",
          8204 => x"73",
          8205 => x"38",
          8206 => x"83",
          8207 => x"56",
          8208 => x"75",
          8209 => x"82",
          8210 => x"33",
          8211 => x"2e",
          8212 => x"52",
          8213 => x"51",
          8214 => x"3f",
          8215 => x"08",
          8216 => x"ff",
          8217 => x"38",
          8218 => x"88",
          8219 => x"8a",
          8220 => x"38",
          8221 => x"ec",
          8222 => x"75",
          8223 => x"74",
          8224 => x"73",
          8225 => x"05",
          8226 => x"17",
          8227 => x"70",
          8228 => x"34",
          8229 => x"70",
          8230 => x"ff",
          8231 => x"55",
          8232 => x"26",
          8233 => x"8b",
          8234 => x"86",
          8235 => x"e5",
          8236 => x"38",
          8237 => x"99",
          8238 => x"05",
          8239 => x"70",
          8240 => x"73",
          8241 => x"81",
          8242 => x"ff",
          8243 => x"ed",
          8244 => x"80",
          8245 => x"91",
          8246 => x"55",
          8247 => x"3f",
          8248 => x"08",
          8249 => x"a8",
          8250 => x"38",
          8251 => x"51",
          8252 => x"3f",
          8253 => x"08",
          8254 => x"a8",
          8255 => x"76",
          8256 => x"67",
          8257 => x"34",
          8258 => x"82",
          8259 => x"84",
          8260 => x"06",
          8261 => x"80",
          8262 => x"2e",
          8263 => x"81",
          8264 => x"ff",
          8265 => x"82",
          8266 => x"54",
          8267 => x"08",
          8268 => x"53",
          8269 => x"08",
          8270 => x"ff",
          8271 => x"67",
          8272 => x"8b",
          8273 => x"53",
          8274 => x"51",
          8275 => x"3f",
          8276 => x"0b",
          8277 => x"79",
          8278 => x"ee",
          8279 => x"a8",
          8280 => x"55",
          8281 => x"a8",
          8282 => x"0d",
          8283 => x"0d",
          8284 => x"88",
          8285 => x"05",
          8286 => x"fc",
          8287 => x"54",
          8288 => x"d2",
          8289 => x"b5",
          8290 => x"82",
          8291 => x"82",
          8292 => x"1a",
          8293 => x"82",
          8294 => x"80",
          8295 => x"8c",
          8296 => x"78",
          8297 => x"1a",
          8298 => x"2a",
          8299 => x"51",
          8300 => x"90",
          8301 => x"82",
          8302 => x"58",
          8303 => x"81",
          8304 => x"39",
          8305 => x"22",
          8306 => x"70",
          8307 => x"56",
          8308 => x"ce",
          8309 => x"14",
          8310 => x"30",
          8311 => x"9f",
          8312 => x"a8",
          8313 => x"19",
          8314 => x"5a",
          8315 => x"81",
          8316 => x"38",
          8317 => x"77",
          8318 => x"82",
          8319 => x"56",
          8320 => x"74",
          8321 => x"ff",
          8322 => x"81",
          8323 => x"55",
          8324 => x"75",
          8325 => x"82",
          8326 => x"a8",
          8327 => x"ff",
          8328 => x"b5",
          8329 => x"2e",
          8330 => x"82",
          8331 => x"8e",
          8332 => x"56",
          8333 => x"09",
          8334 => x"38",
          8335 => x"59",
          8336 => x"77",
          8337 => x"06",
          8338 => x"87",
          8339 => x"39",
          8340 => x"ba",
          8341 => x"55",
          8342 => x"2e",
          8343 => x"15",
          8344 => x"2e",
          8345 => x"83",
          8346 => x"75",
          8347 => x"7e",
          8348 => x"a8",
          8349 => x"a8",
          8350 => x"b5",
          8351 => x"ce",
          8352 => x"16",
          8353 => x"56",
          8354 => x"38",
          8355 => x"19",
          8356 => x"8c",
          8357 => x"7d",
          8358 => x"38",
          8359 => x"0c",
          8360 => x"0c",
          8361 => x"80",
          8362 => x"73",
          8363 => x"98",
          8364 => x"05",
          8365 => x"57",
          8366 => x"26",
          8367 => x"7b",
          8368 => x"0c",
          8369 => x"81",
          8370 => x"84",
          8371 => x"54",
          8372 => x"a8",
          8373 => x"0d",
          8374 => x"0d",
          8375 => x"88",
          8376 => x"05",
          8377 => x"54",
          8378 => x"c5",
          8379 => x"56",
          8380 => x"b5",
          8381 => x"8b",
          8382 => x"b5",
          8383 => x"29",
          8384 => x"05",
          8385 => x"55",
          8386 => x"84",
          8387 => x"34",
          8388 => x"08",
          8389 => x"5f",
          8390 => x"51",
          8391 => x"3f",
          8392 => x"08",
          8393 => x"70",
          8394 => x"57",
          8395 => x"8b",
          8396 => x"82",
          8397 => x"06",
          8398 => x"56",
          8399 => x"38",
          8400 => x"05",
          8401 => x"7e",
          8402 => x"f0",
          8403 => x"a8",
          8404 => x"67",
          8405 => x"2e",
          8406 => x"82",
          8407 => x"8b",
          8408 => x"75",
          8409 => x"80",
          8410 => x"81",
          8411 => x"2e",
          8412 => x"80",
          8413 => x"38",
          8414 => x"0a",
          8415 => x"ff",
          8416 => x"55",
          8417 => x"86",
          8418 => x"8a",
          8419 => x"89",
          8420 => x"2a",
          8421 => x"77",
          8422 => x"59",
          8423 => x"81",
          8424 => x"70",
          8425 => x"07",
          8426 => x"56",
          8427 => x"38",
          8428 => x"05",
          8429 => x"7e",
          8430 => x"80",
          8431 => x"82",
          8432 => x"8a",
          8433 => x"83",
          8434 => x"06",
          8435 => x"08",
          8436 => x"74",
          8437 => x"41",
          8438 => x"56",
          8439 => x"8a",
          8440 => x"61",
          8441 => x"55",
          8442 => x"27",
          8443 => x"93",
          8444 => x"80",
          8445 => x"38",
          8446 => x"70",
          8447 => x"43",
          8448 => x"95",
          8449 => x"06",
          8450 => x"2e",
          8451 => x"77",
          8452 => x"74",
          8453 => x"83",
          8454 => x"06",
          8455 => x"82",
          8456 => x"2e",
          8457 => x"78",
          8458 => x"2e",
          8459 => x"80",
          8460 => x"ae",
          8461 => x"2a",
          8462 => x"82",
          8463 => x"56",
          8464 => x"2e",
          8465 => x"77",
          8466 => x"82",
          8467 => x"79",
          8468 => x"70",
          8469 => x"5a",
          8470 => x"86",
          8471 => x"27",
          8472 => x"52",
          8473 => x"c9",
          8474 => x"b5",
          8475 => x"29",
          8476 => x"70",
          8477 => x"55",
          8478 => x"0b",
          8479 => x"08",
          8480 => x"05",
          8481 => x"ff",
          8482 => x"27",
          8483 => x"88",
          8484 => x"ae",
          8485 => x"2a",
          8486 => x"82",
          8487 => x"56",
          8488 => x"2e",
          8489 => x"77",
          8490 => x"82",
          8491 => x"79",
          8492 => x"70",
          8493 => x"5a",
          8494 => x"86",
          8495 => x"27",
          8496 => x"52",
          8497 => x"c8",
          8498 => x"b5",
          8499 => x"84",
          8500 => x"b5",
          8501 => x"f5",
          8502 => x"81",
          8503 => x"a8",
          8504 => x"b5",
          8505 => x"71",
          8506 => x"83",
          8507 => x"5e",
          8508 => x"89",
          8509 => x"5c",
          8510 => x"1c",
          8511 => x"05",
          8512 => x"ff",
          8513 => x"70",
          8514 => x"31",
          8515 => x"57",
          8516 => x"83",
          8517 => x"06",
          8518 => x"1c",
          8519 => x"5c",
          8520 => x"1d",
          8521 => x"29",
          8522 => x"31",
          8523 => x"55",
          8524 => x"87",
          8525 => x"7c",
          8526 => x"7a",
          8527 => x"31",
          8528 => x"c7",
          8529 => x"b5",
          8530 => x"7d",
          8531 => x"81",
          8532 => x"82",
          8533 => x"83",
          8534 => x"80",
          8535 => x"87",
          8536 => x"81",
          8537 => x"fd",
          8538 => x"f8",
          8539 => x"2e",
          8540 => x"80",
          8541 => x"ff",
          8542 => x"b5",
          8543 => x"a0",
          8544 => x"38",
          8545 => x"74",
          8546 => x"86",
          8547 => x"fd",
          8548 => x"81",
          8549 => x"80",
          8550 => x"83",
          8551 => x"39",
          8552 => x"08",
          8553 => x"92",
          8554 => x"b8",
          8555 => x"59",
          8556 => x"27",
          8557 => x"86",
          8558 => x"55",
          8559 => x"09",
          8560 => x"38",
          8561 => x"f5",
          8562 => x"38",
          8563 => x"55",
          8564 => x"86",
          8565 => x"80",
          8566 => x"7a",
          8567 => x"b9",
          8568 => x"82",
          8569 => x"7a",
          8570 => x"8a",
          8571 => x"52",
          8572 => x"ff",
          8573 => x"79",
          8574 => x"7b",
          8575 => x"06",
          8576 => x"51",
          8577 => x"3f",
          8578 => x"1c",
          8579 => x"32",
          8580 => x"96",
          8581 => x"06",
          8582 => x"91",
          8583 => x"a1",
          8584 => x"55",
          8585 => x"ff",
          8586 => x"74",
          8587 => x"06",
          8588 => x"51",
          8589 => x"3f",
          8590 => x"52",
          8591 => x"ff",
          8592 => x"f8",
          8593 => x"34",
          8594 => x"1b",
          8595 => x"d9",
          8596 => x"52",
          8597 => x"ff",
          8598 => x"60",
          8599 => x"51",
          8600 => x"3f",
          8601 => x"09",
          8602 => x"cb",
          8603 => x"b2",
          8604 => x"c3",
          8605 => x"a0",
          8606 => x"52",
          8607 => x"ff",
          8608 => x"82",
          8609 => x"51",
          8610 => x"3f",
          8611 => x"1b",
          8612 => x"95",
          8613 => x"b2",
          8614 => x"a0",
          8615 => x"80",
          8616 => x"1c",
          8617 => x"80",
          8618 => x"93",
          8619 => x"b8",
          8620 => x"1b",
          8621 => x"82",
          8622 => x"52",
          8623 => x"ff",
          8624 => x"7c",
          8625 => x"06",
          8626 => x"51",
          8627 => x"3f",
          8628 => x"a4",
          8629 => x"0b",
          8630 => x"93",
          8631 => x"cc",
          8632 => x"51",
          8633 => x"3f",
          8634 => x"52",
          8635 => x"70",
          8636 => x"9f",
          8637 => x"54",
          8638 => x"52",
          8639 => x"9b",
          8640 => x"56",
          8641 => x"08",
          8642 => x"7d",
          8643 => x"81",
          8644 => x"38",
          8645 => x"86",
          8646 => x"52",
          8647 => x"9b",
          8648 => x"80",
          8649 => x"7a",
          8650 => x"ed",
          8651 => x"85",
          8652 => x"7a",
          8653 => x"8f",
          8654 => x"85",
          8655 => x"83",
          8656 => x"ff",
          8657 => x"ff",
          8658 => x"e8",
          8659 => x"9e",
          8660 => x"52",
          8661 => x"51",
          8662 => x"3f",
          8663 => x"52",
          8664 => x"9e",
          8665 => x"54",
          8666 => x"53",
          8667 => x"51",
          8668 => x"3f",
          8669 => x"16",
          8670 => x"7e",
          8671 => x"d8",
          8672 => x"80",
          8673 => x"ff",
          8674 => x"7f",
          8675 => x"7d",
          8676 => x"81",
          8677 => x"f8",
          8678 => x"ff",
          8679 => x"ff",
          8680 => x"51",
          8681 => x"3f",
          8682 => x"88",
          8683 => x"39",
          8684 => x"f8",
          8685 => x"2e",
          8686 => x"55",
          8687 => x"51",
          8688 => x"3f",
          8689 => x"57",
          8690 => x"83",
          8691 => x"76",
          8692 => x"7a",
          8693 => x"ff",
          8694 => x"82",
          8695 => x"82",
          8696 => x"80",
          8697 => x"a8",
          8698 => x"51",
          8699 => x"3f",
          8700 => x"78",
          8701 => x"74",
          8702 => x"18",
          8703 => x"2e",
          8704 => x"79",
          8705 => x"2e",
          8706 => x"55",
          8707 => x"62",
          8708 => x"74",
          8709 => x"75",
          8710 => x"7e",
          8711 => x"b8",
          8712 => x"a8",
          8713 => x"38",
          8714 => x"78",
          8715 => x"74",
          8716 => x"56",
          8717 => x"93",
          8718 => x"66",
          8719 => x"26",
          8720 => x"56",
          8721 => x"83",
          8722 => x"64",
          8723 => x"77",
          8724 => x"84",
          8725 => x"52",
          8726 => x"9d",
          8727 => x"d4",
          8728 => x"51",
          8729 => x"3f",
          8730 => x"55",
          8731 => x"81",
          8732 => x"34",
          8733 => x"16",
          8734 => x"16",
          8735 => x"16",
          8736 => x"05",
          8737 => x"c1",
          8738 => x"fe",
          8739 => x"fe",
          8740 => x"34",
          8741 => x"08",
          8742 => x"07",
          8743 => x"16",
          8744 => x"a8",
          8745 => x"34",
          8746 => x"c6",
          8747 => x"9c",
          8748 => x"52",
          8749 => x"51",
          8750 => x"3f",
          8751 => x"53",
          8752 => x"51",
          8753 => x"3f",
          8754 => x"b5",
          8755 => x"38",
          8756 => x"52",
          8757 => x"99",
          8758 => x"56",
          8759 => x"08",
          8760 => x"39",
          8761 => x"39",
          8762 => x"39",
          8763 => x"08",
          8764 => x"b5",
          8765 => x"3d",
          8766 => x"3d",
          8767 => x"5b",
          8768 => x"60",
          8769 => x"57",
          8770 => x"25",
          8771 => x"3d",
          8772 => x"55",
          8773 => x"15",
          8774 => x"c9",
          8775 => x"81",
          8776 => x"06",
          8777 => x"3d",
          8778 => x"8d",
          8779 => x"74",
          8780 => x"05",
          8781 => x"17",
          8782 => x"2e",
          8783 => x"c9",
          8784 => x"34",
          8785 => x"83",
          8786 => x"74",
          8787 => x"0c",
          8788 => x"04",
          8789 => x"7b",
          8790 => x"b3",
          8791 => x"57",
          8792 => x"09",
          8793 => x"38",
          8794 => x"51",
          8795 => x"17",
          8796 => x"76",
          8797 => x"88",
          8798 => x"17",
          8799 => x"59",
          8800 => x"81",
          8801 => x"76",
          8802 => x"8b",
          8803 => x"54",
          8804 => x"17",
          8805 => x"51",
          8806 => x"79",
          8807 => x"30",
          8808 => x"9f",
          8809 => x"53",
          8810 => x"75",
          8811 => x"81",
          8812 => x"0c",
          8813 => x"04",
          8814 => x"79",
          8815 => x"56",
          8816 => x"24",
          8817 => x"3d",
          8818 => x"74",
          8819 => x"52",
          8820 => x"cb",
          8821 => x"b5",
          8822 => x"38",
          8823 => x"78",
          8824 => x"06",
          8825 => x"16",
          8826 => x"39",
          8827 => x"82",
          8828 => x"89",
          8829 => x"fd",
          8830 => x"54",
          8831 => x"80",
          8832 => x"ff",
          8833 => x"76",
          8834 => x"3d",
          8835 => x"3d",
          8836 => x"e3",
          8837 => x"53",
          8838 => x"53",
          8839 => x"3f",
          8840 => x"51",
          8841 => x"72",
          8842 => x"3f",
          8843 => x"04",
          8844 => x"00",
          8845 => x"ff",
          8846 => x"ff",
          8847 => x"ff",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"64",
          8985 => x"74",
          8986 => x"64",
          8987 => x"74",
          8988 => x"66",
          8989 => x"74",
          8990 => x"66",
          8991 => x"64",
          8992 => x"66",
          8993 => x"63",
          8994 => x"6d",
          8995 => x"61",
          8996 => x"6d",
          8997 => x"79",
          8998 => x"6d",
          8999 => x"66",
          9000 => x"6d",
          9001 => x"70",
          9002 => x"6d",
          9003 => x"6d",
          9004 => x"6d",
          9005 => x"68",
          9006 => x"68",
          9007 => x"68",
          9008 => x"68",
          9009 => x"63",
          9010 => x"00",
          9011 => x"6a",
          9012 => x"72",
          9013 => x"61",
          9014 => x"72",
          9015 => x"74",
          9016 => x"69",
          9017 => x"00",
          9018 => x"74",
          9019 => x"00",
          9020 => x"74",
          9021 => x"69",
          9022 => x"6d",
          9023 => x"69",
          9024 => x"6b",
          9025 => x"00",
          9026 => x"65",
          9027 => x"44",
          9028 => x"20",
          9029 => x"6f",
          9030 => x"49",
          9031 => x"72",
          9032 => x"20",
          9033 => x"6f",
          9034 => x"00",
          9035 => x"44",
          9036 => x"20",
          9037 => x"20",
          9038 => x"64",
          9039 => x"00",
          9040 => x"4e",
          9041 => x"69",
          9042 => x"66",
          9043 => x"64",
          9044 => x"4e",
          9045 => x"61",
          9046 => x"66",
          9047 => x"64",
          9048 => x"49",
          9049 => x"6c",
          9050 => x"66",
          9051 => x"6e",
          9052 => x"2e",
          9053 => x"41",
          9054 => x"73",
          9055 => x"65",
          9056 => x"64",
          9057 => x"46",
          9058 => x"20",
          9059 => x"65",
          9060 => x"20",
          9061 => x"73",
          9062 => x"0a",
          9063 => x"46",
          9064 => x"20",
          9065 => x"64",
          9066 => x"69",
          9067 => x"6c",
          9068 => x"0a",
          9069 => x"53",
          9070 => x"73",
          9071 => x"69",
          9072 => x"70",
          9073 => x"65",
          9074 => x"64",
          9075 => x"44",
          9076 => x"65",
          9077 => x"6d",
          9078 => x"20",
          9079 => x"69",
          9080 => x"6c",
          9081 => x"0a",
          9082 => x"44",
          9083 => x"20",
          9084 => x"20",
          9085 => x"62",
          9086 => x"2e",
          9087 => x"4e",
          9088 => x"6f",
          9089 => x"74",
          9090 => x"65",
          9091 => x"6c",
          9092 => x"73",
          9093 => x"20",
          9094 => x"6e",
          9095 => x"6e",
          9096 => x"73",
          9097 => x"00",
          9098 => x"46",
          9099 => x"61",
          9100 => x"62",
          9101 => x"65",
          9102 => x"00",
          9103 => x"54",
          9104 => x"6f",
          9105 => x"20",
          9106 => x"72",
          9107 => x"6f",
          9108 => x"61",
          9109 => x"6c",
          9110 => x"2e",
          9111 => x"46",
          9112 => x"20",
          9113 => x"6c",
          9114 => x"65",
          9115 => x"00",
          9116 => x"49",
          9117 => x"66",
          9118 => x"69",
          9119 => x"20",
          9120 => x"6f",
          9121 => x"0a",
          9122 => x"54",
          9123 => x"6d",
          9124 => x"20",
          9125 => x"6e",
          9126 => x"6c",
          9127 => x"0a",
          9128 => x"50",
          9129 => x"6d",
          9130 => x"72",
          9131 => x"6e",
          9132 => x"72",
          9133 => x"2e",
          9134 => x"53",
          9135 => x"65",
          9136 => x"0a",
          9137 => x"55",
          9138 => x"6f",
          9139 => x"65",
          9140 => x"72",
          9141 => x"0a",
          9142 => x"20",
          9143 => x"65",
          9144 => x"73",
          9145 => x"20",
          9146 => x"20",
          9147 => x"65",
          9148 => x"65",
          9149 => x"00",
          9150 => x"72",
          9151 => x"00",
          9152 => x"25",
          9153 => x"00",
          9154 => x"3a",
          9155 => x"25",
          9156 => x"00",
          9157 => x"20",
          9158 => x"20",
          9159 => x"00",
          9160 => x"25",
          9161 => x"00",
          9162 => x"20",
          9163 => x"20",
          9164 => x"7c",
          9165 => x"7a",
          9166 => x"0a",
          9167 => x"25",
          9168 => x"00",
          9169 => x"30",
          9170 => x"35",
          9171 => x"32",
          9172 => x"76",
          9173 => x"32",
          9174 => x"20",
          9175 => x"2c",
          9176 => x"76",
          9177 => x"32",
          9178 => x"25",
          9179 => x"73",
          9180 => x"0a",
          9181 => x"5a",
          9182 => x"49",
          9183 => x"72",
          9184 => x"74",
          9185 => x"6e",
          9186 => x"72",
          9187 => x"54",
          9188 => x"72",
          9189 => x"74",
          9190 => x"75",
          9191 => x"00",
          9192 => x"50",
          9193 => x"69",
          9194 => x"72",
          9195 => x"74",
          9196 => x"49",
          9197 => x"4c",
          9198 => x"20",
          9199 => x"65",
          9200 => x"70",
          9201 => x"49",
          9202 => x"4c",
          9203 => x"20",
          9204 => x"65",
          9205 => x"70",
          9206 => x"55",
          9207 => x"30",
          9208 => x"20",
          9209 => x"65",
          9210 => x"70",
          9211 => x"55",
          9212 => x"30",
          9213 => x"20",
          9214 => x"65",
          9215 => x"70",
          9216 => x"55",
          9217 => x"31",
          9218 => x"20",
          9219 => x"65",
          9220 => x"70",
          9221 => x"55",
          9222 => x"31",
          9223 => x"20",
          9224 => x"65",
          9225 => x"70",
          9226 => x"53",
          9227 => x"69",
          9228 => x"75",
          9229 => x"69",
          9230 => x"2e",
          9231 => x"00",
          9232 => x"45",
          9233 => x"6c",
          9234 => x"20",
          9235 => x"65",
          9236 => x"2e",
          9237 => x"61",
          9238 => x"65",
          9239 => x"2e",
          9240 => x"00",
          9241 => x"7a",
          9242 => x"68",
          9243 => x"30",
          9244 => x"46",
          9245 => x"65",
          9246 => x"6f",
          9247 => x"69",
          9248 => x"6c",
          9249 => x"20",
          9250 => x"63",
          9251 => x"20",
          9252 => x"70",
          9253 => x"73",
          9254 => x"6e",
          9255 => x"6d",
          9256 => x"61",
          9257 => x"2e",
          9258 => x"2a",
          9259 => x"43",
          9260 => x"72",
          9261 => x"2e",
          9262 => x"00",
          9263 => x"43",
          9264 => x"69",
          9265 => x"2e",
          9266 => x"43",
          9267 => x"61",
          9268 => x"67",
          9269 => x"00",
          9270 => x"25",
          9271 => x"78",
          9272 => x"38",
          9273 => x"3e",
          9274 => x"6c",
          9275 => x"30",
          9276 => x"0a",
          9277 => x"44",
          9278 => x"20",
          9279 => x"6f",
          9280 => x"00",
          9281 => x"0a",
          9282 => x"70",
          9283 => x"65",
          9284 => x"25",
          9285 => x"20",
          9286 => x"58",
          9287 => x"3f",
          9288 => x"00",
          9289 => x"25",
          9290 => x"20",
          9291 => x"58",
          9292 => x"25",
          9293 => x"20",
          9294 => x"58",
          9295 => x"45",
          9296 => x"75",
          9297 => x"67",
          9298 => x"64",
          9299 => x"20",
          9300 => x"78",
          9301 => x"2e",
          9302 => x"43",
          9303 => x"69",
          9304 => x"63",
          9305 => x"20",
          9306 => x"30",
          9307 => x"2e",
          9308 => x"00",
          9309 => x"43",
          9310 => x"20",
          9311 => x"75",
          9312 => x"64",
          9313 => x"64",
          9314 => x"25",
          9315 => x"0a",
          9316 => x"52",
          9317 => x"61",
          9318 => x"6e",
          9319 => x"70",
          9320 => x"63",
          9321 => x"6f",
          9322 => x"2e",
          9323 => x"43",
          9324 => x"20",
          9325 => x"6f",
          9326 => x"6e",
          9327 => x"2e",
          9328 => x"5a",
          9329 => x"62",
          9330 => x"25",
          9331 => x"25",
          9332 => x"73",
          9333 => x"00",
          9334 => x"25",
          9335 => x"25",
          9336 => x"73",
          9337 => x"25",
          9338 => x"25",
          9339 => x"42",
          9340 => x"63",
          9341 => x"61",
          9342 => x"00",
          9343 => x"48",
          9344 => x"4f",
          9345 => x"46",
          9346 => x"20",
          9347 => x"4e",
          9348 => x"48",
          9349 => x"4f",
          9350 => x"46",
          9351 => x"20",
          9352 => x"4e",
          9353 => x"52",
          9354 => x"69",
          9355 => x"2e",
          9356 => x"45",
          9357 => x"6c",
          9358 => x"20",
          9359 => x"65",
          9360 => x"70",
          9361 => x"2e",
          9362 => x"25",
          9363 => x"64",
          9364 => x"20",
          9365 => x"25",
          9366 => x"64",
          9367 => x"25",
          9368 => x"53",
          9369 => x"43",
          9370 => x"69",
          9371 => x"61",
          9372 => x"6e",
          9373 => x"20",
          9374 => x"6f",
          9375 => x"6f",
          9376 => x"6f",
          9377 => x"67",
          9378 => x"3a",
          9379 => x"76",
          9380 => x"73",
          9381 => x"70",
          9382 => x"65",
          9383 => x"64",
          9384 => x"20",
          9385 => x"57",
          9386 => x"44",
          9387 => x"20",
          9388 => x"30",
          9389 => x"25",
          9390 => x"29",
          9391 => x"20",
          9392 => x"53",
          9393 => x"4d",
          9394 => x"20",
          9395 => x"30",
          9396 => x"25",
          9397 => x"29",
          9398 => x"20",
          9399 => x"49",
          9400 => x"20",
          9401 => x"4d",
          9402 => x"30",
          9403 => x"25",
          9404 => x"29",
          9405 => x"20",
          9406 => x"42",
          9407 => x"20",
          9408 => x"20",
          9409 => x"30",
          9410 => x"25",
          9411 => x"29",
          9412 => x"20",
          9413 => x"52",
          9414 => x"20",
          9415 => x"20",
          9416 => x"30",
          9417 => x"25",
          9418 => x"29",
          9419 => x"20",
          9420 => x"53",
          9421 => x"41",
          9422 => x"20",
          9423 => x"65",
          9424 => x"65",
          9425 => x"25",
          9426 => x"29",
          9427 => x"20",
          9428 => x"54",
          9429 => x"52",
          9430 => x"20",
          9431 => x"69",
          9432 => x"73",
          9433 => x"25",
          9434 => x"29",
          9435 => x"20",
          9436 => x"49",
          9437 => x"20",
          9438 => x"4c",
          9439 => x"68",
          9440 => x"65",
          9441 => x"25",
          9442 => x"29",
          9443 => x"20",
          9444 => x"57",
          9445 => x"42",
          9446 => x"20",
          9447 => x"0a",
          9448 => x"20",
          9449 => x"57",
          9450 => x"32",
          9451 => x"20",
          9452 => x"49",
          9453 => x"4c",
          9454 => x"20",
          9455 => x"50",
          9456 => x"00",
          9457 => x"20",
          9458 => x"53",
          9459 => x"00",
          9460 => x"41",
          9461 => x"65",
          9462 => x"73",
          9463 => x"20",
          9464 => x"43",
          9465 => x"52",
          9466 => x"74",
          9467 => x"63",
          9468 => x"20",
          9469 => x"72",
          9470 => x"20",
          9471 => x"30",
          9472 => x"00",
          9473 => x"20",
          9474 => x"43",
          9475 => x"4d",
          9476 => x"72",
          9477 => x"74",
          9478 => x"20",
          9479 => x"72",
          9480 => x"20",
          9481 => x"30",
          9482 => x"00",
          9483 => x"20",
          9484 => x"53",
          9485 => x"6b",
          9486 => x"61",
          9487 => x"41",
          9488 => x"65",
          9489 => x"20",
          9490 => x"20",
          9491 => x"30",
          9492 => x"00",
          9493 => x"4d",
          9494 => x"3a",
          9495 => x"20",
          9496 => x"5a",
          9497 => x"49",
          9498 => x"20",
          9499 => x"20",
          9500 => x"20",
          9501 => x"20",
          9502 => x"20",
          9503 => x"30",
          9504 => x"00",
          9505 => x"20",
          9506 => x"53",
          9507 => x"65",
          9508 => x"6c",
          9509 => x"20",
          9510 => x"71",
          9511 => x"20",
          9512 => x"20",
          9513 => x"64",
          9514 => x"34",
          9515 => x"7a",
          9516 => x"20",
          9517 => x"53",
          9518 => x"4d",
          9519 => x"6f",
          9520 => x"46",
          9521 => x"20",
          9522 => x"20",
          9523 => x"20",
          9524 => x"64",
          9525 => x"34",
          9526 => x"7a",
          9527 => x"20",
          9528 => x"57",
          9529 => x"62",
          9530 => x"20",
          9531 => x"41",
          9532 => x"6c",
          9533 => x"20",
          9534 => x"71",
          9535 => x"64",
          9536 => x"34",
          9537 => x"7a",
          9538 => x"53",
          9539 => x"6c",
          9540 => x"4d",
          9541 => x"75",
          9542 => x"46",
          9543 => x"00",
          9544 => x"45",
          9545 => x"45",
          9546 => x"69",
          9547 => x"55",
          9548 => x"6f",
          9549 => x"00",
          9550 => x"01",
          9551 => x"00",
          9552 => x"00",
          9553 => x"01",
          9554 => x"00",
          9555 => x"00",
          9556 => x"01",
          9557 => x"00",
          9558 => x"00",
          9559 => x"01",
          9560 => x"00",
          9561 => x"00",
          9562 => x"01",
          9563 => x"00",
          9564 => x"00",
          9565 => x"01",
          9566 => x"00",
          9567 => x"00",
          9568 => x"01",
          9569 => x"00",
          9570 => x"00",
          9571 => x"01",
          9572 => x"00",
          9573 => x"00",
          9574 => x"01",
          9575 => x"00",
          9576 => x"00",
          9577 => x"01",
          9578 => x"00",
          9579 => x"00",
          9580 => x"01",
          9581 => x"00",
          9582 => x"00",
          9583 => x"04",
          9584 => x"00",
          9585 => x"00",
          9586 => x"04",
          9587 => x"00",
          9588 => x"00",
          9589 => x"04",
          9590 => x"00",
          9591 => x"00",
          9592 => x"03",
          9593 => x"00",
          9594 => x"00",
          9595 => x"04",
          9596 => x"00",
          9597 => x"00",
          9598 => x"04",
          9599 => x"00",
          9600 => x"00",
          9601 => x"04",
          9602 => x"00",
          9603 => x"00",
          9604 => x"03",
          9605 => x"00",
          9606 => x"00",
          9607 => x"03",
          9608 => x"00",
          9609 => x"00",
          9610 => x"03",
          9611 => x"00",
          9612 => x"00",
          9613 => x"03",
          9614 => x"00",
          9615 => x"1b",
          9616 => x"1b",
          9617 => x"1b",
          9618 => x"1b",
          9619 => x"1b",
          9620 => x"1b",
          9621 => x"1b",
          9622 => x"1b",
          9623 => x"1b",
          9624 => x"1b",
          9625 => x"1b",
          9626 => x"10",
          9627 => x"0e",
          9628 => x"0d",
          9629 => x"0b",
          9630 => x"08",
          9631 => x"06",
          9632 => x"05",
          9633 => x"04",
          9634 => x"03",
          9635 => x"02",
          9636 => x"01",
          9637 => x"68",
          9638 => x"6f",
          9639 => x"68",
          9640 => x"00",
          9641 => x"21",
          9642 => x"25",
          9643 => x"20",
          9644 => x"0a",
          9645 => x"46",
          9646 => x"65",
          9647 => x"6f",
          9648 => x"73",
          9649 => x"74",
          9650 => x"68",
          9651 => x"6f",
          9652 => x"66",
          9653 => x"20",
          9654 => x"45",
          9655 => x"0a",
          9656 => x"43",
          9657 => x"6f",
          9658 => x"70",
          9659 => x"63",
          9660 => x"74",
          9661 => x"69",
          9662 => x"72",
          9663 => x"69",
          9664 => x"20",
          9665 => x"61",
          9666 => x"6e",
          9667 => x"53",
          9668 => x"22",
          9669 => x"3a",
          9670 => x"3e",
          9671 => x"7c",
          9672 => x"46",
          9673 => x"46",
          9674 => x"32",
          9675 => x"eb",
          9676 => x"53",
          9677 => x"35",
          9678 => x"4e",
          9679 => x"41",
          9680 => x"20",
          9681 => x"41",
          9682 => x"20",
          9683 => x"4e",
          9684 => x"41",
          9685 => x"20",
          9686 => x"41",
          9687 => x"20",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"80",
          9693 => x"8e",
          9694 => x"45",
          9695 => x"49",
          9696 => x"90",
          9697 => x"99",
          9698 => x"59",
          9699 => x"9c",
          9700 => x"41",
          9701 => x"a5",
          9702 => x"a8",
          9703 => x"ac",
          9704 => x"b0",
          9705 => x"b4",
          9706 => x"b8",
          9707 => x"bc",
          9708 => x"c0",
          9709 => x"c4",
          9710 => x"c8",
          9711 => x"cc",
          9712 => x"d0",
          9713 => x"d4",
          9714 => x"d8",
          9715 => x"dc",
          9716 => x"e0",
          9717 => x"e4",
          9718 => x"e8",
          9719 => x"ec",
          9720 => x"f0",
          9721 => x"f4",
          9722 => x"f8",
          9723 => x"fc",
          9724 => x"2b",
          9725 => x"3d",
          9726 => x"5c",
          9727 => x"3c",
          9728 => x"7f",
          9729 => x"00",
          9730 => x"00",
          9731 => x"01",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"01",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"01",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"01",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"01",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"01",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"01",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"01",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"01",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"01",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"01",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"01",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"01",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"01",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"01",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"01",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"01",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"01",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"01",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"01",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"01",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"01",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"01",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"01",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"01",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"01",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"01",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"00",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"00",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"01",
          9852 => x"01",
          9853 => x"00",
          9854 => x"00",
          9855 => x"00",
          9856 => x"00",
          9857 => x"05",
          9858 => x"05",
          9859 => x"05",
          9860 => x"00",
          9861 => x"01",
          9862 => x"01",
          9863 => x"01",
          9864 => x"01",
          9865 => x"00",
          9866 => x"00",
          9867 => x"00",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"00",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"00",
          9890 => x"01",
          9891 => x"00",
          9892 => x"01",
          9893 => x"00",
          9894 => x"02",
          9895 => x"00",
          9896 => x"00",
          9897 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
