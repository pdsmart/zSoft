-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"93",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"d3",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"dc",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"94",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"95",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"d4",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"81",
           391 => x"83",
           392 => x"81",
           393 => x"b5",
           394 => x"f8",
           395 => x"80",
           396 => x"f8",
           397 => x"e4",
           398 => x"d4",
           399 => x"90",
           400 => x"d4",
           401 => x"2d",
           402 => x"08",
           403 => x"04",
           404 => x"0c",
           405 => x"81",
           406 => x"83",
           407 => x"81",
           408 => x"b6",
           409 => x"f8",
           410 => x"80",
           411 => x"f8",
           412 => x"bd",
           413 => x"d4",
           414 => x"90",
           415 => x"d4",
           416 => x"2d",
           417 => x"08",
           418 => x"04",
           419 => x"0c",
           420 => x"81",
           421 => x"83",
           422 => x"81",
           423 => x"b6",
           424 => x"f8",
           425 => x"80",
           426 => x"f8",
           427 => x"de",
           428 => x"d4",
           429 => x"90",
           430 => x"d4",
           431 => x"2d",
           432 => x"08",
           433 => x"04",
           434 => x"0c",
           435 => x"81",
           436 => x"83",
           437 => x"81",
           438 => x"a6",
           439 => x"f8",
           440 => x"80",
           441 => x"f8",
           442 => x"f9",
           443 => x"d4",
           444 => x"90",
           445 => x"d4",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"81",
           451 => x"83",
           452 => x"81",
           453 => x"81",
           454 => x"81",
           455 => x"83",
           456 => x"81",
           457 => x"81",
           458 => x"81",
           459 => x"83",
           460 => x"81",
           461 => x"81",
           462 => x"81",
           463 => x"83",
           464 => x"81",
           465 => x"81",
           466 => x"81",
           467 => x"83",
           468 => x"81",
           469 => x"81",
           470 => x"81",
           471 => x"83",
           472 => x"81",
           473 => x"81",
           474 => x"81",
           475 => x"83",
           476 => x"81",
           477 => x"81",
           478 => x"81",
           479 => x"83",
           480 => x"81",
           481 => x"81",
           482 => x"81",
           483 => x"83",
           484 => x"81",
           485 => x"81",
           486 => x"81",
           487 => x"83",
           488 => x"81",
           489 => x"81",
           490 => x"81",
           491 => x"83",
           492 => x"81",
           493 => x"81",
           494 => x"81",
           495 => x"83",
           496 => x"81",
           497 => x"81",
           498 => x"81",
           499 => x"83",
           500 => x"81",
           501 => x"81",
           502 => x"81",
           503 => x"83",
           504 => x"81",
           505 => x"81",
           506 => x"81",
           507 => x"83",
           508 => x"81",
           509 => x"81",
           510 => x"81",
           511 => x"83",
           512 => x"81",
           513 => x"81",
           514 => x"81",
           515 => x"83",
           516 => x"81",
           517 => x"81",
           518 => x"81",
           519 => x"83",
           520 => x"81",
           521 => x"81",
           522 => x"81",
           523 => x"83",
           524 => x"81",
           525 => x"81",
           526 => x"81",
           527 => x"83",
           528 => x"81",
           529 => x"81",
           530 => x"81",
           531 => x"83",
           532 => x"81",
           533 => x"81",
           534 => x"81",
           535 => x"83",
           536 => x"81",
           537 => x"81",
           538 => x"81",
           539 => x"83",
           540 => x"81",
           541 => x"81",
           542 => x"81",
           543 => x"83",
           544 => x"81",
           545 => x"81",
           546 => x"81",
           547 => x"83",
           548 => x"81",
           549 => x"81",
           550 => x"81",
           551 => x"83",
           552 => x"81",
           553 => x"81",
           554 => x"81",
           555 => x"83",
           556 => x"81",
           557 => x"81",
           558 => x"81",
           559 => x"83",
           560 => x"81",
           561 => x"80",
           562 => x"81",
           563 => x"83",
           564 => x"81",
           565 => x"80",
           566 => x"81",
           567 => x"83",
           568 => x"81",
           569 => x"80",
           570 => x"81",
           571 => x"83",
           572 => x"81",
           573 => x"9f",
           574 => x"f8",
           575 => x"80",
           576 => x"f8",
           577 => x"84",
           578 => x"d4",
           579 => x"90",
           580 => x"d4",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"00",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"53",
           597 => x"00",
           598 => x"06",
           599 => x"09",
           600 => x"05",
           601 => x"2b",
           602 => x"06",
           603 => x"04",
           604 => x"72",
           605 => x"05",
           606 => x"05",
           607 => x"72",
           608 => x"53",
           609 => x"51",
           610 => x"04",
           611 => x"70",
           612 => x"27",
           613 => x"71",
           614 => x"53",
           615 => x"0b",
           616 => x"8c",
           617 => x"da",
           618 => x"81",
           619 => x"02",
           620 => x"0c",
           621 => x"80",
           622 => x"d4",
           623 => x"08",
           624 => x"d4",
           625 => x"08",
           626 => x"3f",
           627 => x"08",
           628 => x"c8",
           629 => x"3d",
           630 => x"d4",
           631 => x"f8",
           632 => x"81",
           633 => x"fd",
           634 => x"53",
           635 => x"08",
           636 => x"52",
           637 => x"08",
           638 => x"51",
           639 => x"81",
           640 => x"70",
           641 => x"0c",
           642 => x"0d",
           643 => x"0c",
           644 => x"d4",
           645 => x"f8",
           646 => x"3d",
           647 => x"81",
           648 => x"fc",
           649 => x"f8",
           650 => x"05",
           651 => x"b9",
           652 => x"d4",
           653 => x"08",
           654 => x"d4",
           655 => x"0c",
           656 => x"f8",
           657 => x"05",
           658 => x"d4",
           659 => x"08",
           660 => x"0b",
           661 => x"08",
           662 => x"81",
           663 => x"f4",
           664 => x"f8",
           665 => x"05",
           666 => x"d4",
           667 => x"08",
           668 => x"38",
           669 => x"08",
           670 => x"30",
           671 => x"08",
           672 => x"80",
           673 => x"d4",
           674 => x"0c",
           675 => x"08",
           676 => x"8a",
           677 => x"81",
           678 => x"f0",
           679 => x"f8",
           680 => x"05",
           681 => x"d4",
           682 => x"0c",
           683 => x"f8",
           684 => x"05",
           685 => x"f8",
           686 => x"05",
           687 => x"df",
           688 => x"c8",
           689 => x"f8",
           690 => x"05",
           691 => x"f8",
           692 => x"05",
           693 => x"90",
           694 => x"d4",
           695 => x"08",
           696 => x"d4",
           697 => x"0c",
           698 => x"08",
           699 => x"70",
           700 => x"0c",
           701 => x"0d",
           702 => x"0c",
           703 => x"d4",
           704 => x"f8",
           705 => x"3d",
           706 => x"81",
           707 => x"fc",
           708 => x"f8",
           709 => x"05",
           710 => x"99",
           711 => x"d4",
           712 => x"08",
           713 => x"d4",
           714 => x"0c",
           715 => x"f8",
           716 => x"05",
           717 => x"d4",
           718 => x"08",
           719 => x"38",
           720 => x"08",
           721 => x"30",
           722 => x"08",
           723 => x"81",
           724 => x"d4",
           725 => x"08",
           726 => x"d4",
           727 => x"08",
           728 => x"81",
           729 => x"70",
           730 => x"08",
           731 => x"54",
           732 => x"08",
           733 => x"80",
           734 => x"81",
           735 => x"f8",
           736 => x"81",
           737 => x"f8",
           738 => x"f8",
           739 => x"05",
           740 => x"f8",
           741 => x"87",
           742 => x"f8",
           743 => x"81",
           744 => x"02",
           745 => x"0c",
           746 => x"81",
           747 => x"d4",
           748 => x"0c",
           749 => x"f8",
           750 => x"05",
           751 => x"d4",
           752 => x"08",
           753 => x"08",
           754 => x"27",
           755 => x"f8",
           756 => x"05",
           757 => x"ae",
           758 => x"81",
           759 => x"8c",
           760 => x"a2",
           761 => x"d4",
           762 => x"08",
           763 => x"d4",
           764 => x"0c",
           765 => x"08",
           766 => x"10",
           767 => x"08",
           768 => x"ff",
           769 => x"f8",
           770 => x"05",
           771 => x"80",
           772 => x"f8",
           773 => x"05",
           774 => x"d4",
           775 => x"08",
           776 => x"81",
           777 => x"88",
           778 => x"f8",
           779 => x"05",
           780 => x"f8",
           781 => x"05",
           782 => x"d4",
           783 => x"08",
           784 => x"08",
           785 => x"07",
           786 => x"08",
           787 => x"81",
           788 => x"fc",
           789 => x"2a",
           790 => x"08",
           791 => x"81",
           792 => x"8c",
           793 => x"2a",
           794 => x"08",
           795 => x"ff",
           796 => x"f8",
           797 => x"05",
           798 => x"93",
           799 => x"d4",
           800 => x"08",
           801 => x"d4",
           802 => x"0c",
           803 => x"81",
           804 => x"f8",
           805 => x"81",
           806 => x"f4",
           807 => x"81",
           808 => x"f4",
           809 => x"f8",
           810 => x"3d",
           811 => x"d4",
           812 => x"3d",
           813 => x"79",
           814 => x"55",
           815 => x"27",
           816 => x"75",
           817 => x"51",
           818 => x"a9",
           819 => x"52",
           820 => x"98",
           821 => x"81",
           822 => x"74",
           823 => x"56",
           824 => x"52",
           825 => x"09",
           826 => x"38",
           827 => x"c8",
           828 => x"0d",
           829 => x"72",
           830 => x"54",
           831 => x"84",
           832 => x"72",
           833 => x"54",
           834 => x"84",
           835 => x"72",
           836 => x"54",
           837 => x"84",
           838 => x"72",
           839 => x"54",
           840 => x"84",
           841 => x"f0",
           842 => x"8f",
           843 => x"83",
           844 => x"38",
           845 => x"05",
           846 => x"70",
           847 => x"0c",
           848 => x"71",
           849 => x"38",
           850 => x"81",
           851 => x"0d",
           852 => x"02",
           853 => x"05",
           854 => x"53",
           855 => x"27",
           856 => x"83",
           857 => x"80",
           858 => x"ff",
           859 => x"ff",
           860 => x"73",
           861 => x"05",
           862 => x"12",
           863 => x"2e",
           864 => x"ef",
           865 => x"f8",
           866 => x"3d",
           867 => x"74",
           868 => x"07",
           869 => x"2b",
           870 => x"51",
           871 => x"a5",
           872 => x"70",
           873 => x"0c",
           874 => x"84",
           875 => x"72",
           876 => x"05",
           877 => x"71",
           878 => x"53",
           879 => x"52",
           880 => x"dd",
           881 => x"27",
           882 => x"71",
           883 => x"53",
           884 => x"52",
           885 => x"f2",
           886 => x"ff",
           887 => x"3d",
           888 => x"79",
           889 => x"83",
           890 => x"54",
           891 => x"c3",
           892 => x"08",
           893 => x"f7",
           894 => x"13",
           895 => x"84",
           896 => x"06",
           897 => x"53",
           898 => x"38",
           899 => x"74",
           900 => x"56",
           901 => x"70",
           902 => x"fb",
           903 => x"06",
           904 => x"82",
           905 => x"51",
           906 => x"54",
           907 => x"dc",
           908 => x"71",
           909 => x"53",
           910 => x"73",
           911 => x"55",
           912 => x"38",
           913 => x"c8",
           914 => x"0d",
           915 => x"0d",
           916 => x"83",
           917 => x"52",
           918 => x"71",
           919 => x"09",
           920 => x"ff",
           921 => x"f8",
           922 => x"80",
           923 => x"52",
           924 => x"38",
           925 => x"08",
           926 => x"fb",
           927 => x"06",
           928 => x"82",
           929 => x"51",
           930 => x"70",
           931 => x"38",
           932 => x"33",
           933 => x"2e",
           934 => x"12",
           935 => x"52",
           936 => x"71",
           937 => x"f8",
           938 => x"3d",
           939 => x"3d",
           940 => x"7c",
           941 => x"55",
           942 => x"2e",
           943 => x"71",
           944 => x"06",
           945 => x"2e",
           946 => x"ff",
           947 => x"ff",
           948 => x"71",
           949 => x"56",
           950 => x"2e",
           951 => x"a9",
           952 => x"2e",
           953 => x"70",
           954 => x"51",
           955 => x"80",
           956 => x"12",
           957 => x"15",
           958 => x"72",
           959 => x"81",
           960 => x"71",
           961 => x"56",
           962 => x"ff",
           963 => x"ff",
           964 => x"31",
           965 => x"70",
           966 => x"0c",
           967 => x"04",
           968 => x"55",
           969 => x"88",
           970 => x"74",
           971 => x"38",
           972 => x"52",
           973 => x"fc",
           974 => x"80",
           975 => x"74",
           976 => x"f7",
           977 => x"12",
           978 => x"84",
           979 => x"06",
           980 => x"70",
           981 => x"15",
           982 => x"55",
           983 => x"d0",
           984 => x"76",
           985 => x"38",
           986 => x"52",
           987 => x"80",
           988 => x"c8",
           989 => x"0d",
           990 => x"0d",
           991 => x"53",
           992 => x"52",
           993 => x"81",
           994 => x"81",
           995 => x"07",
           996 => x"52",
           997 => x"e8",
           998 => x"f8",
           999 => x"3d",
          1000 => x"3d",
          1001 => x"08",
          1002 => x"56",
          1003 => x"80",
          1004 => x"33",
          1005 => x"2e",
          1006 => x"86",
          1007 => x"52",
          1008 => x"53",
          1009 => x"13",
          1010 => x"33",
          1011 => x"06",
          1012 => x"70",
          1013 => x"38",
          1014 => x"80",
          1015 => x"74",
          1016 => x"81",
          1017 => x"70",
          1018 => x"81",
          1019 => x"80",
          1020 => x"05",
          1021 => x"76",
          1022 => x"70",
          1023 => x"0c",
          1024 => x"04",
          1025 => x"76",
          1026 => x"80",
          1027 => x"86",
          1028 => x"52",
          1029 => x"97",
          1030 => x"c8",
          1031 => x"80",
          1032 => x"74",
          1033 => x"f8",
          1034 => x"3d",
          1035 => x"3d",
          1036 => x"11",
          1037 => x"52",
          1038 => x"70",
          1039 => x"98",
          1040 => x"33",
          1041 => x"82",
          1042 => x"26",
          1043 => x"84",
          1044 => x"83",
          1045 => x"26",
          1046 => x"85",
          1047 => x"84",
          1048 => x"26",
          1049 => x"86",
          1050 => x"85",
          1051 => x"26",
          1052 => x"88",
          1053 => x"86",
          1054 => x"e7",
          1055 => x"38",
          1056 => x"54",
          1057 => x"87",
          1058 => x"cc",
          1059 => x"87",
          1060 => x"0c",
          1061 => x"c0",
          1062 => x"82",
          1063 => x"c0",
          1064 => x"83",
          1065 => x"c0",
          1066 => x"84",
          1067 => x"c0",
          1068 => x"85",
          1069 => x"c0",
          1070 => x"86",
          1071 => x"c0",
          1072 => x"74",
          1073 => x"a4",
          1074 => x"c0",
          1075 => x"80",
          1076 => x"98",
          1077 => x"52",
          1078 => x"c8",
          1079 => x"0d",
          1080 => x"0d",
          1081 => x"c0",
          1082 => x"81",
          1083 => x"c0",
          1084 => x"5e",
          1085 => x"87",
          1086 => x"08",
          1087 => x"1c",
          1088 => x"98",
          1089 => x"79",
          1090 => x"87",
          1091 => x"08",
          1092 => x"1c",
          1093 => x"98",
          1094 => x"79",
          1095 => x"87",
          1096 => x"08",
          1097 => x"1c",
          1098 => x"98",
          1099 => x"7b",
          1100 => x"87",
          1101 => x"08",
          1102 => x"1c",
          1103 => x"0c",
          1104 => x"ff",
          1105 => x"83",
          1106 => x"58",
          1107 => x"57",
          1108 => x"56",
          1109 => x"55",
          1110 => x"54",
          1111 => x"53",
          1112 => x"ff",
          1113 => x"dd",
          1114 => x"dc",
          1115 => x"0d",
          1116 => x"0d",
          1117 => x"33",
          1118 => x"9f",
          1119 => x"52",
          1120 => x"81",
          1121 => x"83",
          1122 => x"fb",
          1123 => x"0b",
          1124 => x"c0",
          1125 => x"ff",
          1126 => x"56",
          1127 => x"84",
          1128 => x"2e",
          1129 => x"c0",
          1130 => x"70",
          1131 => x"2a",
          1132 => x"53",
          1133 => x"80",
          1134 => x"71",
          1135 => x"81",
          1136 => x"70",
          1137 => x"81",
          1138 => x"06",
          1139 => x"80",
          1140 => x"71",
          1141 => x"81",
          1142 => x"70",
          1143 => x"73",
          1144 => x"51",
          1145 => x"80",
          1146 => x"2e",
          1147 => x"c0",
          1148 => x"75",
          1149 => x"81",
          1150 => x"87",
          1151 => x"fb",
          1152 => x"9f",
          1153 => x"0b",
          1154 => x"33",
          1155 => x"06",
          1156 => x"87",
          1157 => x"51",
          1158 => x"86",
          1159 => x"94",
          1160 => x"08",
          1161 => x"70",
          1162 => x"54",
          1163 => x"2e",
          1164 => x"91",
          1165 => x"06",
          1166 => x"d7",
          1167 => x"32",
          1168 => x"51",
          1169 => x"2e",
          1170 => x"93",
          1171 => x"06",
          1172 => x"ff",
          1173 => x"81",
          1174 => x"87",
          1175 => x"52",
          1176 => x"86",
          1177 => x"94",
          1178 => x"72",
          1179 => x"0d",
          1180 => x"0d",
          1181 => x"74",
          1182 => x"ff",
          1183 => x"57",
          1184 => x"80",
          1185 => x"81",
          1186 => x"15",
          1187 => x"f3",
          1188 => x"81",
          1189 => x"57",
          1190 => x"c0",
          1191 => x"75",
          1192 => x"38",
          1193 => x"94",
          1194 => x"70",
          1195 => x"81",
          1196 => x"52",
          1197 => x"8c",
          1198 => x"2a",
          1199 => x"51",
          1200 => x"38",
          1201 => x"70",
          1202 => x"51",
          1203 => x"8d",
          1204 => x"2a",
          1205 => x"51",
          1206 => x"be",
          1207 => x"ff",
          1208 => x"c0",
          1209 => x"70",
          1210 => x"38",
          1211 => x"90",
          1212 => x"0c",
          1213 => x"33",
          1214 => x"06",
          1215 => x"70",
          1216 => x"76",
          1217 => x"0c",
          1218 => x"04",
          1219 => x"0b",
          1220 => x"c0",
          1221 => x"ff",
          1222 => x"87",
          1223 => x"51",
          1224 => x"86",
          1225 => x"94",
          1226 => x"08",
          1227 => x"70",
          1228 => x"51",
          1229 => x"2e",
          1230 => x"81",
          1231 => x"87",
          1232 => x"52",
          1233 => x"86",
          1234 => x"94",
          1235 => x"08",
          1236 => x"06",
          1237 => x"0c",
          1238 => x"0d",
          1239 => x"0d",
          1240 => x"f3",
          1241 => x"81",
          1242 => x"53",
          1243 => x"84",
          1244 => x"2e",
          1245 => x"c0",
          1246 => x"71",
          1247 => x"2a",
          1248 => x"51",
          1249 => x"52",
          1250 => x"a0",
          1251 => x"ff",
          1252 => x"c0",
          1253 => x"70",
          1254 => x"38",
          1255 => x"90",
          1256 => x"70",
          1257 => x"98",
          1258 => x"51",
          1259 => x"c8",
          1260 => x"0d",
          1261 => x"0d",
          1262 => x"80",
          1263 => x"2a",
          1264 => x"51",
          1265 => x"84",
          1266 => x"c0",
          1267 => x"81",
          1268 => x"87",
          1269 => x"08",
          1270 => x"0c",
          1271 => x"94",
          1272 => x"cc",
          1273 => x"9e",
          1274 => x"f3",
          1275 => x"c0",
          1276 => x"81",
          1277 => x"87",
          1278 => x"08",
          1279 => x"0c",
          1280 => x"ac",
          1281 => x"dc",
          1282 => x"9e",
          1283 => x"f3",
          1284 => x"c0",
          1285 => x"81",
          1286 => x"87",
          1287 => x"08",
          1288 => x"0c",
          1289 => x"bc",
          1290 => x"ec",
          1291 => x"9e",
          1292 => x"f3",
          1293 => x"c0",
          1294 => x"81",
          1295 => x"87",
          1296 => x"08",
          1297 => x"f3",
          1298 => x"c0",
          1299 => x"81",
          1300 => x"87",
          1301 => x"08",
          1302 => x"0c",
          1303 => x"8c",
          1304 => x"84",
          1305 => x"81",
          1306 => x"80",
          1307 => x"9e",
          1308 => x"84",
          1309 => x"51",
          1310 => x"80",
          1311 => x"81",
          1312 => x"f4",
          1313 => x"0b",
          1314 => x"90",
          1315 => x"80",
          1316 => x"52",
          1317 => x"2e",
          1318 => x"52",
          1319 => x"8a",
          1320 => x"87",
          1321 => x"08",
          1322 => x"0a",
          1323 => x"52",
          1324 => x"83",
          1325 => x"71",
          1326 => x"34",
          1327 => x"c0",
          1328 => x"70",
          1329 => x"06",
          1330 => x"70",
          1331 => x"38",
          1332 => x"81",
          1333 => x"80",
          1334 => x"9e",
          1335 => x"a0",
          1336 => x"51",
          1337 => x"80",
          1338 => x"81",
          1339 => x"f4",
          1340 => x"0b",
          1341 => x"90",
          1342 => x"80",
          1343 => x"52",
          1344 => x"2e",
          1345 => x"52",
          1346 => x"8e",
          1347 => x"87",
          1348 => x"08",
          1349 => x"80",
          1350 => x"52",
          1351 => x"83",
          1352 => x"71",
          1353 => x"34",
          1354 => x"c0",
          1355 => x"70",
          1356 => x"06",
          1357 => x"70",
          1358 => x"38",
          1359 => x"81",
          1360 => x"80",
          1361 => x"9e",
          1362 => x"81",
          1363 => x"51",
          1364 => x"80",
          1365 => x"81",
          1366 => x"f4",
          1367 => x"0b",
          1368 => x"90",
          1369 => x"c0",
          1370 => x"52",
          1371 => x"2e",
          1372 => x"52",
          1373 => x"92",
          1374 => x"87",
          1375 => x"08",
          1376 => x"06",
          1377 => x"70",
          1378 => x"38",
          1379 => x"81",
          1380 => x"87",
          1381 => x"08",
          1382 => x"06",
          1383 => x"51",
          1384 => x"81",
          1385 => x"80",
          1386 => x"9e",
          1387 => x"84",
          1388 => x"52",
          1389 => x"2e",
          1390 => x"52",
          1391 => x"95",
          1392 => x"9e",
          1393 => x"83",
          1394 => x"84",
          1395 => x"51",
          1396 => x"96",
          1397 => x"87",
          1398 => x"08",
          1399 => x"51",
          1400 => x"80",
          1401 => x"81",
          1402 => x"f4",
          1403 => x"c0",
          1404 => x"70",
          1405 => x"51",
          1406 => x"98",
          1407 => x"0d",
          1408 => x"0d",
          1409 => x"51",
          1410 => x"81",
          1411 => x"54",
          1412 => x"88",
          1413 => x"fc",
          1414 => x"3f",
          1415 => x"51",
          1416 => x"81",
          1417 => x"54",
          1418 => x"93",
          1419 => x"e4",
          1420 => x"e8",
          1421 => x"52",
          1422 => x"51",
          1423 => x"81",
          1424 => x"54",
          1425 => x"93",
          1426 => x"dc",
          1427 => x"e0",
          1428 => x"52",
          1429 => x"51",
          1430 => x"81",
          1431 => x"54",
          1432 => x"93",
          1433 => x"c4",
          1434 => x"c8",
          1435 => x"52",
          1436 => x"51",
          1437 => x"81",
          1438 => x"54",
          1439 => x"93",
          1440 => x"cc",
          1441 => x"d0",
          1442 => x"52",
          1443 => x"51",
          1444 => x"81",
          1445 => x"54",
          1446 => x"93",
          1447 => x"d4",
          1448 => x"d8",
          1449 => x"52",
          1450 => x"51",
          1451 => x"81",
          1452 => x"54",
          1453 => x"8d",
          1454 => x"94",
          1455 => x"df",
          1456 => x"84",
          1457 => x"97",
          1458 => x"80",
          1459 => x"81",
          1460 => x"52",
          1461 => x"51",
          1462 => x"81",
          1463 => x"54",
          1464 => x"8d",
          1465 => x"96",
          1466 => x"df",
          1467 => x"d8",
          1468 => x"89",
          1469 => x"80",
          1470 => x"81",
          1471 => x"87",
          1472 => x"f4",
          1473 => x"73",
          1474 => x"38",
          1475 => x"51",
          1476 => x"81",
          1477 => x"54",
          1478 => x"88",
          1479 => x"b4",
          1480 => x"3f",
          1481 => x"33",
          1482 => x"2e",
          1483 => x"e0",
          1484 => x"b0",
          1485 => x"92",
          1486 => x"80",
          1487 => x"81",
          1488 => x"87",
          1489 => x"e0",
          1490 => x"98",
          1491 => x"ec",
          1492 => x"e0",
          1493 => x"f0",
          1494 => x"f0",
          1495 => x"e1",
          1496 => x"e4",
          1497 => x"f4",
          1498 => x"e1",
          1499 => x"d8",
          1500 => x"dc",
          1501 => x"3f",
          1502 => x"22",
          1503 => x"e4",
          1504 => x"3f",
          1505 => x"08",
          1506 => x"c0",
          1507 => x"e4",
          1508 => x"f8",
          1509 => x"84",
          1510 => x"71",
          1511 => x"81",
          1512 => x"52",
          1513 => x"51",
          1514 => x"81",
          1515 => x"54",
          1516 => x"a8",
          1517 => x"80",
          1518 => x"84",
          1519 => x"51",
          1520 => x"81",
          1521 => x"bd",
          1522 => x"76",
          1523 => x"54",
          1524 => x"08",
          1525 => x"b8",
          1526 => x"3f",
          1527 => x"33",
          1528 => x"2e",
          1529 => x"f4",
          1530 => x"bd",
          1531 => x"75",
          1532 => x"3f",
          1533 => x"08",
          1534 => x"29",
          1535 => x"54",
          1536 => x"c8",
          1537 => x"e2",
          1538 => x"bc",
          1539 => x"90",
          1540 => x"3f",
          1541 => x"04",
          1542 => x"02",
          1543 => x"ff",
          1544 => x"84",
          1545 => x"71",
          1546 => x"dc",
          1547 => x"71",
          1548 => x"e3",
          1549 => x"39",
          1550 => x"51",
          1551 => x"e3",
          1552 => x"39",
          1553 => x"51",
          1554 => x"e3",
          1555 => x"39",
          1556 => x"51",
          1557 => x"84",
          1558 => x"71",
          1559 => x"04",
          1560 => x"c0",
          1561 => x"04",
          1562 => x"08",
          1563 => x"84",
          1564 => x"3d",
          1565 => x"d8",
          1566 => x"82",
          1567 => x"81",
          1568 => x"81",
          1569 => x"75",
          1570 => x"ff",
          1571 => x"b7",
          1572 => x"38",
          1573 => x"d8",
          1574 => x"72",
          1575 => x"0c",
          1576 => x"04",
          1577 => x"79",
          1578 => x"08",
          1579 => x"14",
          1580 => x"08",
          1581 => x"5a",
          1582 => x"57",
          1583 => x"26",
          1584 => x"13",
          1585 => x"53",
          1586 => x"0c",
          1587 => x"84",
          1588 => x"73",
          1589 => x"14",
          1590 => x"12",
          1591 => x"12",
          1592 => x"13",
          1593 => x"14",
          1594 => x"12",
          1595 => x"12",
          1596 => x"15",
          1597 => x"16",
          1598 => x"80",
          1599 => x"90",
          1600 => x"94",
          1601 => x"81",
          1602 => x"89",
          1603 => x"fc",
          1604 => x"8c",
          1605 => x"12",
          1606 => x"53",
          1607 => x"2e",
          1608 => x"a3",
          1609 => x"08",
          1610 => x"55",
          1611 => x"09",
          1612 => x"38",
          1613 => x"15",
          1614 => x"73",
          1615 => x"71",
          1616 => x"71",
          1617 => x"81",
          1618 => x"f4",
          1619 => x"14",
          1620 => x"a0",
          1621 => x"0c",
          1622 => x"b0",
          1623 => x"08",
          1624 => x"0c",
          1625 => x"81",
          1626 => x"06",
          1627 => x"13",
          1628 => x"52",
          1629 => x"2e",
          1630 => x"a4",
          1631 => x"08",
          1632 => x"0c",
          1633 => x"90",
          1634 => x"90",
          1635 => x"94",
          1636 => x"14",
          1637 => x"08",
          1638 => x"0c",
          1639 => x"0c",
          1640 => x"c8",
          1641 => x"0d",
          1642 => x"0d",
          1643 => x"57",
          1644 => x"81",
          1645 => x"17",
          1646 => x"f4",
          1647 => x"57",
          1648 => x"2e",
          1649 => x"16",
          1650 => x"80",
          1651 => x"16",
          1652 => x"39",
          1653 => x"17",
          1654 => x"06",
          1655 => x"fd",
          1656 => x"f8",
          1657 => x"f8",
          1658 => x"70",
          1659 => x"08",
          1660 => x"81",
          1661 => x"09",
          1662 => x"72",
          1663 => x"73",
          1664 => x"58",
          1665 => x"80",
          1666 => x"2e",
          1667 => x"80",
          1668 => x"39",
          1669 => x"51",
          1670 => x"81",
          1671 => x"c8",
          1672 => x"81",
          1673 => x"84",
          1674 => x"f4",
          1675 => x"72",
          1676 => x"8c",
          1677 => x"26",
          1678 => x"13",
          1679 => x"39",
          1680 => x"88",
          1681 => x"8c",
          1682 => x"88",
          1683 => x"16",
          1684 => x"12",
          1685 => x"51",
          1686 => x"76",
          1687 => x"c8",
          1688 => x"c0",
          1689 => x"c8",
          1690 => x"81",
          1691 => x"89",
          1692 => x"ff",
          1693 => x"52",
          1694 => x"87",
          1695 => x"51",
          1696 => x"83",
          1697 => x"fe",
          1698 => x"93",
          1699 => x"72",
          1700 => x"81",
          1701 => x"8d",
          1702 => x"81",
          1703 => x"52",
          1704 => x"90",
          1705 => x"34",
          1706 => x"08",
          1707 => x"f8",
          1708 => x"39",
          1709 => x"08",
          1710 => x"2e",
          1711 => x"51",
          1712 => x"3d",
          1713 => x"3d",
          1714 => x"05",
          1715 => x"dc",
          1716 => x"f8",
          1717 => x"51",
          1718 => x"72",
          1719 => x"0c",
          1720 => x"04",
          1721 => x"75",
          1722 => x"70",
          1723 => x"53",
          1724 => x"2e",
          1725 => x"81",
          1726 => x"81",
          1727 => x"87",
          1728 => x"85",
          1729 => x"fc",
          1730 => x"81",
          1731 => x"78",
          1732 => x"0c",
          1733 => x"33",
          1734 => x"06",
          1735 => x"80",
          1736 => x"72",
          1737 => x"51",
          1738 => x"fe",
          1739 => x"39",
          1740 => x"dc",
          1741 => x"0d",
          1742 => x"0d",
          1743 => x"59",
          1744 => x"05",
          1745 => x"75",
          1746 => x"f8",
          1747 => x"2e",
          1748 => x"82",
          1749 => x"70",
          1750 => x"05",
          1751 => x"5b",
          1752 => x"2e",
          1753 => x"85",
          1754 => x"8b",
          1755 => x"2e",
          1756 => x"8a",
          1757 => x"78",
          1758 => x"5a",
          1759 => x"aa",
          1760 => x"06",
          1761 => x"84",
          1762 => x"7b",
          1763 => x"5d",
          1764 => x"59",
          1765 => x"d0",
          1766 => x"89",
          1767 => x"7a",
          1768 => x"10",
          1769 => x"d0",
          1770 => x"81",
          1771 => x"57",
          1772 => x"75",
          1773 => x"70",
          1774 => x"07",
          1775 => x"80",
          1776 => x"30",
          1777 => x"80",
          1778 => x"53",
          1779 => x"55",
          1780 => x"2e",
          1781 => x"84",
          1782 => x"81",
          1783 => x"57",
          1784 => x"2e",
          1785 => x"75",
          1786 => x"76",
          1787 => x"e0",
          1788 => x"ff",
          1789 => x"73",
          1790 => x"81",
          1791 => x"80",
          1792 => x"38",
          1793 => x"2e",
          1794 => x"73",
          1795 => x"8b",
          1796 => x"c2",
          1797 => x"38",
          1798 => x"73",
          1799 => x"81",
          1800 => x"8f",
          1801 => x"d5",
          1802 => x"38",
          1803 => x"24",
          1804 => x"80",
          1805 => x"38",
          1806 => x"73",
          1807 => x"80",
          1808 => x"ef",
          1809 => x"19",
          1810 => x"59",
          1811 => x"33",
          1812 => x"75",
          1813 => x"81",
          1814 => x"70",
          1815 => x"55",
          1816 => x"79",
          1817 => x"90",
          1818 => x"16",
          1819 => x"7b",
          1820 => x"a0",
          1821 => x"3f",
          1822 => x"53",
          1823 => x"e9",
          1824 => x"fc",
          1825 => x"81",
          1826 => x"72",
          1827 => x"b0",
          1828 => x"fb",
          1829 => x"39",
          1830 => x"83",
          1831 => x"59",
          1832 => x"82",
          1833 => x"88",
          1834 => x"8a",
          1835 => x"90",
          1836 => x"75",
          1837 => x"3f",
          1838 => x"79",
          1839 => x"81",
          1840 => x"72",
          1841 => x"38",
          1842 => x"59",
          1843 => x"84",
          1844 => x"58",
          1845 => x"80",
          1846 => x"30",
          1847 => x"80",
          1848 => x"55",
          1849 => x"25",
          1850 => x"80",
          1851 => x"74",
          1852 => x"07",
          1853 => x"0b",
          1854 => x"57",
          1855 => x"51",
          1856 => x"81",
          1857 => x"81",
          1858 => x"53",
          1859 => x"d9",
          1860 => x"f8",
          1861 => x"89",
          1862 => x"38",
          1863 => x"75",
          1864 => x"84",
          1865 => x"53",
          1866 => x"06",
          1867 => x"53",
          1868 => x"81",
          1869 => x"81",
          1870 => x"70",
          1871 => x"2a",
          1872 => x"76",
          1873 => x"38",
          1874 => x"38",
          1875 => x"70",
          1876 => x"53",
          1877 => x"8e",
          1878 => x"77",
          1879 => x"53",
          1880 => x"81",
          1881 => x"7a",
          1882 => x"55",
          1883 => x"83",
          1884 => x"79",
          1885 => x"81",
          1886 => x"72",
          1887 => x"17",
          1888 => x"27",
          1889 => x"51",
          1890 => x"75",
          1891 => x"72",
          1892 => x"81",
          1893 => x"7a",
          1894 => x"38",
          1895 => x"05",
          1896 => x"ff",
          1897 => x"70",
          1898 => x"57",
          1899 => x"76",
          1900 => x"81",
          1901 => x"72",
          1902 => x"84",
          1903 => x"f9",
          1904 => x"39",
          1905 => x"04",
          1906 => x"86",
          1907 => x"84",
          1908 => x"55",
          1909 => x"fa",
          1910 => x"3d",
          1911 => x"3d",
          1912 => x"f8",
          1913 => x"3d",
          1914 => x"75",
          1915 => x"3f",
          1916 => x"08",
          1917 => x"34",
          1918 => x"f8",
          1919 => x"3d",
          1920 => x"3d",
          1921 => x"dc",
          1922 => x"f8",
          1923 => x"3d",
          1924 => x"77",
          1925 => x"a1",
          1926 => x"f8",
          1927 => x"3d",
          1928 => x"3d",
          1929 => x"81",
          1930 => x"70",
          1931 => x"55",
          1932 => x"80",
          1933 => x"38",
          1934 => x"08",
          1935 => x"81",
          1936 => x"81",
          1937 => x"72",
          1938 => x"cb",
          1939 => x"2e",
          1940 => x"88",
          1941 => x"70",
          1942 => x"51",
          1943 => x"2e",
          1944 => x"80",
          1945 => x"ff",
          1946 => x"39",
          1947 => x"c8",
          1948 => x"52",
          1949 => x"c0",
          1950 => x"52",
          1951 => x"81",
          1952 => x"51",
          1953 => x"ff",
          1954 => x"15",
          1955 => x"34",
          1956 => x"f3",
          1957 => x"72",
          1958 => x"0c",
          1959 => x"04",
          1960 => x"81",
          1961 => x"75",
          1962 => x"0c",
          1963 => x"52",
          1964 => x"3f",
          1965 => x"e0",
          1966 => x"0d",
          1967 => x"0d",
          1968 => x"56",
          1969 => x"0c",
          1970 => x"70",
          1971 => x"73",
          1972 => x"81",
          1973 => x"81",
          1974 => x"ed",
          1975 => x"2e",
          1976 => x"8e",
          1977 => x"08",
          1978 => x"76",
          1979 => x"56",
          1980 => x"b0",
          1981 => x"06",
          1982 => x"75",
          1983 => x"76",
          1984 => x"70",
          1985 => x"73",
          1986 => x"8b",
          1987 => x"73",
          1988 => x"85",
          1989 => x"82",
          1990 => x"76",
          1991 => x"70",
          1992 => x"ac",
          1993 => x"a0",
          1994 => x"fa",
          1995 => x"53",
          1996 => x"57",
          1997 => x"98",
          1998 => x"39",
          1999 => x"80",
          2000 => x"26",
          2001 => x"86",
          2002 => x"80",
          2003 => x"57",
          2004 => x"74",
          2005 => x"38",
          2006 => x"27",
          2007 => x"14",
          2008 => x"06",
          2009 => x"14",
          2010 => x"06",
          2011 => x"74",
          2012 => x"f9",
          2013 => x"ff",
          2014 => x"89",
          2015 => x"38",
          2016 => x"c5",
          2017 => x"29",
          2018 => x"81",
          2019 => x"76",
          2020 => x"56",
          2021 => x"ba",
          2022 => x"2e",
          2023 => x"30",
          2024 => x"0c",
          2025 => x"81",
          2026 => x"8a",
          2027 => x"f8",
          2028 => x"7c",
          2029 => x"70",
          2030 => x"75",
          2031 => x"55",
          2032 => x"2e",
          2033 => x"87",
          2034 => x"76",
          2035 => x"73",
          2036 => x"81",
          2037 => x"81",
          2038 => x"77",
          2039 => x"70",
          2040 => x"58",
          2041 => x"09",
          2042 => x"c2",
          2043 => x"81",
          2044 => x"75",
          2045 => x"55",
          2046 => x"e2",
          2047 => x"90",
          2048 => x"f8",
          2049 => x"8f",
          2050 => x"81",
          2051 => x"75",
          2052 => x"55",
          2053 => x"81",
          2054 => x"27",
          2055 => x"d0",
          2056 => x"55",
          2057 => x"73",
          2058 => x"80",
          2059 => x"14",
          2060 => x"72",
          2061 => x"e0",
          2062 => x"80",
          2063 => x"39",
          2064 => x"55",
          2065 => x"80",
          2066 => x"e0",
          2067 => x"38",
          2068 => x"81",
          2069 => x"53",
          2070 => x"81",
          2071 => x"53",
          2072 => x"8e",
          2073 => x"70",
          2074 => x"55",
          2075 => x"27",
          2076 => x"77",
          2077 => x"74",
          2078 => x"76",
          2079 => x"77",
          2080 => x"70",
          2081 => x"55",
          2082 => x"77",
          2083 => x"38",
          2084 => x"74",
          2085 => x"55",
          2086 => x"c8",
          2087 => x"0d",
          2088 => x"0d",
          2089 => x"70",
          2090 => x"98",
          2091 => x"2c",
          2092 => x"70",
          2093 => x"53",
          2094 => x"51",
          2095 => x"e4",
          2096 => x"55",
          2097 => x"25",
          2098 => x"e4",
          2099 => x"12",
          2100 => x"97",
          2101 => x"33",
          2102 => x"70",
          2103 => x"81",
          2104 => x"81",
          2105 => x"f8",
          2106 => x"3d",
          2107 => x"3d",
          2108 => x"84",
          2109 => x"33",
          2110 => x"55",
          2111 => x"2e",
          2112 => x"51",
          2113 => x"a0",
          2114 => x"3f",
          2115 => x"f7",
          2116 => x"ff",
          2117 => x"73",
          2118 => x"ff",
          2119 => x"39",
          2120 => x"c0",
          2121 => x"34",
          2122 => x"04",
          2123 => x"7c",
          2124 => x"b7",
          2125 => x"88",
          2126 => x"33",
          2127 => x"33",
          2128 => x"81",
          2129 => x"70",
          2130 => x"59",
          2131 => x"74",
          2132 => x"38",
          2133 => x"9b",
          2134 => x"94",
          2135 => x"29",
          2136 => x"05",
          2137 => x"54",
          2138 => x"f0",
          2139 => x"f8",
          2140 => x"0c",
          2141 => x"33",
          2142 => x"81",
          2143 => x"70",
          2144 => x"5a",
          2145 => x"a6",
          2146 => x"78",
          2147 => x"d6",
          2148 => x"f5",
          2149 => x"05",
          2150 => x"f5",
          2151 => x"81",
          2152 => x"93",
          2153 => x"38",
          2154 => x"f5",
          2155 => x"80",
          2156 => x"81",
          2157 => x"56",
          2158 => x"ac",
          2159 => x"8c",
          2160 => x"a4",
          2161 => x"fc",
          2162 => x"53",
          2163 => x"51",
          2164 => x"3f",
          2165 => x"08",
          2166 => x"80",
          2167 => x"81",
          2168 => x"51",
          2169 => x"3f",
          2170 => x"04",
          2171 => x"81",
          2172 => x"81",
          2173 => x"51",
          2174 => x"3f",
          2175 => x"08",
          2176 => x"81",
          2177 => x"53",
          2178 => x"88",
          2179 => x"56",
          2180 => x"3f",
          2181 => x"08",
          2182 => x"38",
          2183 => x"ad",
          2184 => x"c8",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"81",
          2188 => x"ff",
          2189 => x"55",
          2190 => x"34",
          2191 => x"52",
          2192 => x"e3",
          2193 => x"f6",
          2194 => x"ff",
          2195 => x"06",
          2196 => x"a6",
          2197 => x"d9",
          2198 => x"3d",
          2199 => x"08",
          2200 => x"70",
          2201 => x"52",
          2202 => x"08",
          2203 => x"92",
          2204 => x"c8",
          2205 => x"38",
          2206 => x"f5",
          2207 => x"55",
          2208 => x"8b",
          2209 => x"56",
          2210 => x"3f",
          2211 => x"08",
          2212 => x"38",
          2213 => x"b5",
          2214 => x"c8",
          2215 => x"58",
          2216 => x"81",
          2217 => x"25",
          2218 => x"f8",
          2219 => x"05",
          2220 => x"55",
          2221 => x"74",
          2222 => x"70",
          2223 => x"2a",
          2224 => x"78",
          2225 => x"38",
          2226 => x"38",
          2227 => x"08",
          2228 => x"53",
          2229 => x"aa",
          2230 => x"c8",
          2231 => x"88",
          2232 => x"e8",
          2233 => x"3f",
          2234 => x"09",
          2235 => x"38",
          2236 => x"51",
          2237 => x"79",
          2238 => x"3f",
          2239 => x"54",
          2240 => x"08",
          2241 => x"58",
          2242 => x"c8",
          2243 => x"0d",
          2244 => x"0d",
          2245 => x"5c",
          2246 => x"57",
          2247 => x"73",
          2248 => x"81",
          2249 => x"78",
          2250 => x"56",
          2251 => x"98",
          2252 => x"70",
          2253 => x"33",
          2254 => x"73",
          2255 => x"81",
          2256 => x"75",
          2257 => x"38",
          2258 => x"88",
          2259 => x"98",
          2260 => x"52",
          2261 => x"3f",
          2262 => x"08",
          2263 => x"74",
          2264 => x"ca",
          2265 => x"c8",
          2266 => x"38",
          2267 => x"55",
          2268 => x"88",
          2269 => x"2e",
          2270 => x"39",
          2271 => x"ab",
          2272 => x"5a",
          2273 => x"11",
          2274 => x"51",
          2275 => x"81",
          2276 => x"80",
          2277 => x"7a",
          2278 => x"77",
          2279 => x"3f",
          2280 => x"08",
          2281 => x"55",
          2282 => x"74",
          2283 => x"81",
          2284 => x"ff",
          2285 => x"82",
          2286 => x"8e",
          2287 => x"73",
          2288 => x"0c",
          2289 => x"04",
          2290 => x"b0",
          2291 => x"84",
          2292 => x"05",
          2293 => x"80",
          2294 => x"34",
          2295 => x"33",
          2296 => x"90",
          2297 => x"38",
          2298 => x"33",
          2299 => x"9a",
          2300 => x"eb",
          2301 => x"f8",
          2302 => x"f5",
          2303 => x"f8",
          2304 => x"2e",
          2305 => x"93",
          2306 => x"b8",
          2307 => x"f8",
          2308 => x"bb",
          2309 => x"f8",
          2310 => x"2e",
          2311 => x"e4",
          2312 => x"a4",
          2313 => x"39",
          2314 => x"08",
          2315 => x"52",
          2316 => x"52",
          2317 => x"b0",
          2318 => x"c8",
          2319 => x"f8",
          2320 => x"2e",
          2321 => x"80",
          2322 => x"f8",
          2323 => x"d3",
          2324 => x"f8",
          2325 => x"80",
          2326 => x"c8",
          2327 => x"38",
          2328 => x"08",
          2329 => x"17",
          2330 => x"74",
          2331 => x"74",
          2332 => x"52",
          2333 => x"b4",
          2334 => x"2e",
          2335 => x"ff",
          2336 => x"39",
          2337 => x"f5",
          2338 => x"3d",
          2339 => x"3f",
          2340 => x"08",
          2341 => x"98",
          2342 => x"78",
          2343 => x"38",
          2344 => x"06",
          2345 => x"33",
          2346 => x"70",
          2347 => x"f8",
          2348 => x"98",
          2349 => x"2c",
          2350 => x"05",
          2351 => x"81",
          2352 => x"70",
          2353 => x"33",
          2354 => x"51",
          2355 => x"59",
          2356 => x"56",
          2357 => x"80",
          2358 => x"74",
          2359 => x"74",
          2360 => x"29",
          2361 => x"05",
          2362 => x"51",
          2363 => x"24",
          2364 => x"76",
          2365 => x"77",
          2366 => x"3f",
          2367 => x"08",
          2368 => x"54",
          2369 => x"d7",
          2370 => x"f8",
          2371 => x"56",
          2372 => x"81",
          2373 => x"81",
          2374 => x"70",
          2375 => x"81",
          2376 => x"51",
          2377 => x"26",
          2378 => x"53",
          2379 => x"51",
          2380 => x"81",
          2381 => x"81",
          2382 => x"73",
          2383 => x"39",
          2384 => x"80",
          2385 => x"38",
          2386 => x"74",
          2387 => x"34",
          2388 => x"70",
          2389 => x"f8",
          2390 => x"98",
          2391 => x"2c",
          2392 => x"70",
          2393 => x"e4",
          2394 => x"5e",
          2395 => x"57",
          2396 => x"74",
          2397 => x"81",
          2398 => x"38",
          2399 => x"14",
          2400 => x"80",
          2401 => x"ec",
          2402 => x"81",
          2403 => x"92",
          2404 => x"f8",
          2405 => x"81",
          2406 => x"78",
          2407 => x"75",
          2408 => x"54",
          2409 => x"fd",
          2410 => x"84",
          2411 => x"d0",
          2412 => x"08",
          2413 => x"f4",
          2414 => x"7e",
          2415 => x"38",
          2416 => x"33",
          2417 => x"27",
          2418 => x"98",
          2419 => x"2c",
          2420 => x"75",
          2421 => x"74",
          2422 => x"33",
          2423 => x"74",
          2424 => x"29",
          2425 => x"05",
          2426 => x"81",
          2427 => x"56",
          2428 => x"39",
          2429 => x"33",
          2430 => x"54",
          2431 => x"f4",
          2432 => x"54",
          2433 => x"74",
          2434 => x"f0",
          2435 => x"7e",
          2436 => x"81",
          2437 => x"81",
          2438 => x"81",
          2439 => x"70",
          2440 => x"29",
          2441 => x"05",
          2442 => x"81",
          2443 => x"5a",
          2444 => x"74",
          2445 => x"38",
          2446 => x"33",
          2447 => x"c7",
          2448 => x"80",
          2449 => x"80",
          2450 => x"98",
          2451 => x"f0",
          2452 => x"55",
          2453 => x"e0",
          2454 => x"f4",
          2455 => x"2b",
          2456 => x"81",
          2457 => x"5a",
          2458 => x"74",
          2459 => x"9a",
          2460 => x"e8",
          2461 => x"81",
          2462 => x"81",
          2463 => x"70",
          2464 => x"f8",
          2465 => x"51",
          2466 => x"24",
          2467 => x"fa",
          2468 => x"f4",
          2469 => x"ff",
          2470 => x"73",
          2471 => x"ea",
          2472 => x"f0",
          2473 => x"54",
          2474 => x"f0",
          2475 => x"54",
          2476 => x"f4",
          2477 => x"e7",
          2478 => x"f8",
          2479 => x"98",
          2480 => x"2c",
          2481 => x"33",
          2482 => x"57",
          2483 => x"a7",
          2484 => x"54",
          2485 => x"74",
          2486 => x"51",
          2487 => x"74",
          2488 => x"29",
          2489 => x"05",
          2490 => x"81",
          2491 => x"58",
          2492 => x"75",
          2493 => x"a0",
          2494 => x"3f",
          2495 => x"33",
          2496 => x"70",
          2497 => x"f8",
          2498 => x"51",
          2499 => x"74",
          2500 => x"38",
          2501 => x"ef",
          2502 => x"80",
          2503 => x"80",
          2504 => x"98",
          2505 => x"f0",
          2506 => x"55",
          2507 => x"e4",
          2508 => x"39",
          2509 => x"33",
          2510 => x"80",
          2511 => x"51",
          2512 => x"81",
          2513 => x"79",
          2514 => x"3f",
          2515 => x"08",
          2516 => x"54",
          2517 => x"81",
          2518 => x"54",
          2519 => x"84",
          2520 => x"53",
          2521 => x"51",
          2522 => x"84",
          2523 => x"7a",
          2524 => x"39",
          2525 => x"33",
          2526 => x"2e",
          2527 => x"88",
          2528 => x"3f",
          2529 => x"33",
          2530 => x"73",
          2531 => x"34",
          2532 => x"06",
          2533 => x"81",
          2534 => x"81",
          2535 => x"55",
          2536 => x"2e",
          2537 => x"ff",
          2538 => x"81",
          2539 => x"74",
          2540 => x"98",
          2541 => x"ff",
          2542 => x"55",
          2543 => x"a7",
          2544 => x"54",
          2545 => x"74",
          2546 => x"51",
          2547 => x"74",
          2548 => x"29",
          2549 => x"05",
          2550 => x"81",
          2551 => x"58",
          2552 => x"75",
          2553 => x"a0",
          2554 => x"3f",
          2555 => x"33",
          2556 => x"70",
          2557 => x"f8",
          2558 => x"51",
          2559 => x"74",
          2560 => x"38",
          2561 => x"ff",
          2562 => x"80",
          2563 => x"80",
          2564 => x"98",
          2565 => x"f0",
          2566 => x"55",
          2567 => x"e4",
          2568 => x"39",
          2569 => x"33",
          2570 => x"06",
          2571 => x"33",
          2572 => x"74",
          2573 => x"d2",
          2574 => x"54",
          2575 => x"f4",
          2576 => x"70",
          2577 => x"e4",
          2578 => x"f8",
          2579 => x"81",
          2580 => x"f8",
          2581 => x"56",
          2582 => x"26",
          2583 => x"aa",
          2584 => x"38",
          2585 => x"08",
          2586 => x"2e",
          2587 => x"51",
          2588 => x"81",
          2589 => x"81",
          2590 => x"81",
          2591 => x"81",
          2592 => x"05",
          2593 => x"79",
          2594 => x"3f",
          2595 => x"c1",
          2596 => x"29",
          2597 => x"05",
          2598 => x"56",
          2599 => x"2e",
          2600 => x"51",
          2601 => x"81",
          2602 => x"81",
          2603 => x"81",
          2604 => x"81",
          2605 => x"05",
          2606 => x"79",
          2607 => x"3f",
          2608 => x"80",
          2609 => x"08",
          2610 => x"2e",
          2611 => x"74",
          2612 => x"3f",
          2613 => x"7a",
          2614 => x"81",
          2615 => x"81",
          2616 => x"55",
          2617 => x"89",
          2618 => x"ca",
          2619 => x"c8",
          2620 => x"29",
          2621 => x"05",
          2622 => x"56",
          2623 => x"2e",
          2624 => x"51",
          2625 => x"81",
          2626 => x"81",
          2627 => x"81",
          2628 => x"81",
          2629 => x"05",
          2630 => x"79",
          2631 => x"3f",
          2632 => x"73",
          2633 => x"5b",
          2634 => x"08",
          2635 => x"2e",
          2636 => x"74",
          2637 => x"3f",
          2638 => x"08",
          2639 => x"34",
          2640 => x"08",
          2641 => x"81",
          2642 => x"52",
          2643 => x"e2",
          2644 => x"f4",
          2645 => x"f0",
          2646 => x"51",
          2647 => x"f6",
          2648 => x"f8",
          2649 => x"81",
          2650 => x"f8",
          2651 => x"56",
          2652 => x"27",
          2653 => x"81",
          2654 => x"81",
          2655 => x"74",
          2656 => x"52",
          2657 => x"3f",
          2658 => x"81",
          2659 => x"54",
          2660 => x"f5",
          2661 => x"51",
          2662 => x"81",
          2663 => x"ff",
          2664 => x"81",
          2665 => x"f5",
          2666 => x"0b",
          2667 => x"34",
          2668 => x"f8",
          2669 => x"81",
          2670 => x"af",
          2671 => x"ff",
          2672 => x"8f",
          2673 => x"81",
          2674 => x"26",
          2675 => x"f5",
          2676 => x"52",
          2677 => x"c8",
          2678 => x"0d",
          2679 => x"0d",
          2680 => x"33",
          2681 => x"9f",
          2682 => x"53",
          2683 => x"81",
          2684 => x"38",
          2685 => x"87",
          2686 => x"11",
          2687 => x"54",
          2688 => x"84",
          2689 => x"54",
          2690 => x"87",
          2691 => x"11",
          2692 => x"0c",
          2693 => x"c0",
          2694 => x"70",
          2695 => x"70",
          2696 => x"51",
          2697 => x"8a",
          2698 => x"98",
          2699 => x"70",
          2700 => x"08",
          2701 => x"06",
          2702 => x"38",
          2703 => x"8c",
          2704 => x"80",
          2705 => x"71",
          2706 => x"14",
          2707 => x"b0",
          2708 => x"70",
          2709 => x"0c",
          2710 => x"04",
          2711 => x"60",
          2712 => x"8c",
          2713 => x"33",
          2714 => x"5b",
          2715 => x"5a",
          2716 => x"81",
          2717 => x"81",
          2718 => x"52",
          2719 => x"38",
          2720 => x"84",
          2721 => x"92",
          2722 => x"c0",
          2723 => x"87",
          2724 => x"13",
          2725 => x"57",
          2726 => x"0b",
          2727 => x"8c",
          2728 => x"0c",
          2729 => x"75",
          2730 => x"2a",
          2731 => x"51",
          2732 => x"80",
          2733 => x"7b",
          2734 => x"7b",
          2735 => x"5d",
          2736 => x"59",
          2737 => x"06",
          2738 => x"73",
          2739 => x"81",
          2740 => x"ff",
          2741 => x"72",
          2742 => x"38",
          2743 => x"8c",
          2744 => x"c3",
          2745 => x"98",
          2746 => x"71",
          2747 => x"38",
          2748 => x"2e",
          2749 => x"76",
          2750 => x"92",
          2751 => x"72",
          2752 => x"06",
          2753 => x"f7",
          2754 => x"5a",
          2755 => x"80",
          2756 => x"70",
          2757 => x"5a",
          2758 => x"80",
          2759 => x"73",
          2760 => x"06",
          2761 => x"38",
          2762 => x"fe",
          2763 => x"fc",
          2764 => x"52",
          2765 => x"83",
          2766 => x"71",
          2767 => x"f8",
          2768 => x"3d",
          2769 => x"3d",
          2770 => x"64",
          2771 => x"bf",
          2772 => x"40",
          2773 => x"59",
          2774 => x"58",
          2775 => x"81",
          2776 => x"81",
          2777 => x"52",
          2778 => x"09",
          2779 => x"b1",
          2780 => x"84",
          2781 => x"92",
          2782 => x"c0",
          2783 => x"87",
          2784 => x"13",
          2785 => x"56",
          2786 => x"87",
          2787 => x"0c",
          2788 => x"82",
          2789 => x"58",
          2790 => x"84",
          2791 => x"06",
          2792 => x"71",
          2793 => x"38",
          2794 => x"05",
          2795 => x"0c",
          2796 => x"73",
          2797 => x"81",
          2798 => x"71",
          2799 => x"38",
          2800 => x"8c",
          2801 => x"d0",
          2802 => x"98",
          2803 => x"71",
          2804 => x"38",
          2805 => x"2e",
          2806 => x"76",
          2807 => x"92",
          2808 => x"72",
          2809 => x"06",
          2810 => x"f7",
          2811 => x"59",
          2812 => x"1a",
          2813 => x"06",
          2814 => x"59",
          2815 => x"80",
          2816 => x"73",
          2817 => x"06",
          2818 => x"38",
          2819 => x"fe",
          2820 => x"fc",
          2821 => x"52",
          2822 => x"83",
          2823 => x"71",
          2824 => x"f8",
          2825 => x"3d",
          2826 => x"3d",
          2827 => x"84",
          2828 => x"33",
          2829 => x"a7",
          2830 => x"54",
          2831 => x"fa",
          2832 => x"f8",
          2833 => x"06",
          2834 => x"72",
          2835 => x"85",
          2836 => x"98",
          2837 => x"56",
          2838 => x"80",
          2839 => x"76",
          2840 => x"74",
          2841 => x"c0",
          2842 => x"54",
          2843 => x"2e",
          2844 => x"d4",
          2845 => x"2e",
          2846 => x"80",
          2847 => x"08",
          2848 => x"70",
          2849 => x"51",
          2850 => x"2e",
          2851 => x"c0",
          2852 => x"52",
          2853 => x"87",
          2854 => x"08",
          2855 => x"38",
          2856 => x"87",
          2857 => x"14",
          2858 => x"70",
          2859 => x"52",
          2860 => x"96",
          2861 => x"92",
          2862 => x"0a",
          2863 => x"39",
          2864 => x"0c",
          2865 => x"39",
          2866 => x"54",
          2867 => x"c8",
          2868 => x"0d",
          2869 => x"0d",
          2870 => x"33",
          2871 => x"88",
          2872 => x"f8",
          2873 => x"51",
          2874 => x"04",
          2875 => x"75",
          2876 => x"82",
          2877 => x"90",
          2878 => x"2b",
          2879 => x"33",
          2880 => x"88",
          2881 => x"71",
          2882 => x"c8",
          2883 => x"54",
          2884 => x"85",
          2885 => x"ff",
          2886 => x"02",
          2887 => x"05",
          2888 => x"70",
          2889 => x"05",
          2890 => x"88",
          2891 => x"72",
          2892 => x"0d",
          2893 => x"0d",
          2894 => x"52",
          2895 => x"81",
          2896 => x"70",
          2897 => x"70",
          2898 => x"05",
          2899 => x"88",
          2900 => x"72",
          2901 => x"54",
          2902 => x"2a",
          2903 => x"34",
          2904 => x"04",
          2905 => x"76",
          2906 => x"54",
          2907 => x"2e",
          2908 => x"70",
          2909 => x"33",
          2910 => x"05",
          2911 => x"11",
          2912 => x"84",
          2913 => x"fe",
          2914 => x"77",
          2915 => x"53",
          2916 => x"81",
          2917 => x"ff",
          2918 => x"f4",
          2919 => x"0d",
          2920 => x"0d",
          2921 => x"56",
          2922 => x"70",
          2923 => x"33",
          2924 => x"05",
          2925 => x"71",
          2926 => x"56",
          2927 => x"72",
          2928 => x"38",
          2929 => x"e2",
          2930 => x"f8",
          2931 => x"3d",
          2932 => x"3d",
          2933 => x"54",
          2934 => x"71",
          2935 => x"38",
          2936 => x"70",
          2937 => x"f3",
          2938 => x"81",
          2939 => x"84",
          2940 => x"80",
          2941 => x"c8",
          2942 => x"0b",
          2943 => x"0c",
          2944 => x"0d",
          2945 => x"0b",
          2946 => x"56",
          2947 => x"2e",
          2948 => x"81",
          2949 => x"08",
          2950 => x"70",
          2951 => x"33",
          2952 => x"a2",
          2953 => x"c8",
          2954 => x"09",
          2955 => x"38",
          2956 => x"08",
          2957 => x"b0",
          2958 => x"a4",
          2959 => x"9c",
          2960 => x"56",
          2961 => x"27",
          2962 => x"16",
          2963 => x"82",
          2964 => x"06",
          2965 => x"54",
          2966 => x"78",
          2967 => x"33",
          2968 => x"3f",
          2969 => x"5a",
          2970 => x"c8",
          2971 => x"0d",
          2972 => x"0d",
          2973 => x"56",
          2974 => x"b0",
          2975 => x"af",
          2976 => x"fe",
          2977 => x"f8",
          2978 => x"81",
          2979 => x"9f",
          2980 => x"74",
          2981 => x"52",
          2982 => x"51",
          2983 => x"81",
          2984 => x"80",
          2985 => x"ff",
          2986 => x"74",
          2987 => x"76",
          2988 => x"0c",
          2989 => x"04",
          2990 => x"7a",
          2991 => x"fe",
          2992 => x"f8",
          2993 => x"81",
          2994 => x"81",
          2995 => x"33",
          2996 => x"2e",
          2997 => x"80",
          2998 => x"17",
          2999 => x"81",
          3000 => x"06",
          3001 => x"84",
          3002 => x"f8",
          3003 => x"b4",
          3004 => x"56",
          3005 => x"82",
          3006 => x"84",
          3007 => x"fc",
          3008 => x"8b",
          3009 => x"52",
          3010 => x"a9",
          3011 => x"85",
          3012 => x"84",
          3013 => x"fc",
          3014 => x"17",
          3015 => x"9c",
          3016 => x"91",
          3017 => x"08",
          3018 => x"17",
          3019 => x"3f",
          3020 => x"81",
          3021 => x"19",
          3022 => x"53",
          3023 => x"17",
          3024 => x"82",
          3025 => x"18",
          3026 => x"80",
          3027 => x"33",
          3028 => x"3f",
          3029 => x"08",
          3030 => x"38",
          3031 => x"81",
          3032 => x"8a",
          3033 => x"fb",
          3034 => x"fe",
          3035 => x"08",
          3036 => x"56",
          3037 => x"74",
          3038 => x"38",
          3039 => x"75",
          3040 => x"16",
          3041 => x"53",
          3042 => x"c8",
          3043 => x"0d",
          3044 => x"0d",
          3045 => x"08",
          3046 => x"81",
          3047 => x"df",
          3048 => x"15",
          3049 => x"d7",
          3050 => x"33",
          3051 => x"82",
          3052 => x"38",
          3053 => x"89",
          3054 => x"2e",
          3055 => x"bf",
          3056 => x"2e",
          3057 => x"81",
          3058 => x"81",
          3059 => x"89",
          3060 => x"08",
          3061 => x"52",
          3062 => x"3f",
          3063 => x"08",
          3064 => x"74",
          3065 => x"14",
          3066 => x"81",
          3067 => x"2a",
          3068 => x"05",
          3069 => x"57",
          3070 => x"f5",
          3071 => x"c8",
          3072 => x"38",
          3073 => x"06",
          3074 => x"33",
          3075 => x"78",
          3076 => x"06",
          3077 => x"5c",
          3078 => x"53",
          3079 => x"38",
          3080 => x"06",
          3081 => x"39",
          3082 => x"a4",
          3083 => x"52",
          3084 => x"bd",
          3085 => x"c8",
          3086 => x"38",
          3087 => x"fe",
          3088 => x"b4",
          3089 => x"8d",
          3090 => x"c8",
          3091 => x"ff",
          3092 => x"39",
          3093 => x"a4",
          3094 => x"52",
          3095 => x"91",
          3096 => x"c8",
          3097 => x"76",
          3098 => x"fc",
          3099 => x"b4",
          3100 => x"f8",
          3101 => x"c8",
          3102 => x"06",
          3103 => x"81",
          3104 => x"f8",
          3105 => x"3d",
          3106 => x"3d",
          3107 => x"7e",
          3108 => x"82",
          3109 => x"27",
          3110 => x"76",
          3111 => x"27",
          3112 => x"75",
          3113 => x"79",
          3114 => x"38",
          3115 => x"89",
          3116 => x"2e",
          3117 => x"80",
          3118 => x"2e",
          3119 => x"81",
          3120 => x"81",
          3121 => x"89",
          3122 => x"08",
          3123 => x"52",
          3124 => x"3f",
          3125 => x"08",
          3126 => x"c8",
          3127 => x"38",
          3128 => x"06",
          3129 => x"81",
          3130 => x"06",
          3131 => x"77",
          3132 => x"2e",
          3133 => x"84",
          3134 => x"06",
          3135 => x"06",
          3136 => x"53",
          3137 => x"81",
          3138 => x"34",
          3139 => x"a4",
          3140 => x"52",
          3141 => x"d9",
          3142 => x"c8",
          3143 => x"f8",
          3144 => x"94",
          3145 => x"ff",
          3146 => x"05",
          3147 => x"54",
          3148 => x"38",
          3149 => x"74",
          3150 => x"06",
          3151 => x"07",
          3152 => x"74",
          3153 => x"39",
          3154 => x"a4",
          3155 => x"52",
          3156 => x"9d",
          3157 => x"c8",
          3158 => x"f8",
          3159 => x"d8",
          3160 => x"ff",
          3161 => x"76",
          3162 => x"06",
          3163 => x"05",
          3164 => x"3f",
          3165 => x"87",
          3166 => x"08",
          3167 => x"51",
          3168 => x"81",
          3169 => x"59",
          3170 => x"08",
          3171 => x"f0",
          3172 => x"82",
          3173 => x"06",
          3174 => x"05",
          3175 => x"54",
          3176 => x"3f",
          3177 => x"08",
          3178 => x"74",
          3179 => x"51",
          3180 => x"81",
          3181 => x"34",
          3182 => x"c8",
          3183 => x"0d",
          3184 => x"0d",
          3185 => x"72",
          3186 => x"56",
          3187 => x"27",
          3188 => x"98",
          3189 => x"9d",
          3190 => x"2e",
          3191 => x"53",
          3192 => x"51",
          3193 => x"81",
          3194 => x"54",
          3195 => x"08",
          3196 => x"93",
          3197 => x"80",
          3198 => x"54",
          3199 => x"81",
          3200 => x"54",
          3201 => x"74",
          3202 => x"fb",
          3203 => x"f8",
          3204 => x"81",
          3205 => x"80",
          3206 => x"38",
          3207 => x"08",
          3208 => x"38",
          3209 => x"08",
          3210 => x"38",
          3211 => x"52",
          3212 => x"d6",
          3213 => x"c8",
          3214 => x"98",
          3215 => x"11",
          3216 => x"57",
          3217 => x"74",
          3218 => x"81",
          3219 => x"0c",
          3220 => x"81",
          3221 => x"84",
          3222 => x"55",
          3223 => x"ff",
          3224 => x"54",
          3225 => x"c8",
          3226 => x"0d",
          3227 => x"0d",
          3228 => x"08",
          3229 => x"79",
          3230 => x"17",
          3231 => x"80",
          3232 => x"98",
          3233 => x"26",
          3234 => x"58",
          3235 => x"52",
          3236 => x"fd",
          3237 => x"74",
          3238 => x"08",
          3239 => x"38",
          3240 => x"08",
          3241 => x"c8",
          3242 => x"82",
          3243 => x"17",
          3244 => x"c8",
          3245 => x"c7",
          3246 => x"90",
          3247 => x"56",
          3248 => x"2e",
          3249 => x"77",
          3250 => x"81",
          3251 => x"38",
          3252 => x"98",
          3253 => x"26",
          3254 => x"56",
          3255 => x"51",
          3256 => x"80",
          3257 => x"c8",
          3258 => x"09",
          3259 => x"38",
          3260 => x"08",
          3261 => x"c8",
          3262 => x"30",
          3263 => x"80",
          3264 => x"07",
          3265 => x"08",
          3266 => x"55",
          3267 => x"ef",
          3268 => x"c8",
          3269 => x"95",
          3270 => x"08",
          3271 => x"27",
          3272 => x"98",
          3273 => x"89",
          3274 => x"85",
          3275 => x"db",
          3276 => x"81",
          3277 => x"17",
          3278 => x"89",
          3279 => x"75",
          3280 => x"ac",
          3281 => x"7a",
          3282 => x"3f",
          3283 => x"08",
          3284 => x"38",
          3285 => x"f8",
          3286 => x"2e",
          3287 => x"86",
          3288 => x"c8",
          3289 => x"f8",
          3290 => x"70",
          3291 => x"07",
          3292 => x"7c",
          3293 => x"55",
          3294 => x"f8",
          3295 => x"2e",
          3296 => x"ff",
          3297 => x"55",
          3298 => x"ff",
          3299 => x"76",
          3300 => x"3f",
          3301 => x"08",
          3302 => x"08",
          3303 => x"f8",
          3304 => x"80",
          3305 => x"55",
          3306 => x"94",
          3307 => x"2e",
          3308 => x"53",
          3309 => x"51",
          3310 => x"81",
          3311 => x"55",
          3312 => x"75",
          3313 => x"98",
          3314 => x"05",
          3315 => x"56",
          3316 => x"26",
          3317 => x"15",
          3318 => x"84",
          3319 => x"07",
          3320 => x"18",
          3321 => x"ff",
          3322 => x"2e",
          3323 => x"39",
          3324 => x"39",
          3325 => x"08",
          3326 => x"81",
          3327 => x"74",
          3328 => x"0c",
          3329 => x"04",
          3330 => x"7a",
          3331 => x"f3",
          3332 => x"f8",
          3333 => x"81",
          3334 => x"c8",
          3335 => x"38",
          3336 => x"51",
          3337 => x"81",
          3338 => x"81",
          3339 => x"b0",
          3340 => x"84",
          3341 => x"52",
          3342 => x"52",
          3343 => x"3f",
          3344 => x"39",
          3345 => x"8a",
          3346 => x"75",
          3347 => x"38",
          3348 => x"19",
          3349 => x"81",
          3350 => x"ed",
          3351 => x"f8",
          3352 => x"2e",
          3353 => x"15",
          3354 => x"70",
          3355 => x"07",
          3356 => x"53",
          3357 => x"75",
          3358 => x"0c",
          3359 => x"04",
          3360 => x"7a",
          3361 => x"58",
          3362 => x"f0",
          3363 => x"80",
          3364 => x"9f",
          3365 => x"80",
          3366 => x"90",
          3367 => x"17",
          3368 => x"aa",
          3369 => x"53",
          3370 => x"88",
          3371 => x"08",
          3372 => x"38",
          3373 => x"53",
          3374 => x"17",
          3375 => x"72",
          3376 => x"fe",
          3377 => x"08",
          3378 => x"80",
          3379 => x"16",
          3380 => x"2b",
          3381 => x"75",
          3382 => x"73",
          3383 => x"f5",
          3384 => x"f8",
          3385 => x"81",
          3386 => x"ff",
          3387 => x"81",
          3388 => x"c8",
          3389 => x"38",
          3390 => x"81",
          3391 => x"26",
          3392 => x"58",
          3393 => x"73",
          3394 => x"39",
          3395 => x"51",
          3396 => x"81",
          3397 => x"98",
          3398 => x"94",
          3399 => x"17",
          3400 => x"58",
          3401 => x"9a",
          3402 => x"81",
          3403 => x"74",
          3404 => x"98",
          3405 => x"83",
          3406 => x"b4",
          3407 => x"0c",
          3408 => x"81",
          3409 => x"8a",
          3410 => x"f8",
          3411 => x"70",
          3412 => x"08",
          3413 => x"57",
          3414 => x"0a",
          3415 => x"38",
          3416 => x"15",
          3417 => x"08",
          3418 => x"72",
          3419 => x"cb",
          3420 => x"ff",
          3421 => x"81",
          3422 => x"13",
          3423 => x"94",
          3424 => x"74",
          3425 => x"85",
          3426 => x"22",
          3427 => x"73",
          3428 => x"38",
          3429 => x"8a",
          3430 => x"05",
          3431 => x"06",
          3432 => x"8a",
          3433 => x"73",
          3434 => x"3f",
          3435 => x"08",
          3436 => x"81",
          3437 => x"c8",
          3438 => x"ff",
          3439 => x"81",
          3440 => x"ff",
          3441 => x"38",
          3442 => x"81",
          3443 => x"26",
          3444 => x"7b",
          3445 => x"98",
          3446 => x"55",
          3447 => x"94",
          3448 => x"73",
          3449 => x"3f",
          3450 => x"08",
          3451 => x"81",
          3452 => x"80",
          3453 => x"38",
          3454 => x"f8",
          3455 => x"2e",
          3456 => x"55",
          3457 => x"08",
          3458 => x"38",
          3459 => x"08",
          3460 => x"fb",
          3461 => x"f8",
          3462 => x"38",
          3463 => x"0c",
          3464 => x"51",
          3465 => x"81",
          3466 => x"98",
          3467 => x"90",
          3468 => x"16",
          3469 => x"15",
          3470 => x"74",
          3471 => x"0c",
          3472 => x"04",
          3473 => x"7b",
          3474 => x"5b",
          3475 => x"52",
          3476 => x"ac",
          3477 => x"c8",
          3478 => x"f8",
          3479 => x"ec",
          3480 => x"c8",
          3481 => x"17",
          3482 => x"51",
          3483 => x"81",
          3484 => x"54",
          3485 => x"08",
          3486 => x"81",
          3487 => x"9c",
          3488 => x"33",
          3489 => x"72",
          3490 => x"09",
          3491 => x"38",
          3492 => x"f8",
          3493 => x"72",
          3494 => x"55",
          3495 => x"53",
          3496 => x"8e",
          3497 => x"56",
          3498 => x"09",
          3499 => x"38",
          3500 => x"f8",
          3501 => x"81",
          3502 => x"fd",
          3503 => x"f8",
          3504 => x"81",
          3505 => x"80",
          3506 => x"38",
          3507 => x"09",
          3508 => x"38",
          3509 => x"81",
          3510 => x"8b",
          3511 => x"fd",
          3512 => x"9a",
          3513 => x"eb",
          3514 => x"f8",
          3515 => x"ff",
          3516 => x"70",
          3517 => x"53",
          3518 => x"09",
          3519 => x"38",
          3520 => x"eb",
          3521 => x"f8",
          3522 => x"2b",
          3523 => x"72",
          3524 => x"0c",
          3525 => x"04",
          3526 => x"77",
          3527 => x"ff",
          3528 => x"9a",
          3529 => x"55",
          3530 => x"76",
          3531 => x"53",
          3532 => x"09",
          3533 => x"38",
          3534 => x"52",
          3535 => x"eb",
          3536 => x"3d",
          3537 => x"3d",
          3538 => x"5b",
          3539 => x"08",
          3540 => x"15",
          3541 => x"81",
          3542 => x"15",
          3543 => x"51",
          3544 => x"81",
          3545 => x"58",
          3546 => x"08",
          3547 => x"9c",
          3548 => x"33",
          3549 => x"86",
          3550 => x"80",
          3551 => x"13",
          3552 => x"06",
          3553 => x"06",
          3554 => x"72",
          3555 => x"81",
          3556 => x"53",
          3557 => x"2e",
          3558 => x"53",
          3559 => x"a9",
          3560 => x"74",
          3561 => x"72",
          3562 => x"38",
          3563 => x"99",
          3564 => x"c8",
          3565 => x"06",
          3566 => x"88",
          3567 => x"06",
          3568 => x"54",
          3569 => x"a0",
          3570 => x"74",
          3571 => x"3f",
          3572 => x"08",
          3573 => x"c8",
          3574 => x"98",
          3575 => x"fa",
          3576 => x"80",
          3577 => x"0c",
          3578 => x"c8",
          3579 => x"0d",
          3580 => x"0d",
          3581 => x"57",
          3582 => x"73",
          3583 => x"3f",
          3584 => x"08",
          3585 => x"c8",
          3586 => x"98",
          3587 => x"75",
          3588 => x"3f",
          3589 => x"08",
          3590 => x"c8",
          3591 => x"a0",
          3592 => x"c8",
          3593 => x"14",
          3594 => x"db",
          3595 => x"a0",
          3596 => x"14",
          3597 => x"ac",
          3598 => x"83",
          3599 => x"81",
          3600 => x"87",
          3601 => x"fd",
          3602 => x"70",
          3603 => x"08",
          3604 => x"55",
          3605 => x"3f",
          3606 => x"08",
          3607 => x"13",
          3608 => x"73",
          3609 => x"83",
          3610 => x"3d",
          3611 => x"3d",
          3612 => x"57",
          3613 => x"89",
          3614 => x"17",
          3615 => x"81",
          3616 => x"70",
          3617 => x"55",
          3618 => x"08",
          3619 => x"81",
          3620 => x"52",
          3621 => x"a8",
          3622 => x"2e",
          3623 => x"84",
          3624 => x"52",
          3625 => x"09",
          3626 => x"38",
          3627 => x"81",
          3628 => x"81",
          3629 => x"73",
          3630 => x"55",
          3631 => x"55",
          3632 => x"c5",
          3633 => x"88",
          3634 => x"0b",
          3635 => x"9c",
          3636 => x"8b",
          3637 => x"17",
          3638 => x"08",
          3639 => x"52",
          3640 => x"81",
          3641 => x"76",
          3642 => x"51",
          3643 => x"81",
          3644 => x"86",
          3645 => x"12",
          3646 => x"3f",
          3647 => x"08",
          3648 => x"88",
          3649 => x"f3",
          3650 => x"70",
          3651 => x"80",
          3652 => x"51",
          3653 => x"af",
          3654 => x"81",
          3655 => x"dc",
          3656 => x"74",
          3657 => x"38",
          3658 => x"88",
          3659 => x"39",
          3660 => x"80",
          3661 => x"56",
          3662 => x"af",
          3663 => x"06",
          3664 => x"56",
          3665 => x"32",
          3666 => x"80",
          3667 => x"51",
          3668 => x"dc",
          3669 => x"1c",
          3670 => x"33",
          3671 => x"9f",
          3672 => x"ff",
          3673 => x"1c",
          3674 => x"7a",
          3675 => x"3f",
          3676 => x"08",
          3677 => x"39",
          3678 => x"a0",
          3679 => x"5e",
          3680 => x"52",
          3681 => x"ff",
          3682 => x"59",
          3683 => x"33",
          3684 => x"ae",
          3685 => x"06",
          3686 => x"78",
          3687 => x"81",
          3688 => x"32",
          3689 => x"9f",
          3690 => x"26",
          3691 => x"53",
          3692 => x"73",
          3693 => x"17",
          3694 => x"34",
          3695 => x"db",
          3696 => x"32",
          3697 => x"9f",
          3698 => x"54",
          3699 => x"2e",
          3700 => x"80",
          3701 => x"75",
          3702 => x"bd",
          3703 => x"7e",
          3704 => x"a0",
          3705 => x"bd",
          3706 => x"82",
          3707 => x"18",
          3708 => x"1a",
          3709 => x"a0",
          3710 => x"fc",
          3711 => x"32",
          3712 => x"80",
          3713 => x"30",
          3714 => x"71",
          3715 => x"51",
          3716 => x"55",
          3717 => x"ac",
          3718 => x"81",
          3719 => x"78",
          3720 => x"51",
          3721 => x"af",
          3722 => x"06",
          3723 => x"55",
          3724 => x"32",
          3725 => x"80",
          3726 => x"51",
          3727 => x"db",
          3728 => x"39",
          3729 => x"09",
          3730 => x"38",
          3731 => x"7c",
          3732 => x"54",
          3733 => x"a2",
          3734 => x"32",
          3735 => x"ae",
          3736 => x"72",
          3737 => x"9f",
          3738 => x"51",
          3739 => x"74",
          3740 => x"88",
          3741 => x"fe",
          3742 => x"98",
          3743 => x"80",
          3744 => x"75",
          3745 => x"81",
          3746 => x"33",
          3747 => x"51",
          3748 => x"81",
          3749 => x"80",
          3750 => x"78",
          3751 => x"81",
          3752 => x"5a",
          3753 => x"d2",
          3754 => x"c8",
          3755 => x"80",
          3756 => x"1c",
          3757 => x"27",
          3758 => x"79",
          3759 => x"74",
          3760 => x"7a",
          3761 => x"74",
          3762 => x"39",
          3763 => x"e5",
          3764 => x"fe",
          3765 => x"c8",
          3766 => x"ff",
          3767 => x"73",
          3768 => x"38",
          3769 => x"81",
          3770 => x"54",
          3771 => x"75",
          3772 => x"17",
          3773 => x"39",
          3774 => x"0c",
          3775 => x"99",
          3776 => x"54",
          3777 => x"2e",
          3778 => x"84",
          3779 => x"34",
          3780 => x"76",
          3781 => x"8b",
          3782 => x"81",
          3783 => x"56",
          3784 => x"80",
          3785 => x"1b",
          3786 => x"08",
          3787 => x"51",
          3788 => x"81",
          3789 => x"56",
          3790 => x"08",
          3791 => x"98",
          3792 => x"76",
          3793 => x"3f",
          3794 => x"08",
          3795 => x"c8",
          3796 => x"38",
          3797 => x"70",
          3798 => x"73",
          3799 => x"be",
          3800 => x"33",
          3801 => x"73",
          3802 => x"8b",
          3803 => x"83",
          3804 => x"06",
          3805 => x"73",
          3806 => x"53",
          3807 => x"51",
          3808 => x"81",
          3809 => x"80",
          3810 => x"75",
          3811 => x"f3",
          3812 => x"9f",
          3813 => x"1c",
          3814 => x"74",
          3815 => x"38",
          3816 => x"09",
          3817 => x"e7",
          3818 => x"2a",
          3819 => x"77",
          3820 => x"51",
          3821 => x"2e",
          3822 => x"81",
          3823 => x"80",
          3824 => x"38",
          3825 => x"ab",
          3826 => x"55",
          3827 => x"75",
          3828 => x"73",
          3829 => x"55",
          3830 => x"82",
          3831 => x"06",
          3832 => x"ab",
          3833 => x"33",
          3834 => x"70",
          3835 => x"55",
          3836 => x"2e",
          3837 => x"1b",
          3838 => x"06",
          3839 => x"52",
          3840 => x"db",
          3841 => x"c8",
          3842 => x"0c",
          3843 => x"74",
          3844 => x"0c",
          3845 => x"04",
          3846 => x"7c",
          3847 => x"08",
          3848 => x"55",
          3849 => x"59",
          3850 => x"81",
          3851 => x"70",
          3852 => x"33",
          3853 => x"52",
          3854 => x"2e",
          3855 => x"ee",
          3856 => x"2e",
          3857 => x"81",
          3858 => x"33",
          3859 => x"81",
          3860 => x"52",
          3861 => x"26",
          3862 => x"14",
          3863 => x"06",
          3864 => x"52",
          3865 => x"80",
          3866 => x"0b",
          3867 => x"59",
          3868 => x"7a",
          3869 => x"70",
          3870 => x"33",
          3871 => x"05",
          3872 => x"9f",
          3873 => x"53",
          3874 => x"89",
          3875 => x"70",
          3876 => x"54",
          3877 => x"12",
          3878 => x"26",
          3879 => x"12",
          3880 => x"06",
          3881 => x"30",
          3882 => x"51",
          3883 => x"2e",
          3884 => x"85",
          3885 => x"be",
          3886 => x"74",
          3887 => x"30",
          3888 => x"9f",
          3889 => x"2a",
          3890 => x"54",
          3891 => x"2e",
          3892 => x"15",
          3893 => x"55",
          3894 => x"ff",
          3895 => x"39",
          3896 => x"86",
          3897 => x"7c",
          3898 => x"51",
          3899 => x"f9",
          3900 => x"70",
          3901 => x"0c",
          3902 => x"04",
          3903 => x"78",
          3904 => x"83",
          3905 => x"0b",
          3906 => x"79",
          3907 => x"e2",
          3908 => x"55",
          3909 => x"08",
          3910 => x"84",
          3911 => x"df",
          3912 => x"f8",
          3913 => x"ff",
          3914 => x"83",
          3915 => x"d4",
          3916 => x"81",
          3917 => x"38",
          3918 => x"17",
          3919 => x"74",
          3920 => x"09",
          3921 => x"38",
          3922 => x"81",
          3923 => x"30",
          3924 => x"79",
          3925 => x"54",
          3926 => x"74",
          3927 => x"09",
          3928 => x"38",
          3929 => x"e6",
          3930 => x"ea",
          3931 => x"b1",
          3932 => x"c8",
          3933 => x"f8",
          3934 => x"2e",
          3935 => x"53",
          3936 => x"52",
          3937 => x"51",
          3938 => x"81",
          3939 => x"55",
          3940 => x"08",
          3941 => x"38",
          3942 => x"81",
          3943 => x"88",
          3944 => x"f2",
          3945 => x"02",
          3946 => x"cb",
          3947 => x"55",
          3948 => x"60",
          3949 => x"3f",
          3950 => x"08",
          3951 => x"80",
          3952 => x"c8",
          3953 => x"fc",
          3954 => x"c8",
          3955 => x"81",
          3956 => x"70",
          3957 => x"8c",
          3958 => x"2e",
          3959 => x"73",
          3960 => x"81",
          3961 => x"33",
          3962 => x"80",
          3963 => x"81",
          3964 => x"d7",
          3965 => x"f8",
          3966 => x"ff",
          3967 => x"06",
          3968 => x"98",
          3969 => x"2e",
          3970 => x"74",
          3971 => x"81",
          3972 => x"8a",
          3973 => x"ac",
          3974 => x"39",
          3975 => x"77",
          3976 => x"81",
          3977 => x"33",
          3978 => x"3f",
          3979 => x"08",
          3980 => x"70",
          3981 => x"55",
          3982 => x"86",
          3983 => x"80",
          3984 => x"74",
          3985 => x"81",
          3986 => x"8a",
          3987 => x"f4",
          3988 => x"53",
          3989 => x"fd",
          3990 => x"f8",
          3991 => x"ff",
          3992 => x"82",
          3993 => x"06",
          3994 => x"8c",
          3995 => x"58",
          3996 => x"f6",
          3997 => x"58",
          3998 => x"2e",
          3999 => x"fa",
          4000 => x"e8",
          4001 => x"c8",
          4002 => x"78",
          4003 => x"5a",
          4004 => x"90",
          4005 => x"75",
          4006 => x"38",
          4007 => x"3d",
          4008 => x"70",
          4009 => x"08",
          4010 => x"7a",
          4011 => x"38",
          4012 => x"51",
          4013 => x"81",
          4014 => x"81",
          4015 => x"81",
          4016 => x"38",
          4017 => x"83",
          4018 => x"38",
          4019 => x"84",
          4020 => x"38",
          4021 => x"81",
          4022 => x"38",
          4023 => x"db",
          4024 => x"f8",
          4025 => x"ff",
          4026 => x"72",
          4027 => x"09",
          4028 => x"d0",
          4029 => x"14",
          4030 => x"3f",
          4031 => x"08",
          4032 => x"06",
          4033 => x"38",
          4034 => x"51",
          4035 => x"81",
          4036 => x"58",
          4037 => x"0c",
          4038 => x"33",
          4039 => x"80",
          4040 => x"ff",
          4041 => x"ff",
          4042 => x"55",
          4043 => x"81",
          4044 => x"38",
          4045 => x"06",
          4046 => x"80",
          4047 => x"52",
          4048 => x"8a",
          4049 => x"80",
          4050 => x"ff",
          4051 => x"53",
          4052 => x"86",
          4053 => x"83",
          4054 => x"c5",
          4055 => x"f5",
          4056 => x"c8",
          4057 => x"f8",
          4058 => x"15",
          4059 => x"06",
          4060 => x"76",
          4061 => x"80",
          4062 => x"da",
          4063 => x"f8",
          4064 => x"ff",
          4065 => x"74",
          4066 => x"d4",
          4067 => x"dc",
          4068 => x"c8",
          4069 => x"c2",
          4070 => x"b9",
          4071 => x"c8",
          4072 => x"ff",
          4073 => x"56",
          4074 => x"83",
          4075 => x"14",
          4076 => x"71",
          4077 => x"5a",
          4078 => x"26",
          4079 => x"8a",
          4080 => x"74",
          4081 => x"ff",
          4082 => x"81",
          4083 => x"55",
          4084 => x"08",
          4085 => x"ec",
          4086 => x"c8",
          4087 => x"ff",
          4088 => x"83",
          4089 => x"74",
          4090 => x"26",
          4091 => x"57",
          4092 => x"26",
          4093 => x"57",
          4094 => x"56",
          4095 => x"82",
          4096 => x"15",
          4097 => x"0c",
          4098 => x"0c",
          4099 => x"a4",
          4100 => x"1d",
          4101 => x"54",
          4102 => x"2e",
          4103 => x"af",
          4104 => x"14",
          4105 => x"3f",
          4106 => x"08",
          4107 => x"06",
          4108 => x"72",
          4109 => x"79",
          4110 => x"80",
          4111 => x"d9",
          4112 => x"f8",
          4113 => x"15",
          4114 => x"2b",
          4115 => x"8d",
          4116 => x"2e",
          4117 => x"77",
          4118 => x"0c",
          4119 => x"76",
          4120 => x"38",
          4121 => x"70",
          4122 => x"81",
          4123 => x"53",
          4124 => x"89",
          4125 => x"56",
          4126 => x"08",
          4127 => x"38",
          4128 => x"15",
          4129 => x"8c",
          4130 => x"80",
          4131 => x"34",
          4132 => x"09",
          4133 => x"92",
          4134 => x"14",
          4135 => x"3f",
          4136 => x"08",
          4137 => x"06",
          4138 => x"2e",
          4139 => x"80",
          4140 => x"1b",
          4141 => x"db",
          4142 => x"f8",
          4143 => x"ea",
          4144 => x"c8",
          4145 => x"34",
          4146 => x"51",
          4147 => x"81",
          4148 => x"83",
          4149 => x"53",
          4150 => x"d5",
          4151 => x"06",
          4152 => x"b4",
          4153 => x"84",
          4154 => x"c8",
          4155 => x"85",
          4156 => x"09",
          4157 => x"38",
          4158 => x"51",
          4159 => x"81",
          4160 => x"86",
          4161 => x"f2",
          4162 => x"06",
          4163 => x"9c",
          4164 => x"d8",
          4165 => x"c8",
          4166 => x"0c",
          4167 => x"51",
          4168 => x"81",
          4169 => x"8c",
          4170 => x"74",
          4171 => x"88",
          4172 => x"53",
          4173 => x"88",
          4174 => x"15",
          4175 => x"94",
          4176 => x"56",
          4177 => x"c8",
          4178 => x"0d",
          4179 => x"0d",
          4180 => x"55",
          4181 => x"b9",
          4182 => x"53",
          4183 => x"b1",
          4184 => x"52",
          4185 => x"a9",
          4186 => x"22",
          4187 => x"57",
          4188 => x"2e",
          4189 => x"99",
          4190 => x"33",
          4191 => x"3f",
          4192 => x"08",
          4193 => x"71",
          4194 => x"74",
          4195 => x"83",
          4196 => x"78",
          4197 => x"52",
          4198 => x"c8",
          4199 => x"0d",
          4200 => x"0d",
          4201 => x"33",
          4202 => x"3d",
          4203 => x"56",
          4204 => x"8b",
          4205 => x"81",
          4206 => x"24",
          4207 => x"f8",
          4208 => x"29",
          4209 => x"05",
          4210 => x"55",
          4211 => x"84",
          4212 => x"34",
          4213 => x"80",
          4214 => x"80",
          4215 => x"75",
          4216 => x"75",
          4217 => x"38",
          4218 => x"3d",
          4219 => x"05",
          4220 => x"3f",
          4221 => x"08",
          4222 => x"f8",
          4223 => x"3d",
          4224 => x"3d",
          4225 => x"84",
          4226 => x"05",
          4227 => x"89",
          4228 => x"2e",
          4229 => x"77",
          4230 => x"54",
          4231 => x"05",
          4232 => x"84",
          4233 => x"f6",
          4234 => x"f8",
          4235 => x"81",
          4236 => x"84",
          4237 => x"5c",
          4238 => x"3d",
          4239 => x"ed",
          4240 => x"f8",
          4241 => x"81",
          4242 => x"92",
          4243 => x"d7",
          4244 => x"98",
          4245 => x"73",
          4246 => x"38",
          4247 => x"9c",
          4248 => x"80",
          4249 => x"38",
          4250 => x"95",
          4251 => x"2e",
          4252 => x"aa",
          4253 => x"ea",
          4254 => x"f8",
          4255 => x"9e",
          4256 => x"05",
          4257 => x"54",
          4258 => x"38",
          4259 => x"70",
          4260 => x"54",
          4261 => x"8e",
          4262 => x"83",
          4263 => x"88",
          4264 => x"83",
          4265 => x"83",
          4266 => x"06",
          4267 => x"80",
          4268 => x"38",
          4269 => x"51",
          4270 => x"81",
          4271 => x"56",
          4272 => x"0a",
          4273 => x"05",
          4274 => x"3f",
          4275 => x"0b",
          4276 => x"80",
          4277 => x"7a",
          4278 => x"3f",
          4279 => x"9c",
          4280 => x"d1",
          4281 => x"81",
          4282 => x"34",
          4283 => x"80",
          4284 => x"b0",
          4285 => x"54",
          4286 => x"52",
          4287 => x"05",
          4288 => x"3f",
          4289 => x"08",
          4290 => x"c8",
          4291 => x"38",
          4292 => x"82",
          4293 => x"b2",
          4294 => x"84",
          4295 => x"06",
          4296 => x"73",
          4297 => x"38",
          4298 => x"ad",
          4299 => x"2a",
          4300 => x"51",
          4301 => x"2e",
          4302 => x"81",
          4303 => x"80",
          4304 => x"87",
          4305 => x"39",
          4306 => x"51",
          4307 => x"81",
          4308 => x"7b",
          4309 => x"12",
          4310 => x"81",
          4311 => x"81",
          4312 => x"83",
          4313 => x"06",
          4314 => x"80",
          4315 => x"77",
          4316 => x"58",
          4317 => x"08",
          4318 => x"63",
          4319 => x"63",
          4320 => x"57",
          4321 => x"81",
          4322 => x"81",
          4323 => x"88",
          4324 => x"9c",
          4325 => x"d2",
          4326 => x"f8",
          4327 => x"f8",
          4328 => x"1b",
          4329 => x"0c",
          4330 => x"22",
          4331 => x"77",
          4332 => x"80",
          4333 => x"34",
          4334 => x"1a",
          4335 => x"94",
          4336 => x"85",
          4337 => x"06",
          4338 => x"80",
          4339 => x"38",
          4340 => x"08",
          4341 => x"84",
          4342 => x"c8",
          4343 => x"0c",
          4344 => x"70",
          4345 => x"52",
          4346 => x"39",
          4347 => x"51",
          4348 => x"81",
          4349 => x"57",
          4350 => x"08",
          4351 => x"38",
          4352 => x"f8",
          4353 => x"2e",
          4354 => x"83",
          4355 => x"75",
          4356 => x"74",
          4357 => x"07",
          4358 => x"54",
          4359 => x"8a",
          4360 => x"75",
          4361 => x"73",
          4362 => x"98",
          4363 => x"a9",
          4364 => x"ff",
          4365 => x"80",
          4366 => x"76",
          4367 => x"d6",
          4368 => x"f8",
          4369 => x"38",
          4370 => x"39",
          4371 => x"81",
          4372 => x"05",
          4373 => x"84",
          4374 => x"0c",
          4375 => x"81",
          4376 => x"97",
          4377 => x"f2",
          4378 => x"63",
          4379 => x"40",
          4380 => x"7e",
          4381 => x"fc",
          4382 => x"51",
          4383 => x"81",
          4384 => x"55",
          4385 => x"08",
          4386 => x"19",
          4387 => x"80",
          4388 => x"74",
          4389 => x"39",
          4390 => x"81",
          4391 => x"56",
          4392 => x"82",
          4393 => x"39",
          4394 => x"1a",
          4395 => x"82",
          4396 => x"0b",
          4397 => x"81",
          4398 => x"39",
          4399 => x"94",
          4400 => x"55",
          4401 => x"83",
          4402 => x"7b",
          4403 => x"89",
          4404 => x"08",
          4405 => x"06",
          4406 => x"81",
          4407 => x"8a",
          4408 => x"05",
          4409 => x"06",
          4410 => x"a8",
          4411 => x"38",
          4412 => x"55",
          4413 => x"19",
          4414 => x"51",
          4415 => x"81",
          4416 => x"55",
          4417 => x"ff",
          4418 => x"ff",
          4419 => x"38",
          4420 => x"0c",
          4421 => x"52",
          4422 => x"cb",
          4423 => x"c8",
          4424 => x"ff",
          4425 => x"f8",
          4426 => x"7c",
          4427 => x"57",
          4428 => x"80",
          4429 => x"1a",
          4430 => x"22",
          4431 => x"75",
          4432 => x"38",
          4433 => x"58",
          4434 => x"53",
          4435 => x"1b",
          4436 => x"88",
          4437 => x"c8",
          4438 => x"38",
          4439 => x"33",
          4440 => x"80",
          4441 => x"b0",
          4442 => x"31",
          4443 => x"27",
          4444 => x"80",
          4445 => x"52",
          4446 => x"77",
          4447 => x"7d",
          4448 => x"e0",
          4449 => x"2b",
          4450 => x"76",
          4451 => x"94",
          4452 => x"ff",
          4453 => x"71",
          4454 => x"7b",
          4455 => x"38",
          4456 => x"19",
          4457 => x"51",
          4458 => x"81",
          4459 => x"fe",
          4460 => x"53",
          4461 => x"83",
          4462 => x"b4",
          4463 => x"51",
          4464 => x"7b",
          4465 => x"08",
          4466 => x"76",
          4467 => x"08",
          4468 => x"0c",
          4469 => x"f3",
          4470 => x"75",
          4471 => x"0c",
          4472 => x"04",
          4473 => x"60",
          4474 => x"40",
          4475 => x"80",
          4476 => x"3d",
          4477 => x"77",
          4478 => x"3f",
          4479 => x"08",
          4480 => x"c8",
          4481 => x"91",
          4482 => x"74",
          4483 => x"38",
          4484 => x"b8",
          4485 => x"33",
          4486 => x"70",
          4487 => x"56",
          4488 => x"74",
          4489 => x"a4",
          4490 => x"82",
          4491 => x"34",
          4492 => x"98",
          4493 => x"91",
          4494 => x"56",
          4495 => x"94",
          4496 => x"11",
          4497 => x"76",
          4498 => x"75",
          4499 => x"80",
          4500 => x"38",
          4501 => x"70",
          4502 => x"56",
          4503 => x"fd",
          4504 => x"11",
          4505 => x"77",
          4506 => x"5c",
          4507 => x"38",
          4508 => x"88",
          4509 => x"74",
          4510 => x"52",
          4511 => x"18",
          4512 => x"51",
          4513 => x"81",
          4514 => x"55",
          4515 => x"08",
          4516 => x"ab",
          4517 => x"2e",
          4518 => x"74",
          4519 => x"95",
          4520 => x"19",
          4521 => x"08",
          4522 => x"88",
          4523 => x"55",
          4524 => x"9c",
          4525 => x"09",
          4526 => x"38",
          4527 => x"c1",
          4528 => x"c8",
          4529 => x"38",
          4530 => x"52",
          4531 => x"97",
          4532 => x"c8",
          4533 => x"fe",
          4534 => x"f8",
          4535 => x"7c",
          4536 => x"57",
          4537 => x"80",
          4538 => x"1b",
          4539 => x"22",
          4540 => x"75",
          4541 => x"38",
          4542 => x"59",
          4543 => x"53",
          4544 => x"1a",
          4545 => x"be",
          4546 => x"c8",
          4547 => x"38",
          4548 => x"08",
          4549 => x"56",
          4550 => x"9b",
          4551 => x"53",
          4552 => x"77",
          4553 => x"7d",
          4554 => x"16",
          4555 => x"3f",
          4556 => x"0b",
          4557 => x"78",
          4558 => x"80",
          4559 => x"18",
          4560 => x"08",
          4561 => x"7e",
          4562 => x"3f",
          4563 => x"08",
          4564 => x"7e",
          4565 => x"0c",
          4566 => x"19",
          4567 => x"08",
          4568 => x"84",
          4569 => x"57",
          4570 => x"27",
          4571 => x"56",
          4572 => x"52",
          4573 => x"f9",
          4574 => x"c8",
          4575 => x"38",
          4576 => x"52",
          4577 => x"83",
          4578 => x"b4",
          4579 => x"d4",
          4580 => x"81",
          4581 => x"34",
          4582 => x"7e",
          4583 => x"0c",
          4584 => x"1a",
          4585 => x"94",
          4586 => x"1b",
          4587 => x"5e",
          4588 => x"27",
          4589 => x"55",
          4590 => x"0c",
          4591 => x"90",
          4592 => x"c0",
          4593 => x"90",
          4594 => x"56",
          4595 => x"c8",
          4596 => x"0d",
          4597 => x"0d",
          4598 => x"fc",
          4599 => x"52",
          4600 => x"3f",
          4601 => x"08",
          4602 => x"c8",
          4603 => x"38",
          4604 => x"70",
          4605 => x"81",
          4606 => x"55",
          4607 => x"80",
          4608 => x"16",
          4609 => x"51",
          4610 => x"81",
          4611 => x"57",
          4612 => x"08",
          4613 => x"a4",
          4614 => x"11",
          4615 => x"55",
          4616 => x"16",
          4617 => x"08",
          4618 => x"75",
          4619 => x"e8",
          4620 => x"08",
          4621 => x"51",
          4622 => x"82",
          4623 => x"52",
          4624 => x"c9",
          4625 => x"52",
          4626 => x"c9",
          4627 => x"54",
          4628 => x"15",
          4629 => x"cc",
          4630 => x"f8",
          4631 => x"17",
          4632 => x"06",
          4633 => x"90",
          4634 => x"81",
          4635 => x"8a",
          4636 => x"fc",
          4637 => x"70",
          4638 => x"d9",
          4639 => x"c8",
          4640 => x"f8",
          4641 => x"38",
          4642 => x"05",
          4643 => x"f1",
          4644 => x"f8",
          4645 => x"81",
          4646 => x"87",
          4647 => x"c8",
          4648 => x"72",
          4649 => x"0c",
          4650 => x"04",
          4651 => x"84",
          4652 => x"e4",
          4653 => x"80",
          4654 => x"c8",
          4655 => x"38",
          4656 => x"08",
          4657 => x"34",
          4658 => x"81",
          4659 => x"83",
          4660 => x"ef",
          4661 => x"53",
          4662 => x"05",
          4663 => x"51",
          4664 => x"81",
          4665 => x"55",
          4666 => x"08",
          4667 => x"76",
          4668 => x"93",
          4669 => x"51",
          4670 => x"81",
          4671 => x"55",
          4672 => x"08",
          4673 => x"80",
          4674 => x"70",
          4675 => x"56",
          4676 => x"89",
          4677 => x"94",
          4678 => x"b2",
          4679 => x"05",
          4680 => x"2a",
          4681 => x"51",
          4682 => x"80",
          4683 => x"76",
          4684 => x"52",
          4685 => x"3f",
          4686 => x"08",
          4687 => x"8e",
          4688 => x"c8",
          4689 => x"09",
          4690 => x"38",
          4691 => x"81",
          4692 => x"93",
          4693 => x"e4",
          4694 => x"6f",
          4695 => x"7a",
          4696 => x"9e",
          4697 => x"05",
          4698 => x"51",
          4699 => x"81",
          4700 => x"57",
          4701 => x"08",
          4702 => x"7b",
          4703 => x"94",
          4704 => x"55",
          4705 => x"73",
          4706 => x"ed",
          4707 => x"93",
          4708 => x"55",
          4709 => x"81",
          4710 => x"57",
          4711 => x"08",
          4712 => x"68",
          4713 => x"c9",
          4714 => x"f8",
          4715 => x"81",
          4716 => x"82",
          4717 => x"52",
          4718 => x"a3",
          4719 => x"c8",
          4720 => x"52",
          4721 => x"b8",
          4722 => x"c8",
          4723 => x"f8",
          4724 => x"a2",
          4725 => x"74",
          4726 => x"3f",
          4727 => x"08",
          4728 => x"c8",
          4729 => x"69",
          4730 => x"d9",
          4731 => x"81",
          4732 => x"2e",
          4733 => x"52",
          4734 => x"cf",
          4735 => x"c8",
          4736 => x"f8",
          4737 => x"2e",
          4738 => x"84",
          4739 => x"06",
          4740 => x"57",
          4741 => x"76",
          4742 => x"9e",
          4743 => x"05",
          4744 => x"dc",
          4745 => x"90",
          4746 => x"81",
          4747 => x"56",
          4748 => x"80",
          4749 => x"02",
          4750 => x"81",
          4751 => x"70",
          4752 => x"56",
          4753 => x"81",
          4754 => x"78",
          4755 => x"38",
          4756 => x"99",
          4757 => x"81",
          4758 => x"18",
          4759 => x"18",
          4760 => x"58",
          4761 => x"33",
          4762 => x"ee",
          4763 => x"6f",
          4764 => x"af",
          4765 => x"8d",
          4766 => x"2e",
          4767 => x"8a",
          4768 => x"6f",
          4769 => x"af",
          4770 => x"0b",
          4771 => x"33",
          4772 => x"81",
          4773 => x"70",
          4774 => x"52",
          4775 => x"56",
          4776 => x"8d",
          4777 => x"70",
          4778 => x"51",
          4779 => x"f5",
          4780 => x"54",
          4781 => x"a7",
          4782 => x"74",
          4783 => x"38",
          4784 => x"73",
          4785 => x"81",
          4786 => x"81",
          4787 => x"39",
          4788 => x"81",
          4789 => x"74",
          4790 => x"81",
          4791 => x"91",
          4792 => x"6e",
          4793 => x"59",
          4794 => x"7a",
          4795 => x"5c",
          4796 => x"26",
          4797 => x"7a",
          4798 => x"f8",
          4799 => x"3d",
          4800 => x"3d",
          4801 => x"8d",
          4802 => x"54",
          4803 => x"55",
          4804 => x"81",
          4805 => x"53",
          4806 => x"08",
          4807 => x"91",
          4808 => x"72",
          4809 => x"8c",
          4810 => x"73",
          4811 => x"38",
          4812 => x"70",
          4813 => x"81",
          4814 => x"57",
          4815 => x"73",
          4816 => x"08",
          4817 => x"94",
          4818 => x"75",
          4819 => x"97",
          4820 => x"11",
          4821 => x"2b",
          4822 => x"73",
          4823 => x"38",
          4824 => x"16",
          4825 => x"c3",
          4826 => x"c8",
          4827 => x"78",
          4828 => x"55",
          4829 => x"b3",
          4830 => x"c8",
          4831 => x"96",
          4832 => x"70",
          4833 => x"94",
          4834 => x"71",
          4835 => x"08",
          4836 => x"53",
          4837 => x"15",
          4838 => x"a6",
          4839 => x"74",
          4840 => x"3f",
          4841 => x"08",
          4842 => x"c8",
          4843 => x"81",
          4844 => x"f8",
          4845 => x"2e",
          4846 => x"81",
          4847 => x"88",
          4848 => x"98",
          4849 => x"80",
          4850 => x"38",
          4851 => x"80",
          4852 => x"77",
          4853 => x"08",
          4854 => x"0c",
          4855 => x"70",
          4856 => x"81",
          4857 => x"5a",
          4858 => x"2e",
          4859 => x"52",
          4860 => x"f9",
          4861 => x"c8",
          4862 => x"f8",
          4863 => x"38",
          4864 => x"08",
          4865 => x"73",
          4866 => x"c7",
          4867 => x"f8",
          4868 => x"73",
          4869 => x"38",
          4870 => x"af",
          4871 => x"73",
          4872 => x"27",
          4873 => x"98",
          4874 => x"a0",
          4875 => x"08",
          4876 => x"0c",
          4877 => x"06",
          4878 => x"2e",
          4879 => x"52",
          4880 => x"a3",
          4881 => x"c8",
          4882 => x"82",
          4883 => x"34",
          4884 => x"c4",
          4885 => x"91",
          4886 => x"53",
          4887 => x"89",
          4888 => x"c8",
          4889 => x"94",
          4890 => x"8c",
          4891 => x"27",
          4892 => x"8c",
          4893 => x"15",
          4894 => x"07",
          4895 => x"16",
          4896 => x"ff",
          4897 => x"80",
          4898 => x"77",
          4899 => x"2e",
          4900 => x"9c",
          4901 => x"53",
          4902 => x"c8",
          4903 => x"0d",
          4904 => x"0d",
          4905 => x"54",
          4906 => x"81",
          4907 => x"53",
          4908 => x"05",
          4909 => x"84",
          4910 => x"e7",
          4911 => x"c8",
          4912 => x"f8",
          4913 => x"ea",
          4914 => x"0c",
          4915 => x"51",
          4916 => x"81",
          4917 => x"55",
          4918 => x"08",
          4919 => x"ab",
          4920 => x"98",
          4921 => x"80",
          4922 => x"38",
          4923 => x"70",
          4924 => x"81",
          4925 => x"57",
          4926 => x"ad",
          4927 => x"08",
          4928 => x"d3",
          4929 => x"f8",
          4930 => x"17",
          4931 => x"86",
          4932 => x"17",
          4933 => x"75",
          4934 => x"3f",
          4935 => x"08",
          4936 => x"2e",
          4937 => x"85",
          4938 => x"86",
          4939 => x"2e",
          4940 => x"76",
          4941 => x"73",
          4942 => x"0c",
          4943 => x"04",
          4944 => x"76",
          4945 => x"05",
          4946 => x"53",
          4947 => x"81",
          4948 => x"87",
          4949 => x"c8",
          4950 => x"86",
          4951 => x"fb",
          4952 => x"79",
          4953 => x"05",
          4954 => x"56",
          4955 => x"3f",
          4956 => x"08",
          4957 => x"c8",
          4958 => x"38",
          4959 => x"81",
          4960 => x"52",
          4961 => x"f8",
          4962 => x"c8",
          4963 => x"ca",
          4964 => x"c8",
          4965 => x"51",
          4966 => x"81",
          4967 => x"53",
          4968 => x"08",
          4969 => x"81",
          4970 => x"80",
          4971 => x"81",
          4972 => x"a6",
          4973 => x"73",
          4974 => x"3f",
          4975 => x"51",
          4976 => x"81",
          4977 => x"84",
          4978 => x"70",
          4979 => x"2c",
          4980 => x"c8",
          4981 => x"51",
          4982 => x"81",
          4983 => x"87",
          4984 => x"ee",
          4985 => x"57",
          4986 => x"3d",
          4987 => x"3d",
          4988 => x"af",
          4989 => x"c8",
          4990 => x"f8",
          4991 => x"38",
          4992 => x"51",
          4993 => x"81",
          4994 => x"55",
          4995 => x"08",
          4996 => x"80",
          4997 => x"70",
          4998 => x"58",
          4999 => x"85",
          5000 => x"8d",
          5001 => x"2e",
          5002 => x"52",
          5003 => x"be",
          5004 => x"f8",
          5005 => x"3d",
          5006 => x"3d",
          5007 => x"55",
          5008 => x"92",
          5009 => x"52",
          5010 => x"de",
          5011 => x"f8",
          5012 => x"81",
          5013 => x"82",
          5014 => x"74",
          5015 => x"98",
          5016 => x"11",
          5017 => x"59",
          5018 => x"75",
          5019 => x"38",
          5020 => x"81",
          5021 => x"5b",
          5022 => x"82",
          5023 => x"39",
          5024 => x"08",
          5025 => x"59",
          5026 => x"09",
          5027 => x"38",
          5028 => x"57",
          5029 => x"3d",
          5030 => x"c1",
          5031 => x"f8",
          5032 => x"2e",
          5033 => x"f8",
          5034 => x"2e",
          5035 => x"f8",
          5036 => x"70",
          5037 => x"08",
          5038 => x"7a",
          5039 => x"7f",
          5040 => x"54",
          5041 => x"77",
          5042 => x"80",
          5043 => x"15",
          5044 => x"c8",
          5045 => x"75",
          5046 => x"52",
          5047 => x"52",
          5048 => x"8d",
          5049 => x"c8",
          5050 => x"f8",
          5051 => x"d6",
          5052 => x"33",
          5053 => x"1a",
          5054 => x"54",
          5055 => x"09",
          5056 => x"38",
          5057 => x"ff",
          5058 => x"81",
          5059 => x"83",
          5060 => x"70",
          5061 => x"25",
          5062 => x"59",
          5063 => x"9b",
          5064 => x"51",
          5065 => x"3f",
          5066 => x"08",
          5067 => x"70",
          5068 => x"25",
          5069 => x"59",
          5070 => x"75",
          5071 => x"7a",
          5072 => x"ff",
          5073 => x"7c",
          5074 => x"90",
          5075 => x"11",
          5076 => x"56",
          5077 => x"15",
          5078 => x"f8",
          5079 => x"3d",
          5080 => x"3d",
          5081 => x"3d",
          5082 => x"70",
          5083 => x"dd",
          5084 => x"c8",
          5085 => x"f8",
          5086 => x"a8",
          5087 => x"33",
          5088 => x"a0",
          5089 => x"33",
          5090 => x"70",
          5091 => x"55",
          5092 => x"73",
          5093 => x"8e",
          5094 => x"08",
          5095 => x"18",
          5096 => x"80",
          5097 => x"38",
          5098 => x"08",
          5099 => x"08",
          5100 => x"c4",
          5101 => x"f8",
          5102 => x"88",
          5103 => x"80",
          5104 => x"17",
          5105 => x"51",
          5106 => x"3f",
          5107 => x"08",
          5108 => x"81",
          5109 => x"81",
          5110 => x"c8",
          5111 => x"09",
          5112 => x"38",
          5113 => x"39",
          5114 => x"77",
          5115 => x"c8",
          5116 => x"08",
          5117 => x"98",
          5118 => x"81",
          5119 => x"52",
          5120 => x"bd",
          5121 => x"c8",
          5122 => x"17",
          5123 => x"0c",
          5124 => x"80",
          5125 => x"73",
          5126 => x"75",
          5127 => x"38",
          5128 => x"34",
          5129 => x"81",
          5130 => x"89",
          5131 => x"e2",
          5132 => x"53",
          5133 => x"a4",
          5134 => x"3d",
          5135 => x"3f",
          5136 => x"08",
          5137 => x"c8",
          5138 => x"38",
          5139 => x"3d",
          5140 => x"3d",
          5141 => x"d1",
          5142 => x"f8",
          5143 => x"81",
          5144 => x"81",
          5145 => x"80",
          5146 => x"70",
          5147 => x"81",
          5148 => x"56",
          5149 => x"81",
          5150 => x"98",
          5151 => x"74",
          5152 => x"38",
          5153 => x"05",
          5154 => x"06",
          5155 => x"55",
          5156 => x"38",
          5157 => x"51",
          5158 => x"81",
          5159 => x"74",
          5160 => x"81",
          5161 => x"56",
          5162 => x"80",
          5163 => x"54",
          5164 => x"08",
          5165 => x"2e",
          5166 => x"73",
          5167 => x"c8",
          5168 => x"52",
          5169 => x"52",
          5170 => x"3f",
          5171 => x"08",
          5172 => x"c8",
          5173 => x"38",
          5174 => x"08",
          5175 => x"cc",
          5176 => x"f8",
          5177 => x"81",
          5178 => x"86",
          5179 => x"80",
          5180 => x"f8",
          5181 => x"2e",
          5182 => x"f8",
          5183 => x"c0",
          5184 => x"ce",
          5185 => x"f8",
          5186 => x"f8",
          5187 => x"70",
          5188 => x"08",
          5189 => x"51",
          5190 => x"80",
          5191 => x"73",
          5192 => x"38",
          5193 => x"52",
          5194 => x"95",
          5195 => x"c8",
          5196 => x"8c",
          5197 => x"ff",
          5198 => x"81",
          5199 => x"55",
          5200 => x"c8",
          5201 => x"0d",
          5202 => x"0d",
          5203 => x"3d",
          5204 => x"9a",
          5205 => x"cb",
          5206 => x"c8",
          5207 => x"f8",
          5208 => x"b0",
          5209 => x"69",
          5210 => x"70",
          5211 => x"97",
          5212 => x"c8",
          5213 => x"f8",
          5214 => x"38",
          5215 => x"94",
          5216 => x"c8",
          5217 => x"09",
          5218 => x"88",
          5219 => x"df",
          5220 => x"85",
          5221 => x"51",
          5222 => x"74",
          5223 => x"78",
          5224 => x"8a",
          5225 => x"57",
          5226 => x"81",
          5227 => x"75",
          5228 => x"f8",
          5229 => x"38",
          5230 => x"f8",
          5231 => x"2e",
          5232 => x"83",
          5233 => x"81",
          5234 => x"ff",
          5235 => x"06",
          5236 => x"54",
          5237 => x"73",
          5238 => x"81",
          5239 => x"52",
          5240 => x"a4",
          5241 => x"c8",
          5242 => x"f8",
          5243 => x"9a",
          5244 => x"a0",
          5245 => x"51",
          5246 => x"3f",
          5247 => x"0b",
          5248 => x"78",
          5249 => x"bf",
          5250 => x"88",
          5251 => x"80",
          5252 => x"ff",
          5253 => x"75",
          5254 => x"11",
          5255 => x"f8",
          5256 => x"78",
          5257 => x"80",
          5258 => x"ff",
          5259 => x"78",
          5260 => x"80",
          5261 => x"7f",
          5262 => x"d4",
          5263 => x"c9",
          5264 => x"54",
          5265 => x"15",
          5266 => x"cb",
          5267 => x"f8",
          5268 => x"81",
          5269 => x"b2",
          5270 => x"b2",
          5271 => x"96",
          5272 => x"b5",
          5273 => x"53",
          5274 => x"51",
          5275 => x"64",
          5276 => x"8b",
          5277 => x"54",
          5278 => x"15",
          5279 => x"ff",
          5280 => x"81",
          5281 => x"54",
          5282 => x"53",
          5283 => x"51",
          5284 => x"3f",
          5285 => x"c8",
          5286 => x"0d",
          5287 => x"0d",
          5288 => x"05",
          5289 => x"3f",
          5290 => x"3d",
          5291 => x"52",
          5292 => x"d5",
          5293 => x"f8",
          5294 => x"81",
          5295 => x"82",
          5296 => x"4d",
          5297 => x"52",
          5298 => x"52",
          5299 => x"3f",
          5300 => x"08",
          5301 => x"c8",
          5302 => x"38",
          5303 => x"05",
          5304 => x"06",
          5305 => x"73",
          5306 => x"a0",
          5307 => x"08",
          5308 => x"ff",
          5309 => x"ff",
          5310 => x"ac",
          5311 => x"92",
          5312 => x"54",
          5313 => x"3f",
          5314 => x"52",
          5315 => x"f7",
          5316 => x"c8",
          5317 => x"f8",
          5318 => x"38",
          5319 => x"09",
          5320 => x"38",
          5321 => x"08",
          5322 => x"88",
          5323 => x"39",
          5324 => x"08",
          5325 => x"81",
          5326 => x"38",
          5327 => x"b1",
          5328 => x"c8",
          5329 => x"f8",
          5330 => x"c8",
          5331 => x"93",
          5332 => x"ff",
          5333 => x"8d",
          5334 => x"b4",
          5335 => x"af",
          5336 => x"17",
          5337 => x"33",
          5338 => x"70",
          5339 => x"55",
          5340 => x"38",
          5341 => x"54",
          5342 => x"34",
          5343 => x"0b",
          5344 => x"8b",
          5345 => x"84",
          5346 => x"06",
          5347 => x"73",
          5348 => x"e5",
          5349 => x"2e",
          5350 => x"75",
          5351 => x"c6",
          5352 => x"f8",
          5353 => x"78",
          5354 => x"bb",
          5355 => x"81",
          5356 => x"80",
          5357 => x"38",
          5358 => x"08",
          5359 => x"ff",
          5360 => x"81",
          5361 => x"79",
          5362 => x"58",
          5363 => x"f8",
          5364 => x"c0",
          5365 => x"33",
          5366 => x"2e",
          5367 => x"99",
          5368 => x"75",
          5369 => x"c6",
          5370 => x"54",
          5371 => x"15",
          5372 => x"81",
          5373 => x"9c",
          5374 => x"c8",
          5375 => x"f8",
          5376 => x"81",
          5377 => x"8c",
          5378 => x"ff",
          5379 => x"81",
          5380 => x"55",
          5381 => x"c8",
          5382 => x"0d",
          5383 => x"0d",
          5384 => x"05",
          5385 => x"05",
          5386 => x"33",
          5387 => x"53",
          5388 => x"05",
          5389 => x"51",
          5390 => x"81",
          5391 => x"55",
          5392 => x"08",
          5393 => x"78",
          5394 => x"95",
          5395 => x"51",
          5396 => x"81",
          5397 => x"55",
          5398 => x"08",
          5399 => x"80",
          5400 => x"81",
          5401 => x"86",
          5402 => x"38",
          5403 => x"61",
          5404 => x"12",
          5405 => x"7a",
          5406 => x"51",
          5407 => x"74",
          5408 => x"78",
          5409 => x"83",
          5410 => x"51",
          5411 => x"3f",
          5412 => x"08",
          5413 => x"f8",
          5414 => x"3d",
          5415 => x"3d",
          5416 => x"82",
          5417 => x"d0",
          5418 => x"3d",
          5419 => x"3f",
          5420 => x"08",
          5421 => x"c8",
          5422 => x"38",
          5423 => x"52",
          5424 => x"05",
          5425 => x"3f",
          5426 => x"08",
          5427 => x"c8",
          5428 => x"02",
          5429 => x"33",
          5430 => x"54",
          5431 => x"a6",
          5432 => x"22",
          5433 => x"71",
          5434 => x"53",
          5435 => x"51",
          5436 => x"3f",
          5437 => x"0b",
          5438 => x"76",
          5439 => x"b8",
          5440 => x"c8",
          5441 => x"81",
          5442 => x"93",
          5443 => x"ea",
          5444 => x"6b",
          5445 => x"53",
          5446 => x"05",
          5447 => x"51",
          5448 => x"81",
          5449 => x"81",
          5450 => x"30",
          5451 => x"c8",
          5452 => x"25",
          5453 => x"79",
          5454 => x"85",
          5455 => x"75",
          5456 => x"73",
          5457 => x"f9",
          5458 => x"80",
          5459 => x"8d",
          5460 => x"54",
          5461 => x"3f",
          5462 => x"08",
          5463 => x"c8",
          5464 => x"38",
          5465 => x"51",
          5466 => x"81",
          5467 => x"57",
          5468 => x"08",
          5469 => x"f8",
          5470 => x"f8",
          5471 => x"5b",
          5472 => x"18",
          5473 => x"18",
          5474 => x"74",
          5475 => x"81",
          5476 => x"78",
          5477 => x"8b",
          5478 => x"54",
          5479 => x"75",
          5480 => x"38",
          5481 => x"1b",
          5482 => x"55",
          5483 => x"2e",
          5484 => x"39",
          5485 => x"09",
          5486 => x"38",
          5487 => x"80",
          5488 => x"70",
          5489 => x"25",
          5490 => x"80",
          5491 => x"38",
          5492 => x"bc",
          5493 => x"11",
          5494 => x"ff",
          5495 => x"81",
          5496 => x"57",
          5497 => x"08",
          5498 => x"70",
          5499 => x"80",
          5500 => x"83",
          5501 => x"80",
          5502 => x"84",
          5503 => x"a7",
          5504 => x"b4",
          5505 => x"ad",
          5506 => x"f8",
          5507 => x"0c",
          5508 => x"c8",
          5509 => x"0d",
          5510 => x"0d",
          5511 => x"3d",
          5512 => x"52",
          5513 => x"ce",
          5514 => x"f8",
          5515 => x"f8",
          5516 => x"54",
          5517 => x"08",
          5518 => x"8b",
          5519 => x"8b",
          5520 => x"59",
          5521 => x"3f",
          5522 => x"33",
          5523 => x"06",
          5524 => x"57",
          5525 => x"81",
          5526 => x"58",
          5527 => x"06",
          5528 => x"4e",
          5529 => x"ff",
          5530 => x"81",
          5531 => x"80",
          5532 => x"6c",
          5533 => x"53",
          5534 => x"ae",
          5535 => x"f8",
          5536 => x"2e",
          5537 => x"88",
          5538 => x"6d",
          5539 => x"55",
          5540 => x"f8",
          5541 => x"ff",
          5542 => x"83",
          5543 => x"51",
          5544 => x"26",
          5545 => x"15",
          5546 => x"ff",
          5547 => x"80",
          5548 => x"87",
          5549 => x"d8",
          5550 => x"74",
          5551 => x"38",
          5552 => x"e7",
          5553 => x"ae",
          5554 => x"f8",
          5555 => x"38",
          5556 => x"27",
          5557 => x"89",
          5558 => x"8b",
          5559 => x"27",
          5560 => x"55",
          5561 => x"81",
          5562 => x"8f",
          5563 => x"2a",
          5564 => x"70",
          5565 => x"34",
          5566 => x"74",
          5567 => x"05",
          5568 => x"17",
          5569 => x"70",
          5570 => x"52",
          5571 => x"73",
          5572 => x"c8",
          5573 => x"33",
          5574 => x"73",
          5575 => x"81",
          5576 => x"80",
          5577 => x"02",
          5578 => x"76",
          5579 => x"51",
          5580 => x"2e",
          5581 => x"87",
          5582 => x"57",
          5583 => x"79",
          5584 => x"80",
          5585 => x"70",
          5586 => x"ba",
          5587 => x"f8",
          5588 => x"81",
          5589 => x"80",
          5590 => x"52",
          5591 => x"bf",
          5592 => x"f8",
          5593 => x"81",
          5594 => x"8d",
          5595 => x"c4",
          5596 => x"e5",
          5597 => x"c6",
          5598 => x"c8",
          5599 => x"09",
          5600 => x"cc",
          5601 => x"76",
          5602 => x"c4",
          5603 => x"74",
          5604 => x"b0",
          5605 => x"c8",
          5606 => x"f8",
          5607 => x"38",
          5608 => x"f8",
          5609 => x"67",
          5610 => x"db",
          5611 => x"88",
          5612 => x"34",
          5613 => x"52",
          5614 => x"ab",
          5615 => x"54",
          5616 => x"15",
          5617 => x"ff",
          5618 => x"81",
          5619 => x"54",
          5620 => x"81",
          5621 => x"9c",
          5622 => x"f2",
          5623 => x"62",
          5624 => x"80",
          5625 => x"93",
          5626 => x"55",
          5627 => x"5e",
          5628 => x"3f",
          5629 => x"08",
          5630 => x"c8",
          5631 => x"38",
          5632 => x"58",
          5633 => x"38",
          5634 => x"97",
          5635 => x"08",
          5636 => x"38",
          5637 => x"70",
          5638 => x"81",
          5639 => x"55",
          5640 => x"87",
          5641 => x"39",
          5642 => x"90",
          5643 => x"82",
          5644 => x"8a",
          5645 => x"89",
          5646 => x"7f",
          5647 => x"56",
          5648 => x"3f",
          5649 => x"06",
          5650 => x"72",
          5651 => x"81",
          5652 => x"05",
          5653 => x"7c",
          5654 => x"55",
          5655 => x"27",
          5656 => x"16",
          5657 => x"83",
          5658 => x"76",
          5659 => x"80",
          5660 => x"79",
          5661 => x"99",
          5662 => x"7f",
          5663 => x"14",
          5664 => x"83",
          5665 => x"81",
          5666 => x"81",
          5667 => x"38",
          5668 => x"08",
          5669 => x"95",
          5670 => x"c8",
          5671 => x"81",
          5672 => x"7b",
          5673 => x"06",
          5674 => x"39",
          5675 => x"56",
          5676 => x"09",
          5677 => x"b9",
          5678 => x"80",
          5679 => x"80",
          5680 => x"78",
          5681 => x"7a",
          5682 => x"38",
          5683 => x"73",
          5684 => x"81",
          5685 => x"ff",
          5686 => x"74",
          5687 => x"ff",
          5688 => x"81",
          5689 => x"58",
          5690 => x"08",
          5691 => x"74",
          5692 => x"16",
          5693 => x"73",
          5694 => x"39",
          5695 => x"7e",
          5696 => x"0c",
          5697 => x"2e",
          5698 => x"88",
          5699 => x"8c",
          5700 => x"1a",
          5701 => x"07",
          5702 => x"1b",
          5703 => x"08",
          5704 => x"16",
          5705 => x"75",
          5706 => x"38",
          5707 => x"90",
          5708 => x"15",
          5709 => x"54",
          5710 => x"34",
          5711 => x"81",
          5712 => x"90",
          5713 => x"e9",
          5714 => x"6d",
          5715 => x"80",
          5716 => x"9d",
          5717 => x"5c",
          5718 => x"3f",
          5719 => x"0b",
          5720 => x"08",
          5721 => x"38",
          5722 => x"08",
          5723 => x"f8",
          5724 => x"08",
          5725 => x"80",
          5726 => x"80",
          5727 => x"f8",
          5728 => x"ff",
          5729 => x"52",
          5730 => x"a0",
          5731 => x"f8",
          5732 => x"ff",
          5733 => x"06",
          5734 => x"56",
          5735 => x"38",
          5736 => x"70",
          5737 => x"55",
          5738 => x"8b",
          5739 => x"3d",
          5740 => x"83",
          5741 => x"ff",
          5742 => x"81",
          5743 => x"99",
          5744 => x"74",
          5745 => x"38",
          5746 => x"80",
          5747 => x"ff",
          5748 => x"55",
          5749 => x"83",
          5750 => x"78",
          5751 => x"38",
          5752 => x"26",
          5753 => x"81",
          5754 => x"8b",
          5755 => x"79",
          5756 => x"80",
          5757 => x"93",
          5758 => x"39",
          5759 => x"6e",
          5760 => x"89",
          5761 => x"48",
          5762 => x"83",
          5763 => x"61",
          5764 => x"25",
          5765 => x"55",
          5766 => x"8a",
          5767 => x"3d",
          5768 => x"81",
          5769 => x"ff",
          5770 => x"81",
          5771 => x"c8",
          5772 => x"38",
          5773 => x"70",
          5774 => x"f8",
          5775 => x"56",
          5776 => x"38",
          5777 => x"55",
          5778 => x"75",
          5779 => x"38",
          5780 => x"70",
          5781 => x"ff",
          5782 => x"83",
          5783 => x"78",
          5784 => x"89",
          5785 => x"81",
          5786 => x"06",
          5787 => x"80",
          5788 => x"77",
          5789 => x"74",
          5790 => x"8d",
          5791 => x"06",
          5792 => x"2e",
          5793 => x"77",
          5794 => x"93",
          5795 => x"74",
          5796 => x"cb",
          5797 => x"7d",
          5798 => x"81",
          5799 => x"38",
          5800 => x"66",
          5801 => x"81",
          5802 => x"fc",
          5803 => x"74",
          5804 => x"38",
          5805 => x"98",
          5806 => x"fc",
          5807 => x"82",
          5808 => x"57",
          5809 => x"80",
          5810 => x"76",
          5811 => x"38",
          5812 => x"51",
          5813 => x"3f",
          5814 => x"08",
          5815 => x"87",
          5816 => x"2a",
          5817 => x"5c",
          5818 => x"f8",
          5819 => x"80",
          5820 => x"44",
          5821 => x"0a",
          5822 => x"ec",
          5823 => x"39",
          5824 => x"66",
          5825 => x"81",
          5826 => x"ec",
          5827 => x"74",
          5828 => x"38",
          5829 => x"98",
          5830 => x"ec",
          5831 => x"82",
          5832 => x"57",
          5833 => x"80",
          5834 => x"76",
          5835 => x"38",
          5836 => x"51",
          5837 => x"3f",
          5838 => x"08",
          5839 => x"57",
          5840 => x"08",
          5841 => x"96",
          5842 => x"81",
          5843 => x"10",
          5844 => x"08",
          5845 => x"72",
          5846 => x"59",
          5847 => x"ff",
          5848 => x"5d",
          5849 => x"44",
          5850 => x"11",
          5851 => x"70",
          5852 => x"71",
          5853 => x"06",
          5854 => x"52",
          5855 => x"40",
          5856 => x"09",
          5857 => x"38",
          5858 => x"18",
          5859 => x"39",
          5860 => x"79",
          5861 => x"70",
          5862 => x"58",
          5863 => x"76",
          5864 => x"38",
          5865 => x"7d",
          5866 => x"70",
          5867 => x"55",
          5868 => x"3f",
          5869 => x"08",
          5870 => x"2e",
          5871 => x"9b",
          5872 => x"c8",
          5873 => x"f5",
          5874 => x"38",
          5875 => x"38",
          5876 => x"59",
          5877 => x"38",
          5878 => x"7d",
          5879 => x"81",
          5880 => x"38",
          5881 => x"0b",
          5882 => x"08",
          5883 => x"78",
          5884 => x"1a",
          5885 => x"c0",
          5886 => x"74",
          5887 => x"39",
          5888 => x"55",
          5889 => x"8f",
          5890 => x"fd",
          5891 => x"f8",
          5892 => x"f5",
          5893 => x"78",
          5894 => x"79",
          5895 => x"80",
          5896 => x"f1",
          5897 => x"39",
          5898 => x"81",
          5899 => x"06",
          5900 => x"55",
          5901 => x"27",
          5902 => x"81",
          5903 => x"56",
          5904 => x"38",
          5905 => x"80",
          5906 => x"ff",
          5907 => x"8b",
          5908 => x"94",
          5909 => x"ff",
          5910 => x"84",
          5911 => x"1b",
          5912 => x"b3",
          5913 => x"1c",
          5914 => x"ff",
          5915 => x"8e",
          5916 => x"a1",
          5917 => x"0b",
          5918 => x"7d",
          5919 => x"30",
          5920 => x"84",
          5921 => x"51",
          5922 => x"51",
          5923 => x"3f",
          5924 => x"83",
          5925 => x"90",
          5926 => x"ff",
          5927 => x"93",
          5928 => x"a0",
          5929 => x"39",
          5930 => x"1b",
          5931 => x"85",
          5932 => x"95",
          5933 => x"52",
          5934 => x"ff",
          5935 => x"81",
          5936 => x"1b",
          5937 => x"cf",
          5938 => x"9c",
          5939 => x"a0",
          5940 => x"83",
          5941 => x"06",
          5942 => x"82",
          5943 => x"52",
          5944 => x"51",
          5945 => x"3f",
          5946 => x"1b",
          5947 => x"c5",
          5948 => x"ac",
          5949 => x"a0",
          5950 => x"52",
          5951 => x"ff",
          5952 => x"86",
          5953 => x"51",
          5954 => x"3f",
          5955 => x"80",
          5956 => x"a9",
          5957 => x"1c",
          5958 => x"81",
          5959 => x"80",
          5960 => x"ae",
          5961 => x"b2",
          5962 => x"1b",
          5963 => x"85",
          5964 => x"ff",
          5965 => x"96",
          5966 => x"9f",
          5967 => x"80",
          5968 => x"34",
          5969 => x"1c",
          5970 => x"81",
          5971 => x"ab",
          5972 => x"a0",
          5973 => x"d4",
          5974 => x"fe",
          5975 => x"59",
          5976 => x"3f",
          5977 => x"53",
          5978 => x"51",
          5979 => x"3f",
          5980 => x"f8",
          5981 => x"e7",
          5982 => x"2e",
          5983 => x"80",
          5984 => x"54",
          5985 => x"53",
          5986 => x"51",
          5987 => x"3f",
          5988 => x"80",
          5989 => x"ff",
          5990 => x"84",
          5991 => x"d2",
          5992 => x"ff",
          5993 => x"86",
          5994 => x"f2",
          5995 => x"1b",
          5996 => x"81",
          5997 => x"52",
          5998 => x"51",
          5999 => x"3f",
          6000 => x"ec",
          6001 => x"9e",
          6002 => x"d4",
          6003 => x"51",
          6004 => x"3f",
          6005 => x"87",
          6006 => x"52",
          6007 => x"9a",
          6008 => x"54",
          6009 => x"7a",
          6010 => x"ff",
          6011 => x"65",
          6012 => x"7a",
          6013 => x"8f",
          6014 => x"80",
          6015 => x"2e",
          6016 => x"9a",
          6017 => x"7a",
          6018 => x"a9",
          6019 => x"84",
          6020 => x"9e",
          6021 => x"0a",
          6022 => x"51",
          6023 => x"ff",
          6024 => x"7d",
          6025 => x"38",
          6026 => x"52",
          6027 => x"9e",
          6028 => x"55",
          6029 => x"62",
          6030 => x"74",
          6031 => x"75",
          6032 => x"7e",
          6033 => x"fe",
          6034 => x"c8",
          6035 => x"38",
          6036 => x"81",
          6037 => x"52",
          6038 => x"9e",
          6039 => x"16",
          6040 => x"56",
          6041 => x"38",
          6042 => x"77",
          6043 => x"8d",
          6044 => x"7d",
          6045 => x"38",
          6046 => x"57",
          6047 => x"83",
          6048 => x"76",
          6049 => x"7a",
          6050 => x"ff",
          6051 => x"81",
          6052 => x"81",
          6053 => x"16",
          6054 => x"56",
          6055 => x"38",
          6056 => x"83",
          6057 => x"86",
          6058 => x"ff",
          6059 => x"38",
          6060 => x"82",
          6061 => x"81",
          6062 => x"06",
          6063 => x"fe",
          6064 => x"53",
          6065 => x"51",
          6066 => x"3f",
          6067 => x"52",
          6068 => x"9c",
          6069 => x"be",
          6070 => x"75",
          6071 => x"81",
          6072 => x"0b",
          6073 => x"77",
          6074 => x"75",
          6075 => x"60",
          6076 => x"80",
          6077 => x"75",
          6078 => x"af",
          6079 => x"85",
          6080 => x"f8",
          6081 => x"2a",
          6082 => x"75",
          6083 => x"81",
          6084 => x"87",
          6085 => x"52",
          6086 => x"51",
          6087 => x"3f",
          6088 => x"ca",
          6089 => x"9c",
          6090 => x"54",
          6091 => x"52",
          6092 => x"98",
          6093 => x"56",
          6094 => x"08",
          6095 => x"53",
          6096 => x"51",
          6097 => x"3f",
          6098 => x"f8",
          6099 => x"38",
          6100 => x"56",
          6101 => x"56",
          6102 => x"f8",
          6103 => x"75",
          6104 => x"0c",
          6105 => x"04",
          6106 => x"7d",
          6107 => x"80",
          6108 => x"05",
          6109 => x"76",
          6110 => x"38",
          6111 => x"11",
          6112 => x"53",
          6113 => x"79",
          6114 => x"3f",
          6115 => x"09",
          6116 => x"38",
          6117 => x"55",
          6118 => x"db",
          6119 => x"70",
          6120 => x"34",
          6121 => x"74",
          6122 => x"81",
          6123 => x"80",
          6124 => x"55",
          6125 => x"76",
          6126 => x"f8",
          6127 => x"3d",
          6128 => x"3d",
          6129 => x"84",
          6130 => x"33",
          6131 => x"8a",
          6132 => x"06",
          6133 => x"52",
          6134 => x"3f",
          6135 => x"56",
          6136 => x"be",
          6137 => x"08",
          6138 => x"05",
          6139 => x"75",
          6140 => x"56",
          6141 => x"a1",
          6142 => x"fc",
          6143 => x"53",
          6144 => x"76",
          6145 => x"dc",
          6146 => x"32",
          6147 => x"72",
          6148 => x"70",
          6149 => x"56",
          6150 => x"18",
          6151 => x"88",
          6152 => x"3d",
          6153 => x"3d",
          6154 => x"11",
          6155 => x"80",
          6156 => x"38",
          6157 => x"05",
          6158 => x"8c",
          6159 => x"08",
          6160 => x"3f",
          6161 => x"08",
          6162 => x"16",
          6163 => x"09",
          6164 => x"38",
          6165 => x"55",
          6166 => x"55",
          6167 => x"c8",
          6168 => x"0d",
          6169 => x"0d",
          6170 => x"cc",
          6171 => x"73",
          6172 => x"93",
          6173 => x"0c",
          6174 => x"04",
          6175 => x"02",
          6176 => x"33",
          6177 => x"3d",
          6178 => x"54",
          6179 => x"52",
          6180 => x"ae",
          6181 => x"ff",
          6182 => x"3d",
          6183 => x"3d",
          6184 => x"08",
          6185 => x"59",
          6186 => x"80",
          6187 => x"39",
          6188 => x"0c",
          6189 => x"54",
          6190 => x"74",
          6191 => x"a0",
          6192 => x"06",
          6193 => x"15",
          6194 => x"80",
          6195 => x"29",
          6196 => x"05",
          6197 => x"56",
          6198 => x"3f",
          6199 => x"08",
          6200 => x"08",
          6201 => x"76",
          6202 => x"fe",
          6203 => x"81",
          6204 => x"8b",
          6205 => x"33",
          6206 => x"2e",
          6207 => x"81",
          6208 => x"ff",
          6209 => x"98",
          6210 => x"38",
          6211 => x"81",
          6212 => x"8a",
          6213 => x"ff",
          6214 => x"52",
          6215 => x"81",
          6216 => x"84",
          6217 => x"80",
          6218 => x"08",
          6219 => x"b4",
          6220 => x"39",
          6221 => x"51",
          6222 => x"81",
          6223 => x"80",
          6224 => x"e9",
          6225 => x"eb",
          6226 => x"f8",
          6227 => x"39",
          6228 => x"51",
          6229 => x"81",
          6230 => x"80",
          6231 => x"ea",
          6232 => x"cf",
          6233 => x"c4",
          6234 => x"39",
          6235 => x"51",
          6236 => x"81",
          6237 => x"bb",
          6238 => x"90",
          6239 => x"81",
          6240 => x"af",
          6241 => x"d0",
          6242 => x"81",
          6243 => x"a3",
          6244 => x"84",
          6245 => x"81",
          6246 => x"97",
          6247 => x"b0",
          6248 => x"81",
          6249 => x"8b",
          6250 => x"e0",
          6251 => x"81",
          6252 => x"fe",
          6253 => x"83",
          6254 => x"fb",
          6255 => x"79",
          6256 => x"87",
          6257 => x"38",
          6258 => x"87",
          6259 => x"91",
          6260 => x"52",
          6261 => x"cf",
          6262 => x"f8",
          6263 => x"75",
          6264 => x"c7",
          6265 => x"c8",
          6266 => x"53",
          6267 => x"ec",
          6268 => x"f7",
          6269 => x"3d",
          6270 => x"3d",
          6271 => x"84",
          6272 => x"05",
          6273 => x"80",
          6274 => x"70",
          6275 => x"25",
          6276 => x"59",
          6277 => x"87",
          6278 => x"38",
          6279 => x"76",
          6280 => x"ff",
          6281 => x"93",
          6282 => x"80",
          6283 => x"76",
          6284 => x"70",
          6285 => x"bf",
          6286 => x"f8",
          6287 => x"81",
          6288 => x"b8",
          6289 => x"c8",
          6290 => x"98",
          6291 => x"f8",
          6292 => x"96",
          6293 => x"54",
          6294 => x"77",
          6295 => x"c4",
          6296 => x"f8",
          6297 => x"81",
          6298 => x"90",
          6299 => x"74",
          6300 => x"38",
          6301 => x"19",
          6302 => x"39",
          6303 => x"05",
          6304 => x"3f",
          6305 => x"78",
          6306 => x"7b",
          6307 => x"2a",
          6308 => x"57",
          6309 => x"80",
          6310 => x"81",
          6311 => x"87",
          6312 => x"08",
          6313 => x"fe",
          6314 => x"56",
          6315 => x"c8",
          6316 => x"0d",
          6317 => x"0d",
          6318 => x"05",
          6319 => x"57",
          6320 => x"80",
          6321 => x"79",
          6322 => x"3f",
          6323 => x"08",
          6324 => x"80",
          6325 => x"75",
          6326 => x"38",
          6327 => x"55",
          6328 => x"f8",
          6329 => x"52",
          6330 => x"2d",
          6331 => x"08",
          6332 => x"77",
          6333 => x"f8",
          6334 => x"3d",
          6335 => x"3d",
          6336 => x"63",
          6337 => x"80",
          6338 => x"73",
          6339 => x"41",
          6340 => x"5e",
          6341 => x"52",
          6342 => x"51",
          6343 => x"3f",
          6344 => x"51",
          6345 => x"3f",
          6346 => x"79",
          6347 => x"38",
          6348 => x"89",
          6349 => x"2e",
          6350 => x"c6",
          6351 => x"53",
          6352 => x"8e",
          6353 => x"52",
          6354 => x"51",
          6355 => x"3f",
          6356 => x"ed",
          6357 => x"ef",
          6358 => x"15",
          6359 => x"39",
          6360 => x"72",
          6361 => x"38",
          6362 => x"81",
          6363 => x"fe",
          6364 => x"89",
          6365 => x"bc",
          6366 => x"e8",
          6367 => x"55",
          6368 => x"18",
          6369 => x"27",
          6370 => x"33",
          6371 => x"c8",
          6372 => x"b4",
          6373 => x"81",
          6374 => x"fe",
          6375 => x"81",
          6376 => x"51",
          6377 => x"3f",
          6378 => x"81",
          6379 => x"fe",
          6380 => x"80",
          6381 => x"27",
          6382 => x"18",
          6383 => x"53",
          6384 => x"7a",
          6385 => x"81",
          6386 => x"9f",
          6387 => x"38",
          6388 => x"73",
          6389 => x"ff",
          6390 => x"72",
          6391 => x"38",
          6392 => x"26",
          6393 => x"51",
          6394 => x"51",
          6395 => x"3f",
          6396 => x"c1",
          6397 => x"d8",
          6398 => x"e8",
          6399 => x"79",
          6400 => x"fe",
          6401 => x"81",
          6402 => x"98",
          6403 => x"2c",
          6404 => x"a0",
          6405 => x"06",
          6406 => x"de",
          6407 => x"f8",
          6408 => x"2b",
          6409 => x"70",
          6410 => x"30",
          6411 => x"70",
          6412 => x"07",
          6413 => x"06",
          6414 => x"59",
          6415 => x"80",
          6416 => x"38",
          6417 => x"09",
          6418 => x"38",
          6419 => x"39",
          6420 => x"72",
          6421 => x"be",
          6422 => x"72",
          6423 => x"0c",
          6424 => x"04",
          6425 => x"02",
          6426 => x"81",
          6427 => x"81",
          6428 => x"55",
          6429 => x"3f",
          6430 => x"22",
          6431 => x"98",
          6432 => x"ec",
          6433 => x"f8",
          6434 => x"f9",
          6435 => x"ee",
          6436 => x"f2",
          6437 => x"80",
          6438 => x"fe",
          6439 => x"86",
          6440 => x"fe",
          6441 => x"c0",
          6442 => x"53",
          6443 => x"3f",
          6444 => x"d9",
          6445 => x"ee",
          6446 => x"db",
          6447 => x"51",
          6448 => x"3f",
          6449 => x"70",
          6450 => x"52",
          6451 => x"95",
          6452 => x"fe",
          6453 => x"81",
          6454 => x"fe",
          6455 => x"80",
          6456 => x"8d",
          6457 => x"2a",
          6458 => x"51",
          6459 => x"2e",
          6460 => x"51",
          6461 => x"3f",
          6462 => x"51",
          6463 => x"3f",
          6464 => x"d8",
          6465 => x"83",
          6466 => x"06",
          6467 => x"80",
          6468 => x"81",
          6469 => x"d9",
          6470 => x"d8",
          6471 => x"d1",
          6472 => x"fe",
          6473 => x"72",
          6474 => x"81",
          6475 => x"71",
          6476 => x"38",
          6477 => x"d8",
          6478 => x"ee",
          6479 => x"da",
          6480 => x"51",
          6481 => x"3f",
          6482 => x"70",
          6483 => x"52",
          6484 => x"95",
          6485 => x"fe",
          6486 => x"81",
          6487 => x"fe",
          6488 => x"80",
          6489 => x"89",
          6490 => x"2a",
          6491 => x"51",
          6492 => x"2e",
          6493 => x"51",
          6494 => x"3f",
          6495 => x"51",
          6496 => x"3f",
          6497 => x"d7",
          6498 => x"87",
          6499 => x"06",
          6500 => x"80",
          6501 => x"81",
          6502 => x"d5",
          6503 => x"a8",
          6504 => x"cd",
          6505 => x"fe",
          6506 => x"72",
          6507 => x"81",
          6508 => x"71",
          6509 => x"38",
          6510 => x"d7",
          6511 => x"ef",
          6512 => x"d9",
          6513 => x"51",
          6514 => x"3f",
          6515 => x"3f",
          6516 => x"04",
          6517 => x"77",
          6518 => x"a3",
          6519 => x"55",
          6520 => x"52",
          6521 => x"ce",
          6522 => x"f5",
          6523 => x"73",
          6524 => x"53",
          6525 => x"52",
          6526 => x"51",
          6527 => x"3f",
          6528 => x"08",
          6529 => x"f8",
          6530 => x"80",
          6531 => x"31",
          6532 => x"73",
          6533 => x"34",
          6534 => x"33",
          6535 => x"2e",
          6536 => x"ac",
          6537 => x"e0",
          6538 => x"75",
          6539 => x"3f",
          6540 => x"08",
          6541 => x"38",
          6542 => x"08",
          6543 => x"a4",
          6544 => x"82",
          6545 => x"c4",
          6546 => x"0b",
          6547 => x"34",
          6548 => x"33",
          6549 => x"2e",
          6550 => x"89",
          6551 => x"75",
          6552 => x"e4",
          6553 => x"81",
          6554 => x"87",
          6555 => x"ce",
          6556 => x"70",
          6557 => x"dc",
          6558 => x"81",
          6559 => x"ff",
          6560 => x"81",
          6561 => x"81",
          6562 => x"78",
          6563 => x"81",
          6564 => x"81",
          6565 => x"96",
          6566 => x"59",
          6567 => x"3f",
          6568 => x"52",
          6569 => x"51",
          6570 => x"3f",
          6571 => x"08",
          6572 => x"38",
          6573 => x"51",
          6574 => x"81",
          6575 => x"81",
          6576 => x"fe",
          6577 => x"96",
          6578 => x"5a",
          6579 => x"79",
          6580 => x"3f",
          6581 => x"84",
          6582 => x"c2",
          6583 => x"c8",
          6584 => x"70",
          6585 => x"59",
          6586 => x"2e",
          6587 => x"78",
          6588 => x"b2",
          6589 => x"2e",
          6590 => x"78",
          6591 => x"38",
          6592 => x"ff",
          6593 => x"bc",
          6594 => x"38",
          6595 => x"78",
          6596 => x"83",
          6597 => x"80",
          6598 => x"dd",
          6599 => x"2e",
          6600 => x"8a",
          6601 => x"80",
          6602 => x"ea",
          6603 => x"f9",
          6604 => x"78",
          6605 => x"88",
          6606 => x"80",
          6607 => x"b1",
          6608 => x"39",
          6609 => x"2e",
          6610 => x"78",
          6611 => x"8b",
          6612 => x"82",
          6613 => x"38",
          6614 => x"78",
          6615 => x"8a",
          6616 => x"93",
          6617 => x"ff",
          6618 => x"ff",
          6619 => x"fe",
          6620 => x"81",
          6621 => x"80",
          6622 => x"38",
          6623 => x"fc",
          6624 => x"84",
          6625 => x"ee",
          6626 => x"f8",
          6627 => x"2e",
          6628 => x"b4",
          6629 => x"11",
          6630 => x"05",
          6631 => x"9d",
          6632 => x"c8",
          6633 => x"81",
          6634 => x"42",
          6635 => x"51",
          6636 => x"3f",
          6637 => x"5a",
          6638 => x"81",
          6639 => x"59",
          6640 => x"84",
          6641 => x"7a",
          6642 => x"38",
          6643 => x"b4",
          6644 => x"11",
          6645 => x"05",
          6646 => x"e1",
          6647 => x"c8",
          6648 => x"fd",
          6649 => x"3d",
          6650 => x"53",
          6651 => x"51",
          6652 => x"3f",
          6653 => x"08",
          6654 => x"c3",
          6655 => x"fe",
          6656 => x"ff",
          6657 => x"fe",
          6658 => x"81",
          6659 => x"80",
          6660 => x"38",
          6661 => x"51",
          6662 => x"3f",
          6663 => x"63",
          6664 => x"38",
          6665 => x"70",
          6666 => x"33",
          6667 => x"81",
          6668 => x"39",
          6669 => x"80",
          6670 => x"84",
          6671 => x"ec",
          6672 => x"f8",
          6673 => x"2e",
          6674 => x"b4",
          6675 => x"11",
          6676 => x"05",
          6677 => x"e5",
          6678 => x"c8",
          6679 => x"fc",
          6680 => x"3d",
          6681 => x"53",
          6682 => x"51",
          6683 => x"3f",
          6684 => x"08",
          6685 => x"c7",
          6686 => x"e8",
          6687 => x"e4",
          6688 => x"79",
          6689 => x"38",
          6690 => x"7b",
          6691 => x"5b",
          6692 => x"92",
          6693 => x"7a",
          6694 => x"53",
          6695 => x"f0",
          6696 => x"ea",
          6697 => x"1a",
          6698 => x"43",
          6699 => x"81",
          6700 => x"82",
          6701 => x"3d",
          6702 => x"53",
          6703 => x"51",
          6704 => x"3f",
          6705 => x"08",
          6706 => x"81",
          6707 => x"59",
          6708 => x"89",
          6709 => x"c4",
          6710 => x"cd",
          6711 => x"8d",
          6712 => x"80",
          6713 => x"81",
          6714 => x"44",
          6715 => x"f4",
          6716 => x"78",
          6717 => x"38",
          6718 => x"08",
          6719 => x"81",
          6720 => x"59",
          6721 => x"88",
          6722 => x"dc",
          6723 => x"39",
          6724 => x"33",
          6725 => x"2e",
          6726 => x"f3",
          6727 => x"89",
          6728 => x"f4",
          6729 => x"05",
          6730 => x"fe",
          6731 => x"ff",
          6732 => x"fe",
          6733 => x"81",
          6734 => x"80",
          6735 => x"f4",
          6736 => x"78",
          6737 => x"38",
          6738 => x"08",
          6739 => x"39",
          6740 => x"33",
          6741 => x"2e",
          6742 => x"f3",
          6743 => x"bb",
          6744 => x"8e",
          6745 => x"80",
          6746 => x"81",
          6747 => x"43",
          6748 => x"f4",
          6749 => x"78",
          6750 => x"38",
          6751 => x"08",
          6752 => x"81",
          6753 => x"59",
          6754 => x"88",
          6755 => x"e8",
          6756 => x"39",
          6757 => x"08",
          6758 => x"b4",
          6759 => x"11",
          6760 => x"05",
          6761 => x"95",
          6762 => x"c8",
          6763 => x"a7",
          6764 => x"5c",
          6765 => x"2e",
          6766 => x"5c",
          6767 => x"70",
          6768 => x"07",
          6769 => x"7f",
          6770 => x"5a",
          6771 => x"2e",
          6772 => x"a0",
          6773 => x"88",
          6774 => x"94",
          6775 => x"84",
          6776 => x"63",
          6777 => x"62",
          6778 => x"f2",
          6779 => x"f1",
          6780 => x"e1",
          6781 => x"c7",
          6782 => x"ff",
          6783 => x"ff",
          6784 => x"fe",
          6785 => x"81",
          6786 => x"80",
          6787 => x"38",
          6788 => x"fc",
          6789 => x"84",
          6790 => x"e9",
          6791 => x"f8",
          6792 => x"2e",
          6793 => x"59",
          6794 => x"05",
          6795 => x"63",
          6796 => x"b4",
          6797 => x"11",
          6798 => x"05",
          6799 => x"fd",
          6800 => x"c8",
          6801 => x"f8",
          6802 => x"70",
          6803 => x"81",
          6804 => x"fe",
          6805 => x"80",
          6806 => x"51",
          6807 => x"3f",
          6808 => x"33",
          6809 => x"2e",
          6810 => x"9f",
          6811 => x"38",
          6812 => x"fc",
          6813 => x"84",
          6814 => x"e8",
          6815 => x"f8",
          6816 => x"2e",
          6817 => x"59",
          6818 => x"05",
          6819 => x"63",
          6820 => x"ff",
          6821 => x"f1",
          6822 => x"e0",
          6823 => x"aa",
          6824 => x"fe",
          6825 => x"ff",
          6826 => x"fe",
          6827 => x"81",
          6828 => x"80",
          6829 => x"38",
          6830 => x"f0",
          6831 => x"84",
          6832 => x"e9",
          6833 => x"f8",
          6834 => x"2e",
          6835 => x"59",
          6836 => x"22",
          6837 => x"05",
          6838 => x"41",
          6839 => x"f0",
          6840 => x"84",
          6841 => x"e9",
          6842 => x"f8",
          6843 => x"38",
          6844 => x"60",
          6845 => x"52",
          6846 => x"51",
          6847 => x"3f",
          6848 => x"79",
          6849 => x"9a",
          6850 => x"79",
          6851 => x"ae",
          6852 => x"38",
          6853 => x"87",
          6854 => x"05",
          6855 => x"b4",
          6856 => x"11",
          6857 => x"05",
          6858 => x"83",
          6859 => x"c8",
          6860 => x"92",
          6861 => x"02",
          6862 => x"79",
          6863 => x"5b",
          6864 => x"ff",
          6865 => x"f1",
          6866 => x"df",
          6867 => x"a3",
          6868 => x"fe",
          6869 => x"ff",
          6870 => x"fe",
          6871 => x"81",
          6872 => x"80",
          6873 => x"38",
          6874 => x"f0",
          6875 => x"84",
          6876 => x"e8",
          6877 => x"f8",
          6878 => x"2e",
          6879 => x"60",
          6880 => x"60",
          6881 => x"b4",
          6882 => x"11",
          6883 => x"05",
          6884 => x"9b",
          6885 => x"c8",
          6886 => x"f6",
          6887 => x"70",
          6888 => x"81",
          6889 => x"fe",
          6890 => x"80",
          6891 => x"51",
          6892 => x"3f",
          6893 => x"33",
          6894 => x"2e",
          6895 => x"9f",
          6896 => x"38",
          6897 => x"f0",
          6898 => x"84",
          6899 => x"e7",
          6900 => x"f8",
          6901 => x"2e",
          6902 => x"60",
          6903 => x"60",
          6904 => x"ff",
          6905 => x"f1",
          6906 => x"dd",
          6907 => x"ae",
          6908 => x"ff",
          6909 => x"ff",
          6910 => x"fe",
          6911 => x"81",
          6912 => x"80",
          6913 => x"38",
          6914 => x"f1",
          6915 => x"e3",
          6916 => x"59",
          6917 => x"3d",
          6918 => x"53",
          6919 => x"51",
          6920 => x"3f",
          6921 => x"08",
          6922 => x"93",
          6923 => x"81",
          6924 => x"fe",
          6925 => x"63",
          6926 => x"81",
          6927 => x"80",
          6928 => x"38",
          6929 => x"08",
          6930 => x"94",
          6931 => x"f8",
          6932 => x"39",
          6933 => x"51",
          6934 => x"3f",
          6935 => x"3f",
          6936 => x"81",
          6937 => x"fe",
          6938 => x"80",
          6939 => x"39",
          6940 => x"3f",
          6941 => x"79",
          6942 => x"59",
          6943 => x"f4",
          6944 => x"7d",
          6945 => x"80",
          6946 => x"38",
          6947 => x"84",
          6948 => x"c6",
          6949 => x"f8",
          6950 => x"81",
          6951 => x"2e",
          6952 => x"82",
          6953 => x"7a",
          6954 => x"38",
          6955 => x"7a",
          6956 => x"38",
          6957 => x"81",
          6958 => x"7b",
          6959 => x"e4",
          6960 => x"81",
          6961 => x"b4",
          6962 => x"05",
          6963 => x"8e",
          6964 => x"81",
          6965 => x"b4",
          6966 => x"05",
          6967 => x"fe",
          6968 => x"7b",
          6969 => x"e4",
          6970 => x"81",
          6971 => x"b4",
          6972 => x"05",
          6973 => x"e6",
          6974 => x"7b",
          6975 => x"81",
          6976 => x"b4",
          6977 => x"05",
          6978 => x"d2",
          6979 => x"c4",
          6980 => x"90",
          6981 => x"64",
          6982 => x"83",
          6983 => x"83",
          6984 => x"b4",
          6985 => x"05",
          6986 => x"3f",
          6987 => x"08",
          6988 => x"08",
          6989 => x"70",
          6990 => x"25",
          6991 => x"5f",
          6992 => x"83",
          6993 => x"81",
          6994 => x"06",
          6995 => x"2e",
          6996 => x"1b",
          6997 => x"06",
          6998 => x"fe",
          6999 => x"81",
          7000 => x"32",
          7001 => x"8a",
          7002 => x"2e",
          7003 => x"f2",
          7004 => x"f3",
          7005 => x"e0",
          7006 => x"c3",
          7007 => x"0d",
          7008 => x"f9",
          7009 => x"c0",
          7010 => x"08",
          7011 => x"84",
          7012 => x"51",
          7013 => x"3f",
          7014 => x"08",
          7015 => x"08",
          7016 => x"84",
          7017 => x"51",
          7018 => x"3f",
          7019 => x"c8",
          7020 => x"0c",
          7021 => x"9c",
          7022 => x"55",
          7023 => x"52",
          7024 => x"b7",
          7025 => x"f8",
          7026 => x"2b",
          7027 => x"53",
          7028 => x"52",
          7029 => x"b7",
          7030 => x"81",
          7031 => x"07",
          7032 => x"80",
          7033 => x"c0",
          7034 => x"8c",
          7035 => x"87",
          7036 => x"0c",
          7037 => x"81",
          7038 => x"a6",
          7039 => x"f8",
          7040 => x"cb",
          7041 => x"d4",
          7042 => x"f3",
          7043 => x"d9",
          7044 => x"f3",
          7045 => x"d9",
          7046 => x"c9",
          7047 => x"d4",
          7048 => x"51",
          7049 => x"f0",
          7050 => x"04",
          7051 => x"ff",
          7052 => x"ff",
          7053 => x"ff",
          7054 => x"00",
          7055 => x"32",
          7056 => x"38",
          7057 => x"3e",
          7058 => x"44",
          7059 => x"4a",
          7060 => x"b5",
          7061 => x"91",
          7062 => x"34",
          7063 => x"74",
          7064 => x"97",
          7065 => x"24",
          7066 => x"8a",
          7067 => x"8a",
          7068 => x"61",
          7069 => x"d7",
          7070 => x"62",
          7071 => x"8b",
          7072 => x"a9",
          7073 => x"2d",
          7074 => x"34",
          7075 => x"3b",
          7076 => x"42",
          7077 => x"49",
          7078 => x"50",
          7079 => x"57",
          7080 => x"5e",
          7081 => x"65",
          7082 => x"6c",
          7083 => x"73",
          7084 => x"79",
          7085 => x"7f",
          7086 => x"85",
          7087 => x"8b",
          7088 => x"91",
          7089 => x"97",
          7090 => x"9d",
          7091 => x"a3",
          7092 => x"25",
          7093 => x"64",
          7094 => x"3a",
          7095 => x"25",
          7096 => x"64",
          7097 => x"00",
          7098 => x"20",
          7099 => x"66",
          7100 => x"72",
          7101 => x"6f",
          7102 => x"00",
          7103 => x"72",
          7104 => x"53",
          7105 => x"63",
          7106 => x"69",
          7107 => x"00",
          7108 => x"65",
          7109 => x"65",
          7110 => x"6d",
          7111 => x"6d",
          7112 => x"65",
          7113 => x"00",
          7114 => x"20",
          7115 => x"53",
          7116 => x"4d",
          7117 => x"25",
          7118 => x"3a",
          7119 => x"58",
          7120 => x"00",
          7121 => x"20",
          7122 => x"41",
          7123 => x"20",
          7124 => x"25",
          7125 => x"3a",
          7126 => x"58",
          7127 => x"00",
          7128 => x"20",
          7129 => x"4e",
          7130 => x"41",
          7131 => x"25",
          7132 => x"3a",
          7133 => x"58",
          7134 => x"00",
          7135 => x"20",
          7136 => x"4d",
          7137 => x"20",
          7138 => x"25",
          7139 => x"3a",
          7140 => x"58",
          7141 => x"00",
          7142 => x"20",
          7143 => x"20",
          7144 => x"20",
          7145 => x"25",
          7146 => x"3a",
          7147 => x"58",
          7148 => x"00",
          7149 => x"20",
          7150 => x"43",
          7151 => x"20",
          7152 => x"44",
          7153 => x"63",
          7154 => x"3d",
          7155 => x"64",
          7156 => x"00",
          7157 => x"20",
          7158 => x"45",
          7159 => x"20",
          7160 => x"54",
          7161 => x"72",
          7162 => x"3d",
          7163 => x"64",
          7164 => x"00",
          7165 => x"20",
          7166 => x"52",
          7167 => x"52",
          7168 => x"43",
          7169 => x"6e",
          7170 => x"3d",
          7171 => x"64",
          7172 => x"00",
          7173 => x"20",
          7174 => x"48",
          7175 => x"45",
          7176 => x"53",
          7177 => x"00",
          7178 => x"20",
          7179 => x"49",
          7180 => x"00",
          7181 => x"20",
          7182 => x"54",
          7183 => x"00",
          7184 => x"20",
          7185 => x"0a",
          7186 => x"00",
          7187 => x"20",
          7188 => x"0a",
          7189 => x"00",
          7190 => x"72",
          7191 => x"65",
          7192 => x"00",
          7193 => x"20",
          7194 => x"20",
          7195 => x"65",
          7196 => x"65",
          7197 => x"72",
          7198 => x"64",
          7199 => x"73",
          7200 => x"25",
          7201 => x"0a",
          7202 => x"00",
          7203 => x"20",
          7204 => x"20",
          7205 => x"6f",
          7206 => x"53",
          7207 => x"74",
          7208 => x"64",
          7209 => x"73",
          7210 => x"25",
          7211 => x"0a",
          7212 => x"00",
          7213 => x"20",
          7214 => x"63",
          7215 => x"74",
          7216 => x"20",
          7217 => x"72",
          7218 => x"20",
          7219 => x"20",
          7220 => x"25",
          7221 => x"0a",
          7222 => x"00",
          7223 => x"63",
          7224 => x"00",
          7225 => x"20",
          7226 => x"20",
          7227 => x"20",
          7228 => x"20",
          7229 => x"20",
          7230 => x"20",
          7231 => x"20",
          7232 => x"25",
          7233 => x"0a",
          7234 => x"00",
          7235 => x"20",
          7236 => x"74",
          7237 => x"43",
          7238 => x"6b",
          7239 => x"65",
          7240 => x"20",
          7241 => x"20",
          7242 => x"25",
          7243 => x"30",
          7244 => x"48",
          7245 => x"00",
          7246 => x"20",
          7247 => x"41",
          7248 => x"6c",
          7249 => x"20",
          7250 => x"71",
          7251 => x"20",
          7252 => x"20",
          7253 => x"25",
          7254 => x"30",
          7255 => x"48",
          7256 => x"00",
          7257 => x"20",
          7258 => x"68",
          7259 => x"65",
          7260 => x"52",
          7261 => x"43",
          7262 => x"6b",
          7263 => x"65",
          7264 => x"25",
          7265 => x"30",
          7266 => x"48",
          7267 => x"00",
          7268 => x"6c",
          7269 => x"00",
          7270 => x"69",
          7271 => x"00",
          7272 => x"78",
          7273 => x"00",
          7274 => x"00",
          7275 => x"6d",
          7276 => x"00",
          7277 => x"6e",
          7278 => x"00",
          7279 => x"74",
          7280 => x"2e",
          7281 => x"00",
          7282 => x"74",
          7283 => x"00",
          7284 => x"74",
          7285 => x"00",
          7286 => x"00",
          7287 => x"64",
          7288 => x"73",
          7289 => x"00",
          7290 => x"6c",
          7291 => x"74",
          7292 => x"65",
          7293 => x"20",
          7294 => x"20",
          7295 => x"74",
          7296 => x"20",
          7297 => x"65",
          7298 => x"20",
          7299 => x"2e",
          7300 => x"00",
          7301 => x"6e",
          7302 => x"6f",
          7303 => x"2f",
          7304 => x"61",
          7305 => x"68",
          7306 => x"6f",
          7307 => x"66",
          7308 => x"2c",
          7309 => x"73",
          7310 => x"69",
          7311 => x"0a",
          7312 => x"00",
          7313 => x"f0",
          7314 => x"00",
          7315 => x"01",
          7316 => x"ec",
          7317 => x"00",
          7318 => x"02",
          7319 => x"e8",
          7320 => x"00",
          7321 => x"03",
          7322 => x"e4",
          7323 => x"00",
          7324 => x"04",
          7325 => x"e0",
          7326 => x"00",
          7327 => x"05",
          7328 => x"dc",
          7329 => x"00",
          7330 => x"06",
          7331 => x"d8",
          7332 => x"00",
          7333 => x"07",
          7334 => x"d4",
          7335 => x"00",
          7336 => x"08",
          7337 => x"d0",
          7338 => x"00",
          7339 => x"09",
          7340 => x"cc",
          7341 => x"00",
          7342 => x"0a",
          7343 => x"c8",
          7344 => x"00",
          7345 => x"0b",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"7e",
          7351 => x"7e",
          7352 => x"7e",
          7353 => x"7e",
          7354 => x"7e",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"2c",
          7359 => x"3d",
          7360 => x"5d",
          7361 => x"00",
          7362 => x"00",
          7363 => x"33",
          7364 => x"00",
          7365 => x"4d",
          7366 => x"53",
          7367 => x"00",
          7368 => x"4e",
          7369 => x"20",
          7370 => x"46",
          7371 => x"32",
          7372 => x"00",
          7373 => x"4e",
          7374 => x"20",
          7375 => x"46",
          7376 => x"20",
          7377 => x"00",
          7378 => x"f4",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"41",
          7383 => x"80",
          7384 => x"49",
          7385 => x"8f",
          7386 => x"4f",
          7387 => x"55",
          7388 => x"9b",
          7389 => x"9f",
          7390 => x"55",
          7391 => x"a7",
          7392 => x"ab",
          7393 => x"af",
          7394 => x"b3",
          7395 => x"b7",
          7396 => x"bb",
          7397 => x"bf",
          7398 => x"c3",
          7399 => x"c7",
          7400 => x"cb",
          7401 => x"cf",
          7402 => x"d3",
          7403 => x"d7",
          7404 => x"db",
          7405 => x"df",
          7406 => x"e3",
          7407 => x"e7",
          7408 => x"eb",
          7409 => x"ef",
          7410 => x"f3",
          7411 => x"f7",
          7412 => x"fb",
          7413 => x"ff",
          7414 => x"3b",
          7415 => x"2f",
          7416 => x"3a",
          7417 => x"7c",
          7418 => x"00",
          7419 => x"04",
          7420 => x"40",
          7421 => x"00",
          7422 => x"00",
          7423 => x"02",
          7424 => x"08",
          7425 => x"20",
          7426 => x"00",
          7427 => x"69",
          7428 => x"00",
          7429 => x"63",
          7430 => x"00",
          7431 => x"69",
          7432 => x"00",
          7433 => x"61",
          7434 => x"00",
          7435 => x"65",
          7436 => x"00",
          7437 => x"65",
          7438 => x"00",
          7439 => x"70",
          7440 => x"00",
          7441 => x"66",
          7442 => x"00",
          7443 => x"6d",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"6c",
          7453 => x"00",
          7454 => x"00",
          7455 => x"74",
          7456 => x"00",
          7457 => x"65",
          7458 => x"00",
          7459 => x"6f",
          7460 => x"00",
          7461 => x"74",
          7462 => x"00",
          7463 => x"73",
          7464 => x"00",
          7465 => x"73",
          7466 => x"00",
          7467 => x"6f",
          7468 => x"00",
          7469 => x"6b",
          7470 => x"72",
          7471 => x"00",
          7472 => x"65",
          7473 => x"6c",
          7474 => x"72",
          7475 => x"0a",
          7476 => x"00",
          7477 => x"6b",
          7478 => x"74",
          7479 => x"61",
          7480 => x"0a",
          7481 => x"00",
          7482 => x"66",
          7483 => x"20",
          7484 => x"6e",
          7485 => x"00",
          7486 => x"70",
          7487 => x"20",
          7488 => x"6e",
          7489 => x"00",
          7490 => x"61",
          7491 => x"20",
          7492 => x"65",
          7493 => x"65",
          7494 => x"00",
          7495 => x"65",
          7496 => x"64",
          7497 => x"65",
          7498 => x"00",
          7499 => x"65",
          7500 => x"72",
          7501 => x"79",
          7502 => x"69",
          7503 => x"2e",
          7504 => x"00",
          7505 => x"65",
          7506 => x"6e",
          7507 => x"20",
          7508 => x"61",
          7509 => x"2e",
          7510 => x"00",
          7511 => x"69",
          7512 => x"72",
          7513 => x"20",
          7514 => x"74",
          7515 => x"65",
          7516 => x"00",
          7517 => x"76",
          7518 => x"75",
          7519 => x"72",
          7520 => x"20",
          7521 => x"61",
          7522 => x"2e",
          7523 => x"00",
          7524 => x"6b",
          7525 => x"74",
          7526 => x"61",
          7527 => x"64",
          7528 => x"00",
          7529 => x"63",
          7530 => x"61",
          7531 => x"6c",
          7532 => x"69",
          7533 => x"79",
          7534 => x"6d",
          7535 => x"75",
          7536 => x"6f",
          7537 => x"69",
          7538 => x"0a",
          7539 => x"00",
          7540 => x"6d",
          7541 => x"61",
          7542 => x"74",
          7543 => x"0a",
          7544 => x"00",
          7545 => x"65",
          7546 => x"2c",
          7547 => x"65",
          7548 => x"69",
          7549 => x"63",
          7550 => x"65",
          7551 => x"64",
          7552 => x"00",
          7553 => x"65",
          7554 => x"20",
          7555 => x"6b",
          7556 => x"0a",
          7557 => x"00",
          7558 => x"75",
          7559 => x"63",
          7560 => x"74",
          7561 => x"6d",
          7562 => x"2e",
          7563 => x"00",
          7564 => x"20",
          7565 => x"79",
          7566 => x"65",
          7567 => x"69",
          7568 => x"2e",
          7569 => x"00",
          7570 => x"61",
          7571 => x"65",
          7572 => x"69",
          7573 => x"72",
          7574 => x"74",
          7575 => x"00",
          7576 => x"63",
          7577 => x"2e",
          7578 => x"00",
          7579 => x"6e",
          7580 => x"20",
          7581 => x"6f",
          7582 => x"00",
          7583 => x"75",
          7584 => x"74",
          7585 => x"25",
          7586 => x"74",
          7587 => x"75",
          7588 => x"74",
          7589 => x"73",
          7590 => x"0a",
          7591 => x"00",
          7592 => x"64",
          7593 => x"00",
          7594 => x"58",
          7595 => x"00",
          7596 => x"00",
          7597 => x"58",
          7598 => x"00",
          7599 => x"20",
          7600 => x"20",
          7601 => x"00",
          7602 => x"58",
          7603 => x"00",
          7604 => x"00",
          7605 => x"00",
          7606 => x"00",
          7607 => x"00",
          7608 => x"20",
          7609 => x"28",
          7610 => x"00",
          7611 => x"30",
          7612 => x"30",
          7613 => x"00",
          7614 => x"30",
          7615 => x"00",
          7616 => x"55",
          7617 => x"65",
          7618 => x"30",
          7619 => x"20",
          7620 => x"25",
          7621 => x"2a",
          7622 => x"00",
          7623 => x"20",
          7624 => x"65",
          7625 => x"70",
          7626 => x"61",
          7627 => x"65",
          7628 => x"00",
          7629 => x"65",
          7630 => x"6e",
          7631 => x"72",
          7632 => x"0a",
          7633 => x"00",
          7634 => x"20",
          7635 => x"65",
          7636 => x"70",
          7637 => x"00",
          7638 => x"54",
          7639 => x"44",
          7640 => x"74",
          7641 => x"75",
          7642 => x"00",
          7643 => x"54",
          7644 => x"52",
          7645 => x"74",
          7646 => x"75",
          7647 => x"00",
          7648 => x"54",
          7649 => x"58",
          7650 => x"74",
          7651 => x"75",
          7652 => x"00",
          7653 => x"54",
          7654 => x"58",
          7655 => x"74",
          7656 => x"75",
          7657 => x"00",
          7658 => x"54",
          7659 => x"58",
          7660 => x"74",
          7661 => x"75",
          7662 => x"00",
          7663 => x"54",
          7664 => x"58",
          7665 => x"74",
          7666 => x"75",
          7667 => x"00",
          7668 => x"74",
          7669 => x"20",
          7670 => x"74",
          7671 => x"72",
          7672 => x"0a",
          7673 => x"00",
          7674 => x"62",
          7675 => x"67",
          7676 => x"6d",
          7677 => x"2e",
          7678 => x"00",
          7679 => x"6f",
          7680 => x"63",
          7681 => x"74",
          7682 => x"00",
          7683 => x"00",
          7684 => x"6c",
          7685 => x"74",
          7686 => x"6e",
          7687 => x"61",
          7688 => x"65",
          7689 => x"20",
          7690 => x"64",
          7691 => x"20",
          7692 => x"61",
          7693 => x"69",
          7694 => x"20",
          7695 => x"75",
          7696 => x"79",
          7697 => x"00",
          7698 => x"00",
          7699 => x"61",
          7700 => x"67",
          7701 => x"2e",
          7702 => x"00",
          7703 => x"79",
          7704 => x"2e",
          7705 => x"00",
          7706 => x"70",
          7707 => x"6e",
          7708 => x"2e",
          7709 => x"00",
          7710 => x"6c",
          7711 => x"30",
          7712 => x"2d",
          7713 => x"38",
          7714 => x"25",
          7715 => x"29",
          7716 => x"00",
          7717 => x"70",
          7718 => x"6d",
          7719 => x"0a",
          7720 => x"00",
          7721 => x"6d",
          7722 => x"74",
          7723 => x"00",
          7724 => x"58",
          7725 => x"32",
          7726 => x"00",
          7727 => x"0a",
          7728 => x"00",
          7729 => x"58",
          7730 => x"34",
          7731 => x"00",
          7732 => x"58",
          7733 => x"38",
          7734 => x"00",
          7735 => x"63",
          7736 => x"6e",
          7737 => x"6f",
          7738 => x"40",
          7739 => x"38",
          7740 => x"2e",
          7741 => x"00",
          7742 => x"6c",
          7743 => x"20",
          7744 => x"65",
          7745 => x"25",
          7746 => x"20",
          7747 => x"0a",
          7748 => x"00",
          7749 => x"6c",
          7750 => x"74",
          7751 => x"65",
          7752 => x"6f",
          7753 => x"28",
          7754 => x"2e",
          7755 => x"00",
          7756 => x"74",
          7757 => x"69",
          7758 => x"61",
          7759 => x"69",
          7760 => x"69",
          7761 => x"2e",
          7762 => x"00",
          7763 => x"64",
          7764 => x"62",
          7765 => x"69",
          7766 => x"2e",
          7767 => x"00",
          7768 => x"00",
          7769 => x"00",
          7770 => x"5c",
          7771 => x"25",
          7772 => x"73",
          7773 => x"00",
          7774 => x"5c",
          7775 => x"25",
          7776 => x"00",
          7777 => x"5c",
          7778 => x"00",
          7779 => x"20",
          7780 => x"6d",
          7781 => x"2e",
          7782 => x"00",
          7783 => x"6e",
          7784 => x"2e",
          7785 => x"00",
          7786 => x"62",
          7787 => x"67",
          7788 => x"74",
          7789 => x"75",
          7790 => x"2e",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"ff",
          7795 => x"00",
          7796 => x"ff",
          7797 => x"00",
          7798 => x"ff",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"ff",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"00",
          7810 => x"00",
          7811 => x"01",
          7812 => x"01",
          7813 => x"01",
          7814 => x"00",
          7815 => x"00",
          7816 => x"02",
          7817 => x"00",
          7818 => x"20",
          7819 => x"20",
          7820 => x"20",
          7821 => x"20",
          7822 => x"bc",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"c8",
          7847 => x"00",
          7848 => x"d0",
          7849 => x"00",
          7850 => x"d8",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"0c",
          7855 => x"00",
          7856 => x"00",
          7857 => x"00",
          7858 => x"14",
          7859 => x"00",
          7860 => x"00",
          7861 => x"00",
          7862 => x"1c",
          7863 => x"00",
          7864 => x"00",
          7865 => x"00",
          7866 => x"24",
          7867 => x"00",
          7868 => x"00",
          7869 => x"00",
          7870 => x"2c",
          7871 => x"00",
          7872 => x"00",
          7873 => x"00",
          7874 => x"34",
          7875 => x"00",
          7876 => x"00",
          7877 => x"00",
          7878 => x"3c",
          7879 => x"00",
          7880 => x"00",
          7881 => x"00",
          7882 => x"44",
          7883 => x"00",
          7884 => x"00",
          7885 => x"00",
          7886 => x"4c",
          7887 => x"00",
          7888 => x"00",
          7889 => x"00",
          7890 => x"54",
          7891 => x"00",
          7892 => x"00",
          7893 => x"00",
          7894 => x"58",
          7895 => x"00",
          7896 => x"00",
          7897 => x"00",
          7898 => x"5c",
          7899 => x"00",
          7900 => x"00",
          7901 => x"00",
          7902 => x"60",
          7903 => x"00",
          7904 => x"00",
          7905 => x"00",
          7906 => x"64",
          7907 => x"00",
          7908 => x"00",
          7909 => x"00",
          7910 => x"68",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"6c",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"70",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"78",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"7c",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"84",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"8c",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"94",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"9c",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"a4",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"ac",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a3",
           270 => x"0b",
           271 => x"0b",
           272 => x"c1",
           273 => x"0b",
           274 => x"0b",
           275 => x"df",
           276 => x"0b",
           277 => x"0b",
           278 => x"fd",
           279 => x"0b",
           280 => x"0b",
           281 => x"9b",
           282 => x"0b",
           283 => x"0b",
           284 => x"b9",
           285 => x"0b",
           286 => x"0b",
           287 => x"d7",
           288 => x"0b",
           289 => x"0b",
           290 => x"f5",
           291 => x"0b",
           292 => x"0b",
           293 => x"93",
           294 => x"0b",
           295 => x"0b",
           296 => x"b3",
           297 => x"0b",
           298 => x"0b",
           299 => x"d3",
           300 => x"0b",
           301 => x"0b",
           302 => x"f3",
           303 => x"0b",
           304 => x"0b",
           305 => x"93",
           306 => x"0b",
           307 => x"0b",
           308 => x"b3",
           309 => x"0b",
           310 => x"0b",
           311 => x"d3",
           312 => x"0b",
           313 => x"0b",
           314 => x"f3",
           315 => x"0b",
           316 => x"0b",
           317 => x"93",
           318 => x"0b",
           319 => x"0b",
           320 => x"b3",
           321 => x"0b",
           322 => x"0b",
           323 => x"d3",
           324 => x"0b",
           325 => x"0b",
           326 => x"f3",
           327 => x"0b",
           328 => x"0b",
           329 => x"93",
           330 => x"0b",
           331 => x"0b",
           332 => x"b3",
           333 => x"0b",
           334 => x"0b",
           335 => x"d3",
           336 => x"0b",
           337 => x"0b",
           338 => x"f3",
           339 => x"0b",
           340 => x"0b",
           341 => x"91",
           342 => x"0b",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"f8",
           386 => x"ff",
           387 => x"d4",
           388 => x"90",
           389 => x"d4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"81",
           395 => x"83",
           396 => x"81",
           397 => x"b5",
           398 => x"f8",
           399 => x"80",
           400 => x"f8",
           401 => x"a2",
           402 => x"d4",
           403 => x"90",
           404 => x"d4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"81",
           410 => x"83",
           411 => x"81",
           412 => x"bd",
           413 => x"f8",
           414 => x"80",
           415 => x"f8",
           416 => x"af",
           417 => x"d4",
           418 => x"90",
           419 => x"d4",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"81",
           425 => x"83",
           426 => x"81",
           427 => x"bb",
           428 => x"f8",
           429 => x"80",
           430 => x"f8",
           431 => x"82",
           432 => x"d4",
           433 => x"90",
           434 => x"d4",
           435 => x"2d",
           436 => x"08",
           437 => x"04",
           438 => x"0c",
           439 => x"81",
           440 => x"83",
           441 => x"81",
           442 => x"9e",
           443 => x"f8",
           444 => x"80",
           445 => x"f8",
           446 => x"ae",
           447 => x"d4",
           448 => x"90",
           449 => x"d4",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"04",
           565 => x"0c",
           566 => x"2d",
           567 => x"08",
           568 => x"04",
           569 => x"0c",
           570 => x"2d",
           571 => x"08",
           572 => x"04",
           573 => x"0c",
           574 => x"81",
           575 => x"83",
           576 => x"81",
           577 => x"a0",
           578 => x"f8",
           579 => x"80",
           580 => x"f8",
           581 => x"f1",
           582 => x"d4",
           583 => x"90",
           584 => x"d4",
           585 => x"97",
           586 => x"d4",
           587 => x"90",
           588 => x"00",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"00",
           598 => x"ff",
           599 => x"06",
           600 => x"83",
           601 => x"10",
           602 => x"fc",
           603 => x"51",
           604 => x"80",
           605 => x"ff",
           606 => x"06",
           607 => x"52",
           608 => x"0a",
           609 => x"38",
           610 => x"51",
           611 => x"c8",
           612 => x"88",
           613 => x"80",
           614 => x"05",
           615 => x"0b",
           616 => x"04",
           617 => x"81",
           618 => x"00",
           619 => x"08",
           620 => x"d4",
           621 => x"0d",
           622 => x"f8",
           623 => x"05",
           624 => x"f8",
           625 => x"05",
           626 => x"d4",
           627 => x"c8",
           628 => x"f8",
           629 => x"85",
           630 => x"f8",
           631 => x"81",
           632 => x"02",
           633 => x"0c",
           634 => x"81",
           635 => x"d4",
           636 => x"08",
           637 => x"d4",
           638 => x"08",
           639 => x"3f",
           640 => x"08",
           641 => x"c8",
           642 => x"3d",
           643 => x"d4",
           644 => x"f8",
           645 => x"81",
           646 => x"f9",
           647 => x"0b",
           648 => x"08",
           649 => x"81",
           650 => x"88",
           651 => x"25",
           652 => x"f8",
           653 => x"05",
           654 => x"f8",
           655 => x"05",
           656 => x"81",
           657 => x"f4",
           658 => x"f8",
           659 => x"05",
           660 => x"81",
           661 => x"d4",
           662 => x"0c",
           663 => x"08",
           664 => x"81",
           665 => x"fc",
           666 => x"f8",
           667 => x"05",
           668 => x"b9",
           669 => x"d4",
           670 => x"08",
           671 => x"d4",
           672 => x"0c",
           673 => x"f8",
           674 => x"05",
           675 => x"d4",
           676 => x"08",
           677 => x"0b",
           678 => x"08",
           679 => x"81",
           680 => x"f0",
           681 => x"f8",
           682 => x"05",
           683 => x"81",
           684 => x"8c",
           685 => x"81",
           686 => x"88",
           687 => x"81",
           688 => x"f8",
           689 => x"81",
           690 => x"f8",
           691 => x"81",
           692 => x"fc",
           693 => x"2e",
           694 => x"f8",
           695 => x"05",
           696 => x"f8",
           697 => x"05",
           698 => x"d4",
           699 => x"08",
           700 => x"c8",
           701 => x"3d",
           702 => x"d4",
           703 => x"f8",
           704 => x"81",
           705 => x"fb",
           706 => x"0b",
           707 => x"08",
           708 => x"81",
           709 => x"88",
           710 => x"25",
           711 => x"f8",
           712 => x"05",
           713 => x"f8",
           714 => x"05",
           715 => x"81",
           716 => x"fc",
           717 => x"f8",
           718 => x"05",
           719 => x"90",
           720 => x"d4",
           721 => x"08",
           722 => x"d4",
           723 => x"0c",
           724 => x"f8",
           725 => x"05",
           726 => x"f8",
           727 => x"05",
           728 => x"3f",
           729 => x"08",
           730 => x"d4",
           731 => x"0c",
           732 => x"d4",
           733 => x"08",
           734 => x"38",
           735 => x"08",
           736 => x"30",
           737 => x"08",
           738 => x"81",
           739 => x"f8",
           740 => x"81",
           741 => x"54",
           742 => x"81",
           743 => x"04",
           744 => x"08",
           745 => x"d4",
           746 => x"0d",
           747 => x"f8",
           748 => x"05",
           749 => x"81",
           750 => x"f8",
           751 => x"f8",
           752 => x"05",
           753 => x"d4",
           754 => x"08",
           755 => x"81",
           756 => x"fc",
           757 => x"2e",
           758 => x"0b",
           759 => x"08",
           760 => x"24",
           761 => x"f8",
           762 => x"05",
           763 => x"f8",
           764 => x"05",
           765 => x"d4",
           766 => x"08",
           767 => x"d4",
           768 => x"0c",
           769 => x"81",
           770 => x"fc",
           771 => x"2e",
           772 => x"81",
           773 => x"8c",
           774 => x"f8",
           775 => x"05",
           776 => x"38",
           777 => x"08",
           778 => x"81",
           779 => x"8c",
           780 => x"81",
           781 => x"88",
           782 => x"f8",
           783 => x"05",
           784 => x"d4",
           785 => x"08",
           786 => x"d4",
           787 => x"0c",
           788 => x"08",
           789 => x"81",
           790 => x"d4",
           791 => x"0c",
           792 => x"08",
           793 => x"81",
           794 => x"d4",
           795 => x"0c",
           796 => x"81",
           797 => x"90",
           798 => x"2e",
           799 => x"f8",
           800 => x"05",
           801 => x"f8",
           802 => x"05",
           803 => x"39",
           804 => x"08",
           805 => x"70",
           806 => x"08",
           807 => x"51",
           808 => x"08",
           809 => x"81",
           810 => x"85",
           811 => x"f8",
           812 => x"fc",
           813 => x"70",
           814 => x"55",
           815 => x"72",
           816 => x"72",
           817 => x"06",
           818 => x"2e",
           819 => x"12",
           820 => x"2e",
           821 => x"70",
           822 => x"33",
           823 => x"05",
           824 => x"12",
           825 => x"2e",
           826 => x"ea",
           827 => x"f8",
           828 => x"3d",
           829 => x"51",
           830 => x"05",
           831 => x"70",
           832 => x"0c",
           833 => x"05",
           834 => x"70",
           835 => x"0c",
           836 => x"05",
           837 => x"70",
           838 => x"0c",
           839 => x"05",
           840 => x"70",
           841 => x"0c",
           842 => x"71",
           843 => x"38",
           844 => x"95",
           845 => x"84",
           846 => x"71",
           847 => x"53",
           848 => x"52",
           849 => x"ed",
           850 => x"ff",
           851 => x"3d",
           852 => x"71",
           853 => x"9f",
           854 => x"55",
           855 => x"72",
           856 => x"74",
           857 => x"70",
           858 => x"38",
           859 => x"71",
           860 => x"38",
           861 => x"81",
           862 => x"ff",
           863 => x"ff",
           864 => x"06",
           865 => x"81",
           866 => x"86",
           867 => x"74",
           868 => x"75",
           869 => x"90",
           870 => x"54",
           871 => x"27",
           872 => x"71",
           873 => x"53",
           874 => x"70",
           875 => x"0c",
           876 => x"84",
           877 => x"72",
           878 => x"05",
           879 => x"12",
           880 => x"26",
           881 => x"72",
           882 => x"72",
           883 => x"05",
           884 => x"12",
           885 => x"26",
           886 => x"53",
           887 => x"fc",
           888 => x"70",
           889 => x"07",
           890 => x"54",
           891 => x"80",
           892 => x"70",
           893 => x"70",
           894 => x"ff",
           895 => x"f8",
           896 => x"80",
           897 => x"53",
           898 => x"a6",
           899 => x"72",
           900 => x"05",
           901 => x"08",
           902 => x"f7",
           903 => x"13",
           904 => x"84",
           905 => x"06",
           906 => x"53",
           907 => x"2e",
           908 => x"52",
           909 => x"05",
           910 => x"70",
           911 => x"05",
           912 => x"f0",
           913 => x"f8",
           914 => x"3d",
           915 => x"3d",
           916 => x"71",
           917 => x"55",
           918 => x"38",
           919 => x"70",
           920 => x"fd",
           921 => x"70",
           922 => x"81",
           923 => x"51",
           924 => x"9d",
           925 => x"70",
           926 => x"f7",
           927 => x"12",
           928 => x"84",
           929 => x"06",
           930 => x"53",
           931 => x"e5",
           932 => x"71",
           933 => x"80",
           934 => x"81",
           935 => x"52",
           936 => x"38",
           937 => x"81",
           938 => x"85",
           939 => x"fa",
           940 => x"7a",
           941 => x"55",
           942 => x"80",
           943 => x"38",
           944 => x"83",
           945 => x"80",
           946 => x"38",
           947 => x"72",
           948 => x"38",
           949 => x"33",
           950 => x"71",
           951 => x"06",
           952 => x"80",
           953 => x"38",
           954 => x"06",
           955 => x"2e",
           956 => x"81",
           957 => x"ff",
           958 => x"52",
           959 => x"09",
           960 => x"38",
           961 => x"33",
           962 => x"81",
           963 => x"81",
           964 => x"71",
           965 => x"52",
           966 => x"c8",
           967 => x"0d",
           968 => x"57",
           969 => x"27",
           970 => x"08",
           971 => x"88",
           972 => x"55",
           973 => x"39",
           974 => x"72",
           975 => x"38",
           976 => x"09",
           977 => x"ff",
           978 => x"f8",
           979 => x"80",
           980 => x"51",
           981 => x"84",
           982 => x"57",
           983 => x"27",
           984 => x"08",
           985 => x"d0",
           986 => x"55",
           987 => x"39",
           988 => x"f8",
           989 => x"3d",
           990 => x"3d",
           991 => x"83",
           992 => x"2b",
           993 => x"3f",
           994 => x"08",
           995 => x"72",
           996 => x"54",
           997 => x"25",
           998 => x"81",
           999 => x"84",
          1000 => x"fb",
          1001 => x"70",
          1002 => x"53",
          1003 => x"2e",
          1004 => x"71",
          1005 => x"a0",
          1006 => x"06",
          1007 => x"12",
          1008 => x"71",
          1009 => x"81",
          1010 => x"73",
          1011 => x"ff",
          1012 => x"55",
          1013 => x"83",
          1014 => x"70",
          1015 => x"38",
          1016 => x"73",
          1017 => x"51",
          1018 => x"09",
          1019 => x"38",
          1020 => x"81",
          1021 => x"72",
          1022 => x"51",
          1023 => x"c8",
          1024 => x"0d",
          1025 => x"0d",
          1026 => x"08",
          1027 => x"38",
          1028 => x"05",
          1029 => x"9f",
          1030 => x"f8",
          1031 => x"38",
          1032 => x"39",
          1033 => x"81",
          1034 => x"86",
          1035 => x"fc",
          1036 => x"82",
          1037 => x"05",
          1038 => x"52",
          1039 => x"81",
          1040 => x"13",
          1041 => x"51",
          1042 => x"9e",
          1043 => x"38",
          1044 => x"51",
          1045 => x"97",
          1046 => x"38",
          1047 => x"51",
          1048 => x"bb",
          1049 => x"38",
          1050 => x"51",
          1051 => x"bb",
          1052 => x"38",
          1053 => x"55",
          1054 => x"87",
          1055 => x"d9",
          1056 => x"22",
          1057 => x"73",
          1058 => x"80",
          1059 => x"0b",
          1060 => x"9c",
          1061 => x"87",
          1062 => x"0c",
          1063 => x"87",
          1064 => x"0c",
          1065 => x"87",
          1066 => x"0c",
          1067 => x"87",
          1068 => x"0c",
          1069 => x"87",
          1070 => x"0c",
          1071 => x"87",
          1072 => x"0c",
          1073 => x"98",
          1074 => x"87",
          1075 => x"0c",
          1076 => x"c0",
          1077 => x"80",
          1078 => x"f8",
          1079 => x"3d",
          1080 => x"3d",
          1081 => x"87",
          1082 => x"5d",
          1083 => x"87",
          1084 => x"08",
          1085 => x"23",
          1086 => x"b8",
          1087 => x"82",
          1088 => x"c0",
          1089 => x"5a",
          1090 => x"34",
          1091 => x"b0",
          1092 => x"84",
          1093 => x"c0",
          1094 => x"5a",
          1095 => x"34",
          1096 => x"a8",
          1097 => x"86",
          1098 => x"c0",
          1099 => x"5c",
          1100 => x"23",
          1101 => x"a0",
          1102 => x"8a",
          1103 => x"7d",
          1104 => x"ff",
          1105 => x"7b",
          1106 => x"06",
          1107 => x"33",
          1108 => x"33",
          1109 => x"33",
          1110 => x"33",
          1111 => x"33",
          1112 => x"ff",
          1113 => x"81",
          1114 => x"98",
          1115 => x"3d",
          1116 => x"3d",
          1117 => x"05",
          1118 => x"70",
          1119 => x"52",
          1120 => x"0b",
          1121 => x"34",
          1122 => x"04",
          1123 => x"77",
          1124 => x"f3",
          1125 => x"81",
          1126 => x"55",
          1127 => x"94",
          1128 => x"80",
          1129 => x"87",
          1130 => x"51",
          1131 => x"96",
          1132 => x"06",
          1133 => x"70",
          1134 => x"38",
          1135 => x"70",
          1136 => x"51",
          1137 => x"72",
          1138 => x"81",
          1139 => x"70",
          1140 => x"38",
          1141 => x"70",
          1142 => x"51",
          1143 => x"38",
          1144 => x"06",
          1145 => x"94",
          1146 => x"80",
          1147 => x"87",
          1148 => x"52",
          1149 => x"75",
          1150 => x"0c",
          1151 => x"04",
          1152 => x"02",
          1153 => x"0b",
          1154 => x"c0",
          1155 => x"ff",
          1156 => x"56",
          1157 => x"84",
          1158 => x"2e",
          1159 => x"c0",
          1160 => x"70",
          1161 => x"2a",
          1162 => x"53",
          1163 => x"80",
          1164 => x"71",
          1165 => x"81",
          1166 => x"70",
          1167 => x"81",
          1168 => x"06",
          1169 => x"80",
          1170 => x"71",
          1171 => x"81",
          1172 => x"70",
          1173 => x"73",
          1174 => x"51",
          1175 => x"80",
          1176 => x"2e",
          1177 => x"c0",
          1178 => x"75",
          1179 => x"3d",
          1180 => x"3d",
          1181 => x"80",
          1182 => x"81",
          1183 => x"53",
          1184 => x"2e",
          1185 => x"71",
          1186 => x"81",
          1187 => x"81",
          1188 => x"70",
          1189 => x"59",
          1190 => x"87",
          1191 => x"51",
          1192 => x"86",
          1193 => x"94",
          1194 => x"08",
          1195 => x"70",
          1196 => x"54",
          1197 => x"2e",
          1198 => x"91",
          1199 => x"06",
          1200 => x"d7",
          1201 => x"32",
          1202 => x"51",
          1203 => x"2e",
          1204 => x"93",
          1205 => x"06",
          1206 => x"ff",
          1207 => x"81",
          1208 => x"87",
          1209 => x"52",
          1210 => x"86",
          1211 => x"94",
          1212 => x"72",
          1213 => x"74",
          1214 => x"ff",
          1215 => x"57",
          1216 => x"38",
          1217 => x"c8",
          1218 => x"0d",
          1219 => x"0d",
          1220 => x"f3",
          1221 => x"81",
          1222 => x"52",
          1223 => x"84",
          1224 => x"2e",
          1225 => x"c0",
          1226 => x"70",
          1227 => x"2a",
          1228 => x"51",
          1229 => x"80",
          1230 => x"71",
          1231 => x"51",
          1232 => x"80",
          1233 => x"2e",
          1234 => x"c0",
          1235 => x"71",
          1236 => x"ff",
          1237 => x"c8",
          1238 => x"3d",
          1239 => x"3d",
          1240 => x"81",
          1241 => x"70",
          1242 => x"52",
          1243 => x"94",
          1244 => x"80",
          1245 => x"87",
          1246 => x"52",
          1247 => x"82",
          1248 => x"06",
          1249 => x"ff",
          1250 => x"2e",
          1251 => x"81",
          1252 => x"87",
          1253 => x"52",
          1254 => x"86",
          1255 => x"94",
          1256 => x"08",
          1257 => x"70",
          1258 => x"53",
          1259 => x"f8",
          1260 => x"3d",
          1261 => x"3d",
          1262 => x"9e",
          1263 => x"9c",
          1264 => x"51",
          1265 => x"2e",
          1266 => x"87",
          1267 => x"08",
          1268 => x"0c",
          1269 => x"a8",
          1270 => x"c8",
          1271 => x"9e",
          1272 => x"f3",
          1273 => x"c0",
          1274 => x"81",
          1275 => x"87",
          1276 => x"08",
          1277 => x"0c",
          1278 => x"a0",
          1279 => x"d8",
          1280 => x"9e",
          1281 => x"f3",
          1282 => x"c0",
          1283 => x"81",
          1284 => x"87",
          1285 => x"08",
          1286 => x"0c",
          1287 => x"b8",
          1288 => x"e8",
          1289 => x"9e",
          1290 => x"f3",
          1291 => x"c0",
          1292 => x"81",
          1293 => x"87",
          1294 => x"08",
          1295 => x"0c",
          1296 => x"80",
          1297 => x"81",
          1298 => x"87",
          1299 => x"08",
          1300 => x"0c",
          1301 => x"88",
          1302 => x"80",
          1303 => x"9e",
          1304 => x"f4",
          1305 => x"0b",
          1306 => x"34",
          1307 => x"c0",
          1308 => x"70",
          1309 => x"06",
          1310 => x"70",
          1311 => x"38",
          1312 => x"81",
          1313 => x"80",
          1314 => x"9e",
          1315 => x"88",
          1316 => x"51",
          1317 => x"80",
          1318 => x"81",
          1319 => x"f4",
          1320 => x"0b",
          1321 => x"90",
          1322 => x"80",
          1323 => x"52",
          1324 => x"2e",
          1325 => x"52",
          1326 => x"8b",
          1327 => x"87",
          1328 => x"08",
          1329 => x"80",
          1330 => x"52",
          1331 => x"83",
          1332 => x"71",
          1333 => x"34",
          1334 => x"c0",
          1335 => x"70",
          1336 => x"06",
          1337 => x"70",
          1338 => x"38",
          1339 => x"81",
          1340 => x"80",
          1341 => x"9e",
          1342 => x"90",
          1343 => x"51",
          1344 => x"80",
          1345 => x"81",
          1346 => x"f4",
          1347 => x"0b",
          1348 => x"90",
          1349 => x"80",
          1350 => x"52",
          1351 => x"2e",
          1352 => x"52",
          1353 => x"8f",
          1354 => x"87",
          1355 => x"08",
          1356 => x"80",
          1357 => x"52",
          1358 => x"83",
          1359 => x"71",
          1360 => x"34",
          1361 => x"c0",
          1362 => x"70",
          1363 => x"06",
          1364 => x"70",
          1365 => x"38",
          1366 => x"81",
          1367 => x"80",
          1368 => x"9e",
          1369 => x"80",
          1370 => x"51",
          1371 => x"80",
          1372 => x"81",
          1373 => x"f4",
          1374 => x"0b",
          1375 => x"90",
          1376 => x"80",
          1377 => x"52",
          1378 => x"83",
          1379 => x"71",
          1380 => x"34",
          1381 => x"90",
          1382 => x"80",
          1383 => x"2a",
          1384 => x"70",
          1385 => x"34",
          1386 => x"c0",
          1387 => x"70",
          1388 => x"51",
          1389 => x"80",
          1390 => x"81",
          1391 => x"f4",
          1392 => x"c0",
          1393 => x"70",
          1394 => x"70",
          1395 => x"51",
          1396 => x"f4",
          1397 => x"0b",
          1398 => x"90",
          1399 => x"06",
          1400 => x"70",
          1401 => x"38",
          1402 => x"81",
          1403 => x"87",
          1404 => x"08",
          1405 => x"51",
          1406 => x"f4",
          1407 => x"3d",
          1408 => x"3d",
          1409 => x"e8",
          1410 => x"3f",
          1411 => x"33",
          1412 => x"2e",
          1413 => x"dd",
          1414 => x"c9",
          1415 => x"90",
          1416 => x"3f",
          1417 => x"33",
          1418 => x"2e",
          1419 => x"f3",
          1420 => x"f3",
          1421 => x"54",
          1422 => x"a8",
          1423 => x"3f",
          1424 => x"33",
          1425 => x"2e",
          1426 => x"f3",
          1427 => x"f3",
          1428 => x"54",
          1429 => x"c4",
          1430 => x"3f",
          1431 => x"33",
          1432 => x"2e",
          1433 => x"f3",
          1434 => x"f3",
          1435 => x"54",
          1436 => x"e0",
          1437 => x"3f",
          1438 => x"33",
          1439 => x"2e",
          1440 => x"f3",
          1441 => x"f3",
          1442 => x"54",
          1443 => x"fc",
          1444 => x"3f",
          1445 => x"33",
          1446 => x"2e",
          1447 => x"f3",
          1448 => x"f3",
          1449 => x"54",
          1450 => x"98",
          1451 => x"3f",
          1452 => x"33",
          1453 => x"2e",
          1454 => x"f4",
          1455 => x"81",
          1456 => x"8e",
          1457 => x"f4",
          1458 => x"73",
          1459 => x"38",
          1460 => x"33",
          1461 => x"d4",
          1462 => x"3f",
          1463 => x"33",
          1464 => x"2e",
          1465 => x"f4",
          1466 => x"81",
          1467 => x"8d",
          1468 => x"f4",
          1469 => x"73",
          1470 => x"38",
          1471 => x"51",
          1472 => x"81",
          1473 => x"54",
          1474 => x"88",
          1475 => x"a8",
          1476 => x"3f",
          1477 => x"33",
          1478 => x"2e",
          1479 => x"e0",
          1480 => x"c1",
          1481 => x"91",
          1482 => x"80",
          1483 => x"81",
          1484 => x"87",
          1485 => x"f4",
          1486 => x"73",
          1487 => x"38",
          1488 => x"51",
          1489 => x"81",
          1490 => x"87",
          1491 => x"f3",
          1492 => x"81",
          1493 => x"8c",
          1494 => x"f3",
          1495 => x"81",
          1496 => x"8c",
          1497 => x"f3",
          1498 => x"81",
          1499 => x"8c",
          1500 => x"e1",
          1501 => x"ed",
          1502 => x"f8",
          1503 => x"e1",
          1504 => x"c5",
          1505 => x"fc",
          1506 => x"84",
          1507 => x"51",
          1508 => x"81",
          1509 => x"bd",
          1510 => x"76",
          1511 => x"54",
          1512 => x"08",
          1513 => x"8c",
          1514 => x"3f",
          1515 => x"33",
          1516 => x"2e",
          1517 => x"f4",
          1518 => x"bd",
          1519 => x"75",
          1520 => x"3f",
          1521 => x"08",
          1522 => x"29",
          1523 => x"54",
          1524 => x"c8",
          1525 => x"e2",
          1526 => x"ed",
          1527 => x"8a",
          1528 => x"80",
          1529 => x"81",
          1530 => x"56",
          1531 => x"52",
          1532 => x"b8",
          1533 => x"c8",
          1534 => x"c0",
          1535 => x"31",
          1536 => x"f8",
          1537 => x"81",
          1538 => x"8b",
          1539 => x"f1",
          1540 => x"d1",
          1541 => x"0d",
          1542 => x"0d",
          1543 => x"33",
          1544 => x"71",
          1545 => x"38",
          1546 => x"81",
          1547 => x"52",
          1548 => x"81",
          1549 => x"9d",
          1550 => x"98",
          1551 => x"81",
          1552 => x"91",
          1553 => x"a8",
          1554 => x"81",
          1555 => x"85",
          1556 => x"b4",
          1557 => x"3f",
          1558 => x"04",
          1559 => x"0c",
          1560 => x"87",
          1561 => x"0c",
          1562 => x"9c",
          1563 => x"96",
          1564 => x"fe",
          1565 => x"f8",
          1566 => x"38",
          1567 => x"0b",
          1568 => x"0c",
          1569 => x"08",
          1570 => x"52",
          1571 => x"83",
          1572 => x"88",
          1573 => x"f8",
          1574 => x"53",
          1575 => x"c8",
          1576 => x"0d",
          1577 => x"0d",
          1578 => x"12",
          1579 => x"90",
          1580 => x"15",
          1581 => x"5e",
          1582 => x"59",
          1583 => x"77",
          1584 => x"75",
          1585 => x"08",
          1586 => x"71",
          1587 => x"31",
          1588 => x"80",
          1589 => x"84",
          1590 => x"8c",
          1591 => x"88",
          1592 => x"8c",
          1593 => x"88",
          1594 => x"90",
          1595 => x"94",
          1596 => x"94",
          1597 => x"90",
          1598 => x"39",
          1599 => x"73",
          1600 => x"74",
          1601 => x"77",
          1602 => x"0c",
          1603 => x"04",
          1604 => x"76",
          1605 => x"88",
          1606 => x"53",
          1607 => x"81",
          1608 => x"06",
          1609 => x"12",
          1610 => x"52",
          1611 => x"2e",
          1612 => x"94",
          1613 => x"08",
          1614 => x"0c",
          1615 => x"0c",
          1616 => x"0c",
          1617 => x"39",
          1618 => x"81",
          1619 => x"90",
          1620 => x"f4",
          1621 => x"14",
          1622 => x"f4",
          1623 => x"13",
          1624 => x"12",
          1625 => x"08",
          1626 => x"81",
          1627 => x"84",
          1628 => x"14",
          1629 => x"74",
          1630 => x"06",
          1631 => x"14",
          1632 => x"14",
          1633 => x"08",
          1634 => x"70",
          1635 => x"52",
          1636 => x"8c",
          1637 => x"15",
          1638 => x"13",
          1639 => x"12",
          1640 => x"f8",
          1641 => x"3d",
          1642 => x"3d",
          1643 => x"55",
          1644 => x"2e",
          1645 => x"9f",
          1646 => x"81",
          1647 => x"57",
          1648 => x"82",
          1649 => x"84",
          1650 => x"27",
          1651 => x"90",
          1652 => x"ed",
          1653 => x"ff",
          1654 => x"80",
          1655 => x"58",
          1656 => x"81",
          1657 => x"81",
          1658 => x"30",
          1659 => x"c8",
          1660 => x"25",
          1661 => x"08",
          1662 => x"70",
          1663 => x"25",
          1664 => x"58",
          1665 => x"56",
          1666 => x"74",
          1667 => x"06",
          1668 => x"88",
          1669 => x"75",
          1670 => x"39",
          1671 => x"f8",
          1672 => x"77",
          1673 => x"08",
          1674 => x"81",
          1675 => x"53",
          1676 => x"2e",
          1677 => x"73",
          1678 => x"8c",
          1679 => x"f0",
          1680 => x"08",
          1681 => x"72",
          1682 => x"75",
          1683 => x"88",
          1684 => x"8c",
          1685 => x"75",
          1686 => x"3f",
          1687 => x"f8",
          1688 => x"fc",
          1689 => x"f8",
          1690 => x"73",
          1691 => x"0c",
          1692 => x"04",
          1693 => x"73",
          1694 => x"2e",
          1695 => x"12",
          1696 => x"3f",
          1697 => x"04",
          1698 => x"02",
          1699 => x"53",
          1700 => x"09",
          1701 => x"38",
          1702 => x"3f",
          1703 => x"08",
          1704 => x"2e",
          1705 => x"72",
          1706 => x"e4",
          1707 => x"81",
          1708 => x"8f",
          1709 => x"dc",
          1710 => x"80",
          1711 => x"72",
          1712 => x"84",
          1713 => x"fe",
          1714 => x"97",
          1715 => x"f8",
          1716 => x"81",
          1717 => x"54",
          1718 => x"3f",
          1719 => x"dc",
          1720 => x"0d",
          1721 => x"0d",
          1722 => x"33",
          1723 => x"06",
          1724 => x"80",
          1725 => x"72",
          1726 => x"51",
          1727 => x"ff",
          1728 => x"39",
          1729 => x"04",
          1730 => x"77",
          1731 => x"08",
          1732 => x"dc",
          1733 => x"73",
          1734 => x"ff",
          1735 => x"71",
          1736 => x"38",
          1737 => x"06",
          1738 => x"54",
          1739 => x"e7",
          1740 => x"f8",
          1741 => x"3d",
          1742 => x"3d",
          1743 => x"59",
          1744 => x"81",
          1745 => x"56",
          1746 => x"84",
          1747 => x"a5",
          1748 => x"06",
          1749 => x"80",
          1750 => x"81",
          1751 => x"58",
          1752 => x"b0",
          1753 => x"06",
          1754 => x"5a",
          1755 => x"ad",
          1756 => x"06",
          1757 => x"5a",
          1758 => x"05",
          1759 => x"75",
          1760 => x"81",
          1761 => x"77",
          1762 => x"08",
          1763 => x"05",
          1764 => x"5d",
          1765 => x"39",
          1766 => x"72",
          1767 => x"38",
          1768 => x"7b",
          1769 => x"05",
          1770 => x"70",
          1771 => x"33",
          1772 => x"39",
          1773 => x"32",
          1774 => x"72",
          1775 => x"78",
          1776 => x"70",
          1777 => x"07",
          1778 => x"07",
          1779 => x"51",
          1780 => x"80",
          1781 => x"79",
          1782 => x"70",
          1783 => x"33",
          1784 => x"80",
          1785 => x"38",
          1786 => x"e0",
          1787 => x"38",
          1788 => x"81",
          1789 => x"53",
          1790 => x"2e",
          1791 => x"73",
          1792 => x"a2",
          1793 => x"c3",
          1794 => x"38",
          1795 => x"24",
          1796 => x"80",
          1797 => x"8c",
          1798 => x"39",
          1799 => x"2e",
          1800 => x"81",
          1801 => x"80",
          1802 => x"80",
          1803 => x"d5",
          1804 => x"73",
          1805 => x"8e",
          1806 => x"39",
          1807 => x"2e",
          1808 => x"80",
          1809 => x"84",
          1810 => x"56",
          1811 => x"74",
          1812 => x"72",
          1813 => x"38",
          1814 => x"15",
          1815 => x"54",
          1816 => x"38",
          1817 => x"56",
          1818 => x"81",
          1819 => x"72",
          1820 => x"38",
          1821 => x"90",
          1822 => x"06",
          1823 => x"2e",
          1824 => x"51",
          1825 => x"74",
          1826 => x"53",
          1827 => x"fd",
          1828 => x"51",
          1829 => x"ef",
          1830 => x"19",
          1831 => x"53",
          1832 => x"39",
          1833 => x"39",
          1834 => x"39",
          1835 => x"39",
          1836 => x"39",
          1837 => x"d0",
          1838 => x"39",
          1839 => x"70",
          1840 => x"53",
          1841 => x"88",
          1842 => x"19",
          1843 => x"39",
          1844 => x"54",
          1845 => x"74",
          1846 => x"70",
          1847 => x"07",
          1848 => x"55",
          1849 => x"80",
          1850 => x"72",
          1851 => x"38",
          1852 => x"90",
          1853 => x"80",
          1854 => x"5e",
          1855 => x"74",
          1856 => x"3f",
          1857 => x"08",
          1858 => x"7c",
          1859 => x"54",
          1860 => x"81",
          1861 => x"55",
          1862 => x"92",
          1863 => x"53",
          1864 => x"2e",
          1865 => x"14",
          1866 => x"ff",
          1867 => x"14",
          1868 => x"70",
          1869 => x"34",
          1870 => x"30",
          1871 => x"9f",
          1872 => x"57",
          1873 => x"85",
          1874 => x"b1",
          1875 => x"2a",
          1876 => x"51",
          1877 => x"2e",
          1878 => x"3d",
          1879 => x"05",
          1880 => x"34",
          1881 => x"76",
          1882 => x"54",
          1883 => x"72",
          1884 => x"54",
          1885 => x"70",
          1886 => x"56",
          1887 => x"81",
          1888 => x"7b",
          1889 => x"73",
          1890 => x"3f",
          1891 => x"53",
          1892 => x"74",
          1893 => x"53",
          1894 => x"eb",
          1895 => x"77",
          1896 => x"53",
          1897 => x"14",
          1898 => x"54",
          1899 => x"3f",
          1900 => x"74",
          1901 => x"53",
          1902 => x"fb",
          1903 => x"51",
          1904 => x"ef",
          1905 => x"0d",
          1906 => x"0d",
          1907 => x"70",
          1908 => x"08",
          1909 => x"51",
          1910 => x"85",
          1911 => x"fe",
          1912 => x"81",
          1913 => x"85",
          1914 => x"52",
          1915 => x"ca",
          1916 => x"e4",
          1917 => x"73",
          1918 => x"81",
          1919 => x"84",
          1920 => x"fd",
          1921 => x"f8",
          1922 => x"81",
          1923 => x"87",
          1924 => x"53",
          1925 => x"fa",
          1926 => x"81",
          1927 => x"85",
          1928 => x"fb",
          1929 => x"79",
          1930 => x"08",
          1931 => x"57",
          1932 => x"71",
          1933 => x"e0",
          1934 => x"e0",
          1935 => x"2d",
          1936 => x"08",
          1937 => x"53",
          1938 => x"80",
          1939 => x"8d",
          1940 => x"72",
          1941 => x"30",
          1942 => x"51",
          1943 => x"80",
          1944 => x"71",
          1945 => x"38",
          1946 => x"97",
          1947 => x"25",
          1948 => x"16",
          1949 => x"25",
          1950 => x"14",
          1951 => x"34",
          1952 => x"72",
          1953 => x"3f",
          1954 => x"73",
          1955 => x"72",
          1956 => x"f7",
          1957 => x"53",
          1958 => x"c8",
          1959 => x"0d",
          1960 => x"0d",
          1961 => x"08",
          1962 => x"e0",
          1963 => x"76",
          1964 => x"ef",
          1965 => x"f8",
          1966 => x"3d",
          1967 => x"3d",
          1968 => x"5a",
          1969 => x"7a",
          1970 => x"08",
          1971 => x"53",
          1972 => x"09",
          1973 => x"38",
          1974 => x"0c",
          1975 => x"ad",
          1976 => x"06",
          1977 => x"76",
          1978 => x"0c",
          1979 => x"33",
          1980 => x"73",
          1981 => x"81",
          1982 => x"38",
          1983 => x"05",
          1984 => x"08",
          1985 => x"53",
          1986 => x"2e",
          1987 => x"57",
          1988 => x"2e",
          1989 => x"39",
          1990 => x"13",
          1991 => x"08",
          1992 => x"53",
          1993 => x"55",
          1994 => x"80",
          1995 => x"14",
          1996 => x"88",
          1997 => x"27",
          1998 => x"eb",
          1999 => x"53",
          2000 => x"89",
          2001 => x"38",
          2002 => x"55",
          2003 => x"8a",
          2004 => x"a0",
          2005 => x"c2",
          2006 => x"74",
          2007 => x"e0",
          2008 => x"ff",
          2009 => x"d0",
          2010 => x"ff",
          2011 => x"90",
          2012 => x"38",
          2013 => x"81",
          2014 => x"53",
          2015 => x"ca",
          2016 => x"27",
          2017 => x"77",
          2018 => x"08",
          2019 => x"0c",
          2020 => x"33",
          2021 => x"ff",
          2022 => x"80",
          2023 => x"74",
          2024 => x"79",
          2025 => x"74",
          2026 => x"0c",
          2027 => x"04",
          2028 => x"7a",
          2029 => x"80",
          2030 => x"58",
          2031 => x"33",
          2032 => x"a0",
          2033 => x"06",
          2034 => x"13",
          2035 => x"39",
          2036 => x"09",
          2037 => x"38",
          2038 => x"11",
          2039 => x"08",
          2040 => x"54",
          2041 => x"2e",
          2042 => x"80",
          2043 => x"08",
          2044 => x"0c",
          2045 => x"33",
          2046 => x"80",
          2047 => x"38",
          2048 => x"80",
          2049 => x"38",
          2050 => x"57",
          2051 => x"0c",
          2052 => x"33",
          2053 => x"39",
          2054 => x"74",
          2055 => x"38",
          2056 => x"80",
          2057 => x"89",
          2058 => x"38",
          2059 => x"d0",
          2060 => x"55",
          2061 => x"80",
          2062 => x"39",
          2063 => x"d9",
          2064 => x"80",
          2065 => x"27",
          2066 => x"80",
          2067 => x"89",
          2068 => x"70",
          2069 => x"55",
          2070 => x"70",
          2071 => x"55",
          2072 => x"27",
          2073 => x"14",
          2074 => x"06",
          2075 => x"74",
          2076 => x"73",
          2077 => x"38",
          2078 => x"14",
          2079 => x"05",
          2080 => x"08",
          2081 => x"54",
          2082 => x"39",
          2083 => x"84",
          2084 => x"55",
          2085 => x"81",
          2086 => x"f8",
          2087 => x"3d",
          2088 => x"3d",
          2089 => x"2b",
          2090 => x"79",
          2091 => x"98",
          2092 => x"13",
          2093 => x"51",
          2094 => x"51",
          2095 => x"81",
          2096 => x"33",
          2097 => x"74",
          2098 => x"81",
          2099 => x"08",
          2100 => x"05",
          2101 => x"71",
          2102 => x"52",
          2103 => x"09",
          2104 => x"38",
          2105 => x"81",
          2106 => x"85",
          2107 => x"fc",
          2108 => x"02",
          2109 => x"05",
          2110 => x"54",
          2111 => x"80",
          2112 => x"88",
          2113 => x"3f",
          2114 => x"fc",
          2115 => x"f2",
          2116 => x"33",
          2117 => x"71",
          2118 => x"81",
          2119 => x"de",
          2120 => x"f3",
          2121 => x"73",
          2122 => x"0d",
          2123 => x"0d",
          2124 => x"05",
          2125 => x"02",
          2126 => x"05",
          2127 => x"94",
          2128 => x"29",
          2129 => x"05",
          2130 => x"59",
          2131 => x"59",
          2132 => x"86",
          2133 => x"f2",
          2134 => x"f5",
          2135 => x"84",
          2136 => x"bc",
          2137 => x"70",
          2138 => x"5a",
          2139 => x"81",
          2140 => x"75",
          2141 => x"94",
          2142 => x"29",
          2143 => x"05",
          2144 => x"56",
          2145 => x"2e",
          2146 => x"53",
          2147 => x"51",
          2148 => x"81",
          2149 => x"81",
          2150 => x"81",
          2151 => x"74",
          2152 => x"55",
          2153 => x"87",
          2154 => x"81",
          2155 => x"77",
          2156 => x"38",
          2157 => x"08",
          2158 => x"2e",
          2159 => x"f5",
          2160 => x"74",
          2161 => x"3d",
          2162 => x"76",
          2163 => x"75",
          2164 => x"91",
          2165 => x"90",
          2166 => x"51",
          2167 => x"3f",
          2168 => x"08",
          2169 => x"ee",
          2170 => x"0d",
          2171 => x"0d",
          2172 => x"52",
          2173 => x"08",
          2174 => x"87",
          2175 => x"c8",
          2176 => x"38",
          2177 => x"08",
          2178 => x"52",
          2179 => x"52",
          2180 => x"d5",
          2181 => x"c8",
          2182 => x"b8",
          2183 => x"d8",
          2184 => x"f8",
          2185 => x"80",
          2186 => x"c8",
          2187 => x"38",
          2188 => x"08",
          2189 => x"17",
          2190 => x"74",
          2191 => x"76",
          2192 => x"81",
          2193 => x"57",
          2194 => x"74",
          2195 => x"81",
          2196 => x"38",
          2197 => x"04",
          2198 => x"aa",
          2199 => x"3d",
          2200 => x"81",
          2201 => x"80",
          2202 => x"90",
          2203 => x"d1",
          2204 => x"f8",
          2205 => x"91",
          2206 => x"81",
          2207 => x"54",
          2208 => x"52",
          2209 => x"52",
          2210 => x"dd",
          2211 => x"c8",
          2212 => x"a4",
          2213 => x"d7",
          2214 => x"f8",
          2215 => x"18",
          2216 => x"0b",
          2217 => x"08",
          2218 => x"81",
          2219 => x"ff",
          2220 => x"55",
          2221 => x"34",
          2222 => x"30",
          2223 => x"9f",
          2224 => x"55",
          2225 => x"85",
          2226 => x"ad",
          2227 => x"90",
          2228 => x"08",
          2229 => x"d0",
          2230 => x"f8",
          2231 => x"2e",
          2232 => x"e3",
          2233 => x"fd",
          2234 => x"2e",
          2235 => x"99",
          2236 => x"79",
          2237 => x"3f",
          2238 => x"d2",
          2239 => x"08",
          2240 => x"c8",
          2241 => x"80",
          2242 => x"f8",
          2243 => x"3d",
          2244 => x"3d",
          2245 => x"71",
          2246 => x"33",
          2247 => x"58",
          2248 => x"09",
          2249 => x"38",
          2250 => x"05",
          2251 => x"27",
          2252 => x"17",
          2253 => x"71",
          2254 => x"55",
          2255 => x"09",
          2256 => x"38",
          2257 => x"ea",
          2258 => x"73",
          2259 => x"f5",
          2260 => x"08",
          2261 => x"f6",
          2262 => x"c8",
          2263 => x"52",
          2264 => x"d6",
          2265 => x"f8",
          2266 => x"c4",
          2267 => x"33",
          2268 => x"2e",
          2269 => x"82",
          2270 => x"b4",
          2271 => x"3f",
          2272 => x"1a",
          2273 => x"fc",
          2274 => x"05",
          2275 => x"3f",
          2276 => x"08",
          2277 => x"38",
          2278 => x"52",
          2279 => x"b8",
          2280 => x"c8",
          2281 => x"06",
          2282 => x"38",
          2283 => x"39",
          2284 => x"81",
          2285 => x"54",
          2286 => x"ff",
          2287 => x"54",
          2288 => x"c8",
          2289 => x"0d",
          2290 => x"0d",
          2291 => x"02",
          2292 => x"c3",
          2293 => x"5a",
          2294 => x"3d",
          2295 => x"94",
          2296 => x"f5",
          2297 => x"a3",
          2298 => x"8c",
          2299 => x"81",
          2300 => x"51",
          2301 => x"81",
          2302 => x"81",
          2303 => x"81",
          2304 => x"80",
          2305 => x"38",
          2306 => x"f4",
          2307 => x"81",
          2308 => x"51",
          2309 => x"81",
          2310 => x"80",
          2311 => x"81",
          2312 => x"f3",
          2313 => x"e3",
          2314 => x"90",
          2315 => x"f8",
          2316 => x"70",
          2317 => x"f6",
          2318 => x"f8",
          2319 => x"81",
          2320 => x"74",
          2321 => x"06",
          2322 => x"81",
          2323 => x"51",
          2324 => x"81",
          2325 => x"55",
          2326 => x"f8",
          2327 => x"9a",
          2328 => x"c8",
          2329 => x"70",
          2330 => x"80",
          2331 => x"53",
          2332 => x"06",
          2333 => x"f9",
          2334 => x"ff",
          2335 => x"06",
          2336 => x"87",
          2337 => x"81",
          2338 => x"8f",
          2339 => x"ce",
          2340 => x"c8",
          2341 => x"70",
          2342 => x"59",
          2343 => x"ee",
          2344 => x"ff",
          2345 => x"ec",
          2346 => x"2b",
          2347 => x"81",
          2348 => x"70",
          2349 => x"97",
          2350 => x"2c",
          2351 => x"29",
          2352 => x"05",
          2353 => x"70",
          2354 => x"51",
          2355 => x"51",
          2356 => x"81",
          2357 => x"2e",
          2358 => x"77",
          2359 => x"38",
          2360 => x"0a",
          2361 => x"0a",
          2362 => x"2c",
          2363 => x"75",
          2364 => x"38",
          2365 => x"52",
          2366 => x"a6",
          2367 => x"c8",
          2368 => x"06",
          2369 => x"2e",
          2370 => x"81",
          2371 => x"81",
          2372 => x"74",
          2373 => x"29",
          2374 => x"05",
          2375 => x"70",
          2376 => x"56",
          2377 => x"8a",
          2378 => x"76",
          2379 => x"77",
          2380 => x"3f",
          2381 => x"08",
          2382 => x"54",
          2383 => x"d3",
          2384 => x"75",
          2385 => x"ca",
          2386 => x"55",
          2387 => x"ec",
          2388 => x"2b",
          2389 => x"81",
          2390 => x"70",
          2391 => x"98",
          2392 => x"11",
          2393 => x"81",
          2394 => x"33",
          2395 => x"51",
          2396 => x"55",
          2397 => x"09",
          2398 => x"92",
          2399 => x"cc",
          2400 => x"0c",
          2401 => x"f8",
          2402 => x"0b",
          2403 => x"34",
          2404 => x"81",
          2405 => x"75",
          2406 => x"34",
          2407 => x"34",
          2408 => x"7e",
          2409 => x"26",
          2410 => x"73",
          2411 => x"dc",
          2412 => x"73",
          2413 => x"f8",
          2414 => x"73",
          2415 => x"cb",
          2416 => x"f0",
          2417 => x"75",
          2418 => x"74",
          2419 => x"98",
          2420 => x"73",
          2421 => x"38",
          2422 => x"73",
          2423 => x"34",
          2424 => x"0a",
          2425 => x"0a",
          2426 => x"2c",
          2427 => x"33",
          2428 => x"df",
          2429 => x"f4",
          2430 => x"56",
          2431 => x"f8",
          2432 => x"1a",
          2433 => x"33",
          2434 => x"f8",
          2435 => x"73",
          2436 => x"38",
          2437 => x"73",
          2438 => x"34",
          2439 => x"33",
          2440 => x"0a",
          2441 => x"0a",
          2442 => x"2c",
          2443 => x"33",
          2444 => x"56",
          2445 => x"a2",
          2446 => x"70",
          2447 => x"e8",
          2448 => x"81",
          2449 => x"81",
          2450 => x"70",
          2451 => x"f8",
          2452 => x"51",
          2453 => x"24",
          2454 => x"f8",
          2455 => x"98",
          2456 => x"2c",
          2457 => x"33",
          2458 => x"56",
          2459 => x"fc",
          2460 => x"51",
          2461 => x"74",
          2462 => x"29",
          2463 => x"05",
          2464 => x"81",
          2465 => x"56",
          2466 => x"75",
          2467 => x"fb",
          2468 => x"f8",
          2469 => x"81",
          2470 => x"55",
          2471 => x"fb",
          2472 => x"f8",
          2473 => x"05",
          2474 => x"f8",
          2475 => x"15",
          2476 => x"f8",
          2477 => x"51",
          2478 => x"81",
          2479 => x"70",
          2480 => x"98",
          2481 => x"f0",
          2482 => x"56",
          2483 => x"25",
          2484 => x"1a",
          2485 => x"33",
          2486 => x"33",
          2487 => x"3f",
          2488 => x"0a",
          2489 => x"0a",
          2490 => x"2c",
          2491 => x"33",
          2492 => x"75",
          2493 => x"38",
          2494 => x"8c",
          2495 => x"f4",
          2496 => x"2b",
          2497 => x"81",
          2498 => x"57",
          2499 => x"74",
          2500 => x"f7",
          2501 => x"e6",
          2502 => x"81",
          2503 => x"81",
          2504 => x"70",
          2505 => x"f8",
          2506 => x"51",
          2507 => x"25",
          2508 => x"d7",
          2509 => x"f0",
          2510 => x"54",
          2511 => x"8a",
          2512 => x"3f",
          2513 => x"52",
          2514 => x"c6",
          2515 => x"c8",
          2516 => x"06",
          2517 => x"38",
          2518 => x"33",
          2519 => x"2e",
          2520 => x"81",
          2521 => x"79",
          2522 => x"3f",
          2523 => x"80",
          2524 => x"b7",
          2525 => x"f4",
          2526 => x"80",
          2527 => x"38",
          2528 => x"84",
          2529 => x"f4",
          2530 => x"54",
          2531 => x"f4",
          2532 => x"ff",
          2533 => x"39",
          2534 => x"33",
          2535 => x"33",
          2536 => x"75",
          2537 => x"38",
          2538 => x"73",
          2539 => x"34",
          2540 => x"70",
          2541 => x"81",
          2542 => x"51",
          2543 => x"25",
          2544 => x"1a",
          2545 => x"33",
          2546 => x"33",
          2547 => x"3f",
          2548 => x"0a",
          2549 => x"0a",
          2550 => x"2c",
          2551 => x"33",
          2552 => x"75",
          2553 => x"38",
          2554 => x"9c",
          2555 => x"f4",
          2556 => x"2b",
          2557 => x"81",
          2558 => x"57",
          2559 => x"74",
          2560 => x"87",
          2561 => x"e4",
          2562 => x"81",
          2563 => x"81",
          2564 => x"70",
          2565 => x"f8",
          2566 => x"51",
          2567 => x"25",
          2568 => x"e7",
          2569 => x"f4",
          2570 => x"ff",
          2571 => x"f0",
          2572 => x"54",
          2573 => x"f8",
          2574 => x"14",
          2575 => x"f8",
          2576 => x"1a",
          2577 => x"54",
          2578 => x"81",
          2579 => x"70",
          2580 => x"81",
          2581 => x"58",
          2582 => x"75",
          2583 => x"f8",
          2584 => x"ae",
          2585 => x"88",
          2586 => x"80",
          2587 => x"74",
          2588 => x"3f",
          2589 => x"08",
          2590 => x"34",
          2591 => x"08",
          2592 => x"81",
          2593 => x"52",
          2594 => x"a7",
          2595 => x"81",
          2596 => x"84",
          2597 => x"bc",
          2598 => x"08",
          2599 => x"80",
          2600 => x"74",
          2601 => x"3f",
          2602 => x"08",
          2603 => x"34",
          2604 => x"08",
          2605 => x"81",
          2606 => x"52",
          2607 => x"f3",
          2608 => x"54",
          2609 => x"73",
          2610 => x"80",
          2611 => x"38",
          2612 => x"fa",
          2613 => x"39",
          2614 => x"09",
          2615 => x"38",
          2616 => x"08",
          2617 => x"2e",
          2618 => x"51",
          2619 => x"80",
          2620 => x"84",
          2621 => x"bc",
          2622 => x"08",
          2623 => x"80",
          2624 => x"74",
          2625 => x"3f",
          2626 => x"08",
          2627 => x"34",
          2628 => x"08",
          2629 => x"81",
          2630 => x"52",
          2631 => x"93",
          2632 => x"54",
          2633 => x"06",
          2634 => x"73",
          2635 => x"80",
          2636 => x"38",
          2637 => x"96",
          2638 => x"c8",
          2639 => x"f0",
          2640 => x"c8",
          2641 => x"06",
          2642 => x"74",
          2643 => x"c6",
          2644 => x"f8",
          2645 => x"f8",
          2646 => x"79",
          2647 => x"3f",
          2648 => x"81",
          2649 => x"70",
          2650 => x"81",
          2651 => x"59",
          2652 => x"77",
          2653 => x"38",
          2654 => x"73",
          2655 => x"34",
          2656 => x"33",
          2657 => x"80",
          2658 => x"39",
          2659 => x"33",
          2660 => x"2e",
          2661 => x"88",
          2662 => x"3f",
          2663 => x"33",
          2664 => x"73",
          2665 => x"34",
          2666 => x"80",
          2667 => x"f4",
          2668 => x"81",
          2669 => x"79",
          2670 => x"0c",
          2671 => x"04",
          2672 => x"02",
          2673 => x"51",
          2674 => x"72",
          2675 => x"81",
          2676 => x"33",
          2677 => x"f8",
          2678 => x"3d",
          2679 => x"3d",
          2680 => x"05",
          2681 => x"05",
          2682 => x"56",
          2683 => x"72",
          2684 => x"e0",
          2685 => x"2b",
          2686 => x"8c",
          2687 => x"88",
          2688 => x"2e",
          2689 => x"88",
          2690 => x"0c",
          2691 => x"8c",
          2692 => x"71",
          2693 => x"87",
          2694 => x"0c",
          2695 => x"08",
          2696 => x"51",
          2697 => x"2e",
          2698 => x"c0",
          2699 => x"51",
          2700 => x"71",
          2701 => x"80",
          2702 => x"92",
          2703 => x"98",
          2704 => x"70",
          2705 => x"38",
          2706 => x"b0",
          2707 => x"f5",
          2708 => x"51",
          2709 => x"c8",
          2710 => x"0d",
          2711 => x"0d",
          2712 => x"02",
          2713 => x"05",
          2714 => x"58",
          2715 => x"52",
          2716 => x"3f",
          2717 => x"08",
          2718 => x"54",
          2719 => x"be",
          2720 => x"75",
          2721 => x"c0",
          2722 => x"87",
          2723 => x"12",
          2724 => x"84",
          2725 => x"40",
          2726 => x"85",
          2727 => x"98",
          2728 => x"7d",
          2729 => x"0c",
          2730 => x"85",
          2731 => x"06",
          2732 => x"71",
          2733 => x"38",
          2734 => x"71",
          2735 => x"05",
          2736 => x"19",
          2737 => x"a2",
          2738 => x"71",
          2739 => x"38",
          2740 => x"83",
          2741 => x"38",
          2742 => x"8a",
          2743 => x"98",
          2744 => x"71",
          2745 => x"c0",
          2746 => x"52",
          2747 => x"87",
          2748 => x"80",
          2749 => x"81",
          2750 => x"c0",
          2751 => x"53",
          2752 => x"82",
          2753 => x"71",
          2754 => x"1a",
          2755 => x"84",
          2756 => x"19",
          2757 => x"06",
          2758 => x"79",
          2759 => x"38",
          2760 => x"80",
          2761 => x"87",
          2762 => x"26",
          2763 => x"73",
          2764 => x"06",
          2765 => x"2e",
          2766 => x"52",
          2767 => x"81",
          2768 => x"8f",
          2769 => x"f3",
          2770 => x"62",
          2771 => x"05",
          2772 => x"57",
          2773 => x"83",
          2774 => x"52",
          2775 => x"3f",
          2776 => x"08",
          2777 => x"54",
          2778 => x"2e",
          2779 => x"81",
          2780 => x"74",
          2781 => x"c0",
          2782 => x"87",
          2783 => x"12",
          2784 => x"84",
          2785 => x"5f",
          2786 => x"0b",
          2787 => x"8c",
          2788 => x"0c",
          2789 => x"80",
          2790 => x"70",
          2791 => x"81",
          2792 => x"54",
          2793 => x"8c",
          2794 => x"81",
          2795 => x"7c",
          2796 => x"58",
          2797 => x"70",
          2798 => x"52",
          2799 => x"8a",
          2800 => x"98",
          2801 => x"71",
          2802 => x"c0",
          2803 => x"52",
          2804 => x"87",
          2805 => x"80",
          2806 => x"81",
          2807 => x"c0",
          2808 => x"53",
          2809 => x"82",
          2810 => x"71",
          2811 => x"19",
          2812 => x"81",
          2813 => x"ff",
          2814 => x"19",
          2815 => x"78",
          2816 => x"38",
          2817 => x"80",
          2818 => x"87",
          2819 => x"26",
          2820 => x"73",
          2821 => x"06",
          2822 => x"2e",
          2823 => x"52",
          2824 => x"81",
          2825 => x"8f",
          2826 => x"fa",
          2827 => x"02",
          2828 => x"05",
          2829 => x"05",
          2830 => x"71",
          2831 => x"57",
          2832 => x"81",
          2833 => x"81",
          2834 => x"54",
          2835 => x"38",
          2836 => x"c0",
          2837 => x"81",
          2838 => x"2e",
          2839 => x"71",
          2840 => x"38",
          2841 => x"87",
          2842 => x"11",
          2843 => x"80",
          2844 => x"80",
          2845 => x"83",
          2846 => x"38",
          2847 => x"72",
          2848 => x"2a",
          2849 => x"51",
          2850 => x"80",
          2851 => x"87",
          2852 => x"08",
          2853 => x"38",
          2854 => x"8c",
          2855 => x"96",
          2856 => x"0c",
          2857 => x"8c",
          2858 => x"08",
          2859 => x"51",
          2860 => x"38",
          2861 => x"56",
          2862 => x"80",
          2863 => x"85",
          2864 => x"77",
          2865 => x"83",
          2866 => x"75",
          2867 => x"f8",
          2868 => x"3d",
          2869 => x"3d",
          2870 => x"11",
          2871 => x"71",
          2872 => x"81",
          2873 => x"53",
          2874 => x"0d",
          2875 => x"0d",
          2876 => x"33",
          2877 => x"71",
          2878 => x"88",
          2879 => x"14",
          2880 => x"07",
          2881 => x"33",
          2882 => x"f8",
          2883 => x"53",
          2884 => x"52",
          2885 => x"04",
          2886 => x"73",
          2887 => x"92",
          2888 => x"52",
          2889 => x"81",
          2890 => x"70",
          2891 => x"70",
          2892 => x"3d",
          2893 => x"3d",
          2894 => x"52",
          2895 => x"70",
          2896 => x"34",
          2897 => x"51",
          2898 => x"81",
          2899 => x"70",
          2900 => x"70",
          2901 => x"05",
          2902 => x"88",
          2903 => x"72",
          2904 => x"0d",
          2905 => x"0d",
          2906 => x"54",
          2907 => x"80",
          2908 => x"71",
          2909 => x"53",
          2910 => x"81",
          2911 => x"ff",
          2912 => x"39",
          2913 => x"04",
          2914 => x"75",
          2915 => x"52",
          2916 => x"70",
          2917 => x"34",
          2918 => x"70",
          2919 => x"3d",
          2920 => x"3d",
          2921 => x"79",
          2922 => x"74",
          2923 => x"56",
          2924 => x"81",
          2925 => x"71",
          2926 => x"16",
          2927 => x"52",
          2928 => x"86",
          2929 => x"2e",
          2930 => x"81",
          2931 => x"86",
          2932 => x"fe",
          2933 => x"76",
          2934 => x"39",
          2935 => x"8a",
          2936 => x"51",
          2937 => x"71",
          2938 => x"33",
          2939 => x"0c",
          2940 => x"04",
          2941 => x"f8",
          2942 => x"80",
          2943 => x"c8",
          2944 => x"3d",
          2945 => x"80",
          2946 => x"33",
          2947 => x"7a",
          2948 => x"38",
          2949 => x"16",
          2950 => x"16",
          2951 => x"17",
          2952 => x"fa",
          2953 => x"f8",
          2954 => x"2e",
          2955 => x"b7",
          2956 => x"c8",
          2957 => x"34",
          2958 => x"70",
          2959 => x"31",
          2960 => x"59",
          2961 => x"77",
          2962 => x"82",
          2963 => x"74",
          2964 => x"81",
          2965 => x"81",
          2966 => x"53",
          2967 => x"16",
          2968 => x"e3",
          2969 => x"81",
          2970 => x"f8",
          2971 => x"3d",
          2972 => x"3d",
          2973 => x"56",
          2974 => x"74",
          2975 => x"2e",
          2976 => x"51",
          2977 => x"81",
          2978 => x"57",
          2979 => x"08",
          2980 => x"54",
          2981 => x"16",
          2982 => x"33",
          2983 => x"3f",
          2984 => x"08",
          2985 => x"38",
          2986 => x"57",
          2987 => x"0c",
          2988 => x"c8",
          2989 => x"0d",
          2990 => x"0d",
          2991 => x"57",
          2992 => x"81",
          2993 => x"58",
          2994 => x"08",
          2995 => x"76",
          2996 => x"83",
          2997 => x"06",
          2998 => x"84",
          2999 => x"78",
          3000 => x"81",
          3001 => x"38",
          3002 => x"81",
          3003 => x"52",
          3004 => x"52",
          3005 => x"3f",
          3006 => x"52",
          3007 => x"51",
          3008 => x"84",
          3009 => x"d2",
          3010 => x"fc",
          3011 => x"8a",
          3012 => x"52",
          3013 => x"51",
          3014 => x"90",
          3015 => x"84",
          3016 => x"fc",
          3017 => x"17",
          3018 => x"a0",
          3019 => x"86",
          3020 => x"08",
          3021 => x"b0",
          3022 => x"55",
          3023 => x"81",
          3024 => x"f8",
          3025 => x"84",
          3026 => x"53",
          3027 => x"17",
          3028 => x"d7",
          3029 => x"c8",
          3030 => x"83",
          3031 => x"77",
          3032 => x"0c",
          3033 => x"04",
          3034 => x"77",
          3035 => x"12",
          3036 => x"55",
          3037 => x"56",
          3038 => x"8d",
          3039 => x"22",
          3040 => x"ac",
          3041 => x"57",
          3042 => x"f8",
          3043 => x"3d",
          3044 => x"3d",
          3045 => x"70",
          3046 => x"57",
          3047 => x"81",
          3048 => x"98",
          3049 => x"81",
          3050 => x"74",
          3051 => x"72",
          3052 => x"f5",
          3053 => x"24",
          3054 => x"81",
          3055 => x"81",
          3056 => x"83",
          3057 => x"38",
          3058 => x"76",
          3059 => x"70",
          3060 => x"16",
          3061 => x"74",
          3062 => x"96",
          3063 => x"c8",
          3064 => x"38",
          3065 => x"06",
          3066 => x"33",
          3067 => x"89",
          3068 => x"08",
          3069 => x"54",
          3070 => x"fc",
          3071 => x"f8",
          3072 => x"fe",
          3073 => x"ff",
          3074 => x"11",
          3075 => x"2b",
          3076 => x"81",
          3077 => x"2a",
          3078 => x"51",
          3079 => x"e2",
          3080 => x"ff",
          3081 => x"da",
          3082 => x"2a",
          3083 => x"05",
          3084 => x"fc",
          3085 => x"f8",
          3086 => x"c6",
          3087 => x"83",
          3088 => x"05",
          3089 => x"f9",
          3090 => x"f8",
          3091 => x"ff",
          3092 => x"ae",
          3093 => x"2a",
          3094 => x"05",
          3095 => x"fc",
          3096 => x"f8",
          3097 => x"38",
          3098 => x"83",
          3099 => x"05",
          3100 => x"f8",
          3101 => x"f8",
          3102 => x"0a",
          3103 => x"39",
          3104 => x"81",
          3105 => x"89",
          3106 => x"f8",
          3107 => x"7c",
          3108 => x"56",
          3109 => x"77",
          3110 => x"38",
          3111 => x"08",
          3112 => x"38",
          3113 => x"72",
          3114 => x"9d",
          3115 => x"24",
          3116 => x"81",
          3117 => x"82",
          3118 => x"83",
          3119 => x"38",
          3120 => x"76",
          3121 => x"70",
          3122 => x"18",
          3123 => x"76",
          3124 => x"9e",
          3125 => x"c8",
          3126 => x"f8",
          3127 => x"d9",
          3128 => x"ff",
          3129 => x"05",
          3130 => x"81",
          3131 => x"54",
          3132 => x"80",
          3133 => x"77",
          3134 => x"f0",
          3135 => x"8f",
          3136 => x"51",
          3137 => x"34",
          3138 => x"17",
          3139 => x"2a",
          3140 => x"05",
          3141 => x"fa",
          3142 => x"f8",
          3143 => x"81",
          3144 => x"81",
          3145 => x"83",
          3146 => x"b4",
          3147 => x"2a",
          3148 => x"8f",
          3149 => x"2a",
          3150 => x"f0",
          3151 => x"06",
          3152 => x"72",
          3153 => x"ec",
          3154 => x"2a",
          3155 => x"05",
          3156 => x"fa",
          3157 => x"f8",
          3158 => x"81",
          3159 => x"80",
          3160 => x"83",
          3161 => x"52",
          3162 => x"fe",
          3163 => x"b4",
          3164 => x"a4",
          3165 => x"76",
          3166 => x"17",
          3167 => x"75",
          3168 => x"3f",
          3169 => x"08",
          3170 => x"c8",
          3171 => x"77",
          3172 => x"77",
          3173 => x"fc",
          3174 => x"b4",
          3175 => x"51",
          3176 => x"c9",
          3177 => x"c8",
          3178 => x"06",
          3179 => x"72",
          3180 => x"3f",
          3181 => x"17",
          3182 => x"f8",
          3183 => x"3d",
          3184 => x"3d",
          3185 => x"7e",
          3186 => x"56",
          3187 => x"75",
          3188 => x"74",
          3189 => x"27",
          3190 => x"80",
          3191 => x"ff",
          3192 => x"75",
          3193 => x"3f",
          3194 => x"08",
          3195 => x"c8",
          3196 => x"38",
          3197 => x"54",
          3198 => x"81",
          3199 => x"39",
          3200 => x"08",
          3201 => x"39",
          3202 => x"51",
          3203 => x"81",
          3204 => x"58",
          3205 => x"08",
          3206 => x"c7",
          3207 => x"c8",
          3208 => x"d2",
          3209 => x"c8",
          3210 => x"cf",
          3211 => x"74",
          3212 => x"fc",
          3213 => x"f8",
          3214 => x"38",
          3215 => x"fe",
          3216 => x"08",
          3217 => x"74",
          3218 => x"38",
          3219 => x"17",
          3220 => x"33",
          3221 => x"73",
          3222 => x"77",
          3223 => x"26",
          3224 => x"80",
          3225 => x"f8",
          3226 => x"3d",
          3227 => x"3d",
          3228 => x"71",
          3229 => x"5b",
          3230 => x"8c",
          3231 => x"77",
          3232 => x"38",
          3233 => x"78",
          3234 => x"81",
          3235 => x"79",
          3236 => x"f9",
          3237 => x"55",
          3238 => x"c8",
          3239 => x"e0",
          3240 => x"c8",
          3241 => x"f8",
          3242 => x"2e",
          3243 => x"98",
          3244 => x"f8",
          3245 => x"82",
          3246 => x"58",
          3247 => x"70",
          3248 => x"80",
          3249 => x"38",
          3250 => x"09",
          3251 => x"e2",
          3252 => x"56",
          3253 => x"76",
          3254 => x"82",
          3255 => x"7a",
          3256 => x"3f",
          3257 => x"f8",
          3258 => x"2e",
          3259 => x"86",
          3260 => x"c8",
          3261 => x"f8",
          3262 => x"70",
          3263 => x"07",
          3264 => x"7c",
          3265 => x"c8",
          3266 => x"51",
          3267 => x"81",
          3268 => x"f8",
          3269 => x"2e",
          3270 => x"17",
          3271 => x"74",
          3272 => x"73",
          3273 => x"27",
          3274 => x"58",
          3275 => x"80",
          3276 => x"56",
          3277 => x"98",
          3278 => x"26",
          3279 => x"56",
          3280 => x"81",
          3281 => x"52",
          3282 => x"c6",
          3283 => x"c8",
          3284 => x"b8",
          3285 => x"81",
          3286 => x"81",
          3287 => x"06",
          3288 => x"f8",
          3289 => x"81",
          3290 => x"09",
          3291 => x"72",
          3292 => x"70",
          3293 => x"51",
          3294 => x"80",
          3295 => x"78",
          3296 => x"06",
          3297 => x"73",
          3298 => x"39",
          3299 => x"52",
          3300 => x"f7",
          3301 => x"c8",
          3302 => x"c8",
          3303 => x"81",
          3304 => x"07",
          3305 => x"55",
          3306 => x"2e",
          3307 => x"80",
          3308 => x"75",
          3309 => x"76",
          3310 => x"3f",
          3311 => x"08",
          3312 => x"38",
          3313 => x"0c",
          3314 => x"fe",
          3315 => x"08",
          3316 => x"74",
          3317 => x"ff",
          3318 => x"0c",
          3319 => x"81",
          3320 => x"84",
          3321 => x"39",
          3322 => x"81",
          3323 => x"8c",
          3324 => x"8c",
          3325 => x"c8",
          3326 => x"39",
          3327 => x"55",
          3328 => x"c8",
          3329 => x"0d",
          3330 => x"0d",
          3331 => x"55",
          3332 => x"81",
          3333 => x"58",
          3334 => x"f8",
          3335 => x"d8",
          3336 => x"74",
          3337 => x"3f",
          3338 => x"08",
          3339 => x"08",
          3340 => x"59",
          3341 => x"77",
          3342 => x"70",
          3343 => x"c8",
          3344 => x"84",
          3345 => x"56",
          3346 => x"58",
          3347 => x"97",
          3348 => x"75",
          3349 => x"52",
          3350 => x"51",
          3351 => x"81",
          3352 => x"80",
          3353 => x"8a",
          3354 => x"32",
          3355 => x"72",
          3356 => x"2a",
          3357 => x"56",
          3358 => x"c8",
          3359 => x"0d",
          3360 => x"0d",
          3361 => x"08",
          3362 => x"74",
          3363 => x"26",
          3364 => x"74",
          3365 => x"72",
          3366 => x"74",
          3367 => x"88",
          3368 => x"73",
          3369 => x"33",
          3370 => x"27",
          3371 => x"16",
          3372 => x"9b",
          3373 => x"2a",
          3374 => x"88",
          3375 => x"58",
          3376 => x"80",
          3377 => x"16",
          3378 => x"0c",
          3379 => x"8a",
          3380 => x"89",
          3381 => x"72",
          3382 => x"38",
          3383 => x"51",
          3384 => x"81",
          3385 => x"54",
          3386 => x"08",
          3387 => x"38",
          3388 => x"f8",
          3389 => x"8b",
          3390 => x"08",
          3391 => x"08",
          3392 => x"82",
          3393 => x"74",
          3394 => x"cb",
          3395 => x"75",
          3396 => x"3f",
          3397 => x"08",
          3398 => x"73",
          3399 => x"98",
          3400 => x"82",
          3401 => x"2e",
          3402 => x"39",
          3403 => x"39",
          3404 => x"13",
          3405 => x"74",
          3406 => x"16",
          3407 => x"18",
          3408 => x"77",
          3409 => x"0c",
          3410 => x"04",
          3411 => x"7a",
          3412 => x"12",
          3413 => x"59",
          3414 => x"80",
          3415 => x"86",
          3416 => x"98",
          3417 => x"14",
          3418 => x"55",
          3419 => x"81",
          3420 => x"83",
          3421 => x"77",
          3422 => x"81",
          3423 => x"0c",
          3424 => x"55",
          3425 => x"76",
          3426 => x"17",
          3427 => x"74",
          3428 => x"9b",
          3429 => x"39",
          3430 => x"ff",
          3431 => x"2a",
          3432 => x"81",
          3433 => x"52",
          3434 => x"e6",
          3435 => x"c8",
          3436 => x"55",
          3437 => x"f8",
          3438 => x"80",
          3439 => x"55",
          3440 => x"08",
          3441 => x"f4",
          3442 => x"08",
          3443 => x"08",
          3444 => x"38",
          3445 => x"77",
          3446 => x"84",
          3447 => x"39",
          3448 => x"52",
          3449 => x"86",
          3450 => x"c8",
          3451 => x"55",
          3452 => x"08",
          3453 => x"c4",
          3454 => x"81",
          3455 => x"81",
          3456 => x"81",
          3457 => x"c8",
          3458 => x"b0",
          3459 => x"c8",
          3460 => x"51",
          3461 => x"81",
          3462 => x"a0",
          3463 => x"15",
          3464 => x"75",
          3465 => x"3f",
          3466 => x"08",
          3467 => x"76",
          3468 => x"77",
          3469 => x"9c",
          3470 => x"55",
          3471 => x"c8",
          3472 => x"0d",
          3473 => x"0d",
          3474 => x"08",
          3475 => x"80",
          3476 => x"fc",
          3477 => x"f8",
          3478 => x"81",
          3479 => x"80",
          3480 => x"f8",
          3481 => x"98",
          3482 => x"78",
          3483 => x"3f",
          3484 => x"08",
          3485 => x"c8",
          3486 => x"38",
          3487 => x"08",
          3488 => x"70",
          3489 => x"58",
          3490 => x"2e",
          3491 => x"83",
          3492 => x"81",
          3493 => x"55",
          3494 => x"81",
          3495 => x"07",
          3496 => x"2e",
          3497 => x"16",
          3498 => x"2e",
          3499 => x"88",
          3500 => x"81",
          3501 => x"56",
          3502 => x"51",
          3503 => x"81",
          3504 => x"54",
          3505 => x"08",
          3506 => x"9b",
          3507 => x"2e",
          3508 => x"83",
          3509 => x"73",
          3510 => x"0c",
          3511 => x"04",
          3512 => x"76",
          3513 => x"54",
          3514 => x"81",
          3515 => x"83",
          3516 => x"76",
          3517 => x"53",
          3518 => x"2e",
          3519 => x"90",
          3520 => x"51",
          3521 => x"81",
          3522 => x"90",
          3523 => x"53",
          3524 => x"c8",
          3525 => x"0d",
          3526 => x"0d",
          3527 => x"83",
          3528 => x"54",
          3529 => x"55",
          3530 => x"3f",
          3531 => x"51",
          3532 => x"2e",
          3533 => x"8b",
          3534 => x"2a",
          3535 => x"51",
          3536 => x"86",
          3537 => x"f7",
          3538 => x"7d",
          3539 => x"75",
          3540 => x"98",
          3541 => x"2e",
          3542 => x"98",
          3543 => x"78",
          3544 => x"3f",
          3545 => x"08",
          3546 => x"c8",
          3547 => x"38",
          3548 => x"70",
          3549 => x"73",
          3550 => x"58",
          3551 => x"8b",
          3552 => x"bf",
          3553 => x"ff",
          3554 => x"53",
          3555 => x"34",
          3556 => x"08",
          3557 => x"e5",
          3558 => x"81",
          3559 => x"2e",
          3560 => x"70",
          3561 => x"57",
          3562 => x"9e",
          3563 => x"2e",
          3564 => x"f8",
          3565 => x"df",
          3566 => x"72",
          3567 => x"81",
          3568 => x"76",
          3569 => x"2e",
          3570 => x"52",
          3571 => x"fc",
          3572 => x"c8",
          3573 => x"f8",
          3574 => x"38",
          3575 => x"fe",
          3576 => x"39",
          3577 => x"16",
          3578 => x"f8",
          3579 => x"3d",
          3580 => x"3d",
          3581 => x"08",
          3582 => x"52",
          3583 => x"c5",
          3584 => x"c8",
          3585 => x"f8",
          3586 => x"38",
          3587 => x"52",
          3588 => x"de",
          3589 => x"c8",
          3590 => x"f8",
          3591 => x"38",
          3592 => x"f8",
          3593 => x"9c",
          3594 => x"ea",
          3595 => x"53",
          3596 => x"9c",
          3597 => x"ea",
          3598 => x"0b",
          3599 => x"74",
          3600 => x"0c",
          3601 => x"04",
          3602 => x"75",
          3603 => x"12",
          3604 => x"53",
          3605 => x"9a",
          3606 => x"c8",
          3607 => x"9c",
          3608 => x"e5",
          3609 => x"0b",
          3610 => x"85",
          3611 => x"fa",
          3612 => x"7a",
          3613 => x"0b",
          3614 => x"98",
          3615 => x"2e",
          3616 => x"80",
          3617 => x"55",
          3618 => x"17",
          3619 => x"33",
          3620 => x"51",
          3621 => x"2e",
          3622 => x"85",
          3623 => x"06",
          3624 => x"e5",
          3625 => x"2e",
          3626 => x"8b",
          3627 => x"70",
          3628 => x"34",
          3629 => x"71",
          3630 => x"05",
          3631 => x"15",
          3632 => x"27",
          3633 => x"15",
          3634 => x"80",
          3635 => x"34",
          3636 => x"52",
          3637 => x"88",
          3638 => x"17",
          3639 => x"52",
          3640 => x"3f",
          3641 => x"08",
          3642 => x"12",
          3643 => x"3f",
          3644 => x"08",
          3645 => x"98",
          3646 => x"da",
          3647 => x"c8",
          3648 => x"23",
          3649 => x"04",
          3650 => x"7f",
          3651 => x"5b",
          3652 => x"33",
          3653 => x"73",
          3654 => x"38",
          3655 => x"80",
          3656 => x"38",
          3657 => x"8c",
          3658 => x"08",
          3659 => x"aa",
          3660 => x"41",
          3661 => x"33",
          3662 => x"73",
          3663 => x"81",
          3664 => x"81",
          3665 => x"dc",
          3666 => x"70",
          3667 => x"07",
          3668 => x"73",
          3669 => x"88",
          3670 => x"70",
          3671 => x"73",
          3672 => x"38",
          3673 => x"ab",
          3674 => x"52",
          3675 => x"91",
          3676 => x"c8",
          3677 => x"98",
          3678 => x"61",
          3679 => x"5a",
          3680 => x"a0",
          3681 => x"e7",
          3682 => x"70",
          3683 => x"79",
          3684 => x"73",
          3685 => x"81",
          3686 => x"38",
          3687 => x"33",
          3688 => x"ae",
          3689 => x"70",
          3690 => x"82",
          3691 => x"51",
          3692 => x"54",
          3693 => x"79",
          3694 => x"74",
          3695 => x"57",
          3696 => x"af",
          3697 => x"70",
          3698 => x"51",
          3699 => x"dc",
          3700 => x"73",
          3701 => x"38",
          3702 => x"82",
          3703 => x"19",
          3704 => x"54",
          3705 => x"82",
          3706 => x"54",
          3707 => x"78",
          3708 => x"81",
          3709 => x"54",
          3710 => x"81",
          3711 => x"af",
          3712 => x"77",
          3713 => x"70",
          3714 => x"25",
          3715 => x"07",
          3716 => x"51",
          3717 => x"2e",
          3718 => x"39",
          3719 => x"80",
          3720 => x"33",
          3721 => x"73",
          3722 => x"81",
          3723 => x"81",
          3724 => x"dc",
          3725 => x"70",
          3726 => x"07",
          3727 => x"73",
          3728 => x"b5",
          3729 => x"2e",
          3730 => x"83",
          3731 => x"76",
          3732 => x"07",
          3733 => x"2e",
          3734 => x"8b",
          3735 => x"77",
          3736 => x"30",
          3737 => x"71",
          3738 => x"53",
          3739 => x"55",
          3740 => x"38",
          3741 => x"5c",
          3742 => x"75",
          3743 => x"73",
          3744 => x"38",
          3745 => x"06",
          3746 => x"11",
          3747 => x"75",
          3748 => x"3f",
          3749 => x"08",
          3750 => x"38",
          3751 => x"33",
          3752 => x"54",
          3753 => x"e6",
          3754 => x"f8",
          3755 => x"2e",
          3756 => x"ff",
          3757 => x"74",
          3758 => x"38",
          3759 => x"75",
          3760 => x"17",
          3761 => x"57",
          3762 => x"a7",
          3763 => x"81",
          3764 => x"e5",
          3765 => x"f8",
          3766 => x"38",
          3767 => x"54",
          3768 => x"89",
          3769 => x"70",
          3770 => x"57",
          3771 => x"54",
          3772 => x"81",
          3773 => x"f7",
          3774 => x"7e",
          3775 => x"2e",
          3776 => x"33",
          3777 => x"e5",
          3778 => x"06",
          3779 => x"7a",
          3780 => x"a0",
          3781 => x"38",
          3782 => x"55",
          3783 => x"84",
          3784 => x"39",
          3785 => x"8b",
          3786 => x"7b",
          3787 => x"7a",
          3788 => x"3f",
          3789 => x"08",
          3790 => x"c8",
          3791 => x"38",
          3792 => x"52",
          3793 => x"aa",
          3794 => x"c8",
          3795 => x"f8",
          3796 => x"c2",
          3797 => x"08",
          3798 => x"55",
          3799 => x"ff",
          3800 => x"15",
          3801 => x"54",
          3802 => x"34",
          3803 => x"70",
          3804 => x"81",
          3805 => x"58",
          3806 => x"8b",
          3807 => x"74",
          3808 => x"3f",
          3809 => x"08",
          3810 => x"38",
          3811 => x"51",
          3812 => x"ff",
          3813 => x"ab",
          3814 => x"55",
          3815 => x"bb",
          3816 => x"2e",
          3817 => x"80",
          3818 => x"85",
          3819 => x"06",
          3820 => x"58",
          3821 => x"80",
          3822 => x"75",
          3823 => x"73",
          3824 => x"b5",
          3825 => x"0b",
          3826 => x"80",
          3827 => x"39",
          3828 => x"54",
          3829 => x"85",
          3830 => x"75",
          3831 => x"81",
          3832 => x"73",
          3833 => x"1b",
          3834 => x"2a",
          3835 => x"51",
          3836 => x"80",
          3837 => x"90",
          3838 => x"ff",
          3839 => x"05",
          3840 => x"f5",
          3841 => x"f8",
          3842 => x"1c",
          3843 => x"39",
          3844 => x"c8",
          3845 => x"0d",
          3846 => x"0d",
          3847 => x"7b",
          3848 => x"73",
          3849 => x"55",
          3850 => x"2e",
          3851 => x"75",
          3852 => x"57",
          3853 => x"26",
          3854 => x"ba",
          3855 => x"70",
          3856 => x"ba",
          3857 => x"06",
          3858 => x"73",
          3859 => x"70",
          3860 => x"51",
          3861 => x"89",
          3862 => x"82",
          3863 => x"ff",
          3864 => x"56",
          3865 => x"2e",
          3866 => x"80",
          3867 => x"c8",
          3868 => x"08",
          3869 => x"76",
          3870 => x"58",
          3871 => x"81",
          3872 => x"ff",
          3873 => x"53",
          3874 => x"26",
          3875 => x"13",
          3876 => x"06",
          3877 => x"9f",
          3878 => x"99",
          3879 => x"e0",
          3880 => x"ff",
          3881 => x"72",
          3882 => x"2a",
          3883 => x"72",
          3884 => x"06",
          3885 => x"ff",
          3886 => x"30",
          3887 => x"70",
          3888 => x"07",
          3889 => x"9f",
          3890 => x"54",
          3891 => x"80",
          3892 => x"81",
          3893 => x"59",
          3894 => x"25",
          3895 => x"8b",
          3896 => x"24",
          3897 => x"76",
          3898 => x"78",
          3899 => x"81",
          3900 => x"51",
          3901 => x"c8",
          3902 => x"0d",
          3903 => x"0d",
          3904 => x"0b",
          3905 => x"ff",
          3906 => x"0c",
          3907 => x"51",
          3908 => x"84",
          3909 => x"c8",
          3910 => x"38",
          3911 => x"51",
          3912 => x"81",
          3913 => x"83",
          3914 => x"54",
          3915 => x"82",
          3916 => x"09",
          3917 => x"e3",
          3918 => x"b4",
          3919 => x"57",
          3920 => x"2e",
          3921 => x"83",
          3922 => x"74",
          3923 => x"70",
          3924 => x"25",
          3925 => x"51",
          3926 => x"38",
          3927 => x"2e",
          3928 => x"b5",
          3929 => x"81",
          3930 => x"80",
          3931 => x"e0",
          3932 => x"f8",
          3933 => x"81",
          3934 => x"80",
          3935 => x"85",
          3936 => x"8c",
          3937 => x"16",
          3938 => x"3f",
          3939 => x"08",
          3940 => x"c8",
          3941 => x"83",
          3942 => x"74",
          3943 => x"0c",
          3944 => x"04",
          3945 => x"61",
          3946 => x"80",
          3947 => x"58",
          3948 => x"0c",
          3949 => x"e1",
          3950 => x"c8",
          3951 => x"56",
          3952 => x"f8",
          3953 => x"86",
          3954 => x"f8",
          3955 => x"29",
          3956 => x"05",
          3957 => x"53",
          3958 => x"80",
          3959 => x"38",
          3960 => x"76",
          3961 => x"74",
          3962 => x"72",
          3963 => x"38",
          3964 => x"51",
          3965 => x"81",
          3966 => x"81",
          3967 => x"81",
          3968 => x"72",
          3969 => x"80",
          3970 => x"38",
          3971 => x"70",
          3972 => x"53",
          3973 => x"86",
          3974 => x"a7",
          3975 => x"34",
          3976 => x"34",
          3977 => x"14",
          3978 => x"b2",
          3979 => x"c8",
          3980 => x"06",
          3981 => x"54",
          3982 => x"72",
          3983 => x"76",
          3984 => x"38",
          3985 => x"70",
          3986 => x"53",
          3987 => x"85",
          3988 => x"70",
          3989 => x"5b",
          3990 => x"81",
          3991 => x"81",
          3992 => x"76",
          3993 => x"81",
          3994 => x"38",
          3995 => x"56",
          3996 => x"83",
          3997 => x"70",
          3998 => x"80",
          3999 => x"83",
          4000 => x"dc",
          4001 => x"f8",
          4002 => x"76",
          4003 => x"05",
          4004 => x"16",
          4005 => x"56",
          4006 => x"d7",
          4007 => x"8d",
          4008 => x"72",
          4009 => x"54",
          4010 => x"57",
          4011 => x"95",
          4012 => x"73",
          4013 => x"3f",
          4014 => x"08",
          4015 => x"57",
          4016 => x"89",
          4017 => x"56",
          4018 => x"d7",
          4019 => x"76",
          4020 => x"f1",
          4021 => x"76",
          4022 => x"e9",
          4023 => x"51",
          4024 => x"81",
          4025 => x"83",
          4026 => x"53",
          4027 => x"2e",
          4028 => x"84",
          4029 => x"ca",
          4030 => x"da",
          4031 => x"c8",
          4032 => x"ff",
          4033 => x"8d",
          4034 => x"14",
          4035 => x"3f",
          4036 => x"08",
          4037 => x"15",
          4038 => x"14",
          4039 => x"34",
          4040 => x"33",
          4041 => x"81",
          4042 => x"54",
          4043 => x"72",
          4044 => x"91",
          4045 => x"ff",
          4046 => x"29",
          4047 => x"33",
          4048 => x"72",
          4049 => x"72",
          4050 => x"38",
          4051 => x"06",
          4052 => x"2e",
          4053 => x"56",
          4054 => x"80",
          4055 => x"da",
          4056 => x"f8",
          4057 => x"81",
          4058 => x"88",
          4059 => x"8f",
          4060 => x"56",
          4061 => x"38",
          4062 => x"51",
          4063 => x"81",
          4064 => x"83",
          4065 => x"55",
          4066 => x"80",
          4067 => x"da",
          4068 => x"f8",
          4069 => x"80",
          4070 => x"da",
          4071 => x"f8",
          4072 => x"ff",
          4073 => x"8d",
          4074 => x"2e",
          4075 => x"88",
          4076 => x"14",
          4077 => x"05",
          4078 => x"75",
          4079 => x"38",
          4080 => x"52",
          4081 => x"51",
          4082 => x"3f",
          4083 => x"08",
          4084 => x"c8",
          4085 => x"82",
          4086 => x"f8",
          4087 => x"ff",
          4088 => x"26",
          4089 => x"57",
          4090 => x"f5",
          4091 => x"82",
          4092 => x"f5",
          4093 => x"81",
          4094 => x"8d",
          4095 => x"2e",
          4096 => x"82",
          4097 => x"16",
          4098 => x"16",
          4099 => x"70",
          4100 => x"7a",
          4101 => x"0c",
          4102 => x"83",
          4103 => x"06",
          4104 => x"de",
          4105 => x"ae",
          4106 => x"c8",
          4107 => x"ff",
          4108 => x"56",
          4109 => x"38",
          4110 => x"38",
          4111 => x"51",
          4112 => x"81",
          4113 => x"a8",
          4114 => x"82",
          4115 => x"39",
          4116 => x"80",
          4117 => x"38",
          4118 => x"15",
          4119 => x"53",
          4120 => x"8d",
          4121 => x"15",
          4122 => x"76",
          4123 => x"51",
          4124 => x"13",
          4125 => x"8d",
          4126 => x"15",
          4127 => x"c5",
          4128 => x"90",
          4129 => x"0b",
          4130 => x"ff",
          4131 => x"15",
          4132 => x"2e",
          4133 => x"81",
          4134 => x"e4",
          4135 => x"b6",
          4136 => x"c8",
          4137 => x"ff",
          4138 => x"81",
          4139 => x"06",
          4140 => x"81",
          4141 => x"51",
          4142 => x"81",
          4143 => x"80",
          4144 => x"f8",
          4145 => x"15",
          4146 => x"14",
          4147 => x"3f",
          4148 => x"08",
          4149 => x"06",
          4150 => x"d4",
          4151 => x"81",
          4152 => x"38",
          4153 => x"d8",
          4154 => x"f8",
          4155 => x"8b",
          4156 => x"2e",
          4157 => x"b3",
          4158 => x"14",
          4159 => x"3f",
          4160 => x"08",
          4161 => x"e4",
          4162 => x"81",
          4163 => x"84",
          4164 => x"d7",
          4165 => x"f8",
          4166 => x"15",
          4167 => x"14",
          4168 => x"3f",
          4169 => x"08",
          4170 => x"76",
          4171 => x"f9",
          4172 => x"05",
          4173 => x"f9",
          4174 => x"86",
          4175 => x"0b",
          4176 => x"80",
          4177 => x"f8",
          4178 => x"3d",
          4179 => x"3d",
          4180 => x"89",
          4181 => x"2e",
          4182 => x"08",
          4183 => x"2e",
          4184 => x"33",
          4185 => x"2e",
          4186 => x"13",
          4187 => x"22",
          4188 => x"76",
          4189 => x"06",
          4190 => x"13",
          4191 => x"c0",
          4192 => x"c8",
          4193 => x"52",
          4194 => x"71",
          4195 => x"55",
          4196 => x"53",
          4197 => x"0c",
          4198 => x"f8",
          4199 => x"3d",
          4200 => x"3d",
          4201 => x"05",
          4202 => x"89",
          4203 => x"52",
          4204 => x"3f",
          4205 => x"0b",
          4206 => x"08",
          4207 => x"81",
          4208 => x"84",
          4209 => x"f8",
          4210 => x"55",
          4211 => x"2e",
          4212 => x"74",
          4213 => x"73",
          4214 => x"38",
          4215 => x"78",
          4216 => x"54",
          4217 => x"92",
          4218 => x"89",
          4219 => x"84",
          4220 => x"b0",
          4221 => x"c8",
          4222 => x"81",
          4223 => x"88",
          4224 => x"eb",
          4225 => x"02",
          4226 => x"e7",
          4227 => x"59",
          4228 => x"80",
          4229 => x"38",
          4230 => x"70",
          4231 => x"d0",
          4232 => x"3d",
          4233 => x"58",
          4234 => x"81",
          4235 => x"55",
          4236 => x"08",
          4237 => x"7a",
          4238 => x"8c",
          4239 => x"56",
          4240 => x"81",
          4241 => x"55",
          4242 => x"08",
          4243 => x"80",
          4244 => x"70",
          4245 => x"57",
          4246 => x"83",
          4247 => x"77",
          4248 => x"73",
          4249 => x"ab",
          4250 => x"2e",
          4251 => x"84",
          4252 => x"06",
          4253 => x"51",
          4254 => x"81",
          4255 => x"55",
          4256 => x"b2",
          4257 => x"06",
          4258 => x"b8",
          4259 => x"2a",
          4260 => x"51",
          4261 => x"2e",
          4262 => x"55",
          4263 => x"77",
          4264 => x"74",
          4265 => x"77",
          4266 => x"81",
          4267 => x"73",
          4268 => x"af",
          4269 => x"7a",
          4270 => x"3f",
          4271 => x"08",
          4272 => x"b2",
          4273 => x"8e",
          4274 => x"ea",
          4275 => x"a0",
          4276 => x"34",
          4277 => x"52",
          4278 => x"bd",
          4279 => x"62",
          4280 => x"d4",
          4281 => x"54",
          4282 => x"15",
          4283 => x"2e",
          4284 => x"7a",
          4285 => x"51",
          4286 => x"75",
          4287 => x"d4",
          4288 => x"be",
          4289 => x"c8",
          4290 => x"f8",
          4291 => x"ca",
          4292 => x"74",
          4293 => x"02",
          4294 => x"70",
          4295 => x"81",
          4296 => x"56",
          4297 => x"86",
          4298 => x"82",
          4299 => x"81",
          4300 => x"06",
          4301 => x"80",
          4302 => x"75",
          4303 => x"73",
          4304 => x"38",
          4305 => x"92",
          4306 => x"7a",
          4307 => x"3f",
          4308 => x"08",
          4309 => x"8c",
          4310 => x"55",
          4311 => x"08",
          4312 => x"77",
          4313 => x"81",
          4314 => x"73",
          4315 => x"38",
          4316 => x"07",
          4317 => x"11",
          4318 => x"0c",
          4319 => x"0c",
          4320 => x"52",
          4321 => x"3f",
          4322 => x"08",
          4323 => x"08",
          4324 => x"63",
          4325 => x"5a",
          4326 => x"81",
          4327 => x"81",
          4328 => x"8c",
          4329 => x"7a",
          4330 => x"17",
          4331 => x"23",
          4332 => x"34",
          4333 => x"1a",
          4334 => x"9c",
          4335 => x"0b",
          4336 => x"77",
          4337 => x"81",
          4338 => x"73",
          4339 => x"8d",
          4340 => x"c8",
          4341 => x"81",
          4342 => x"f8",
          4343 => x"1a",
          4344 => x"22",
          4345 => x"7b",
          4346 => x"a8",
          4347 => x"78",
          4348 => x"3f",
          4349 => x"08",
          4350 => x"c8",
          4351 => x"83",
          4352 => x"81",
          4353 => x"ff",
          4354 => x"06",
          4355 => x"55",
          4356 => x"56",
          4357 => x"76",
          4358 => x"51",
          4359 => x"27",
          4360 => x"70",
          4361 => x"5a",
          4362 => x"76",
          4363 => x"74",
          4364 => x"83",
          4365 => x"73",
          4366 => x"38",
          4367 => x"51",
          4368 => x"81",
          4369 => x"85",
          4370 => x"8e",
          4371 => x"2a",
          4372 => x"08",
          4373 => x"0c",
          4374 => x"79",
          4375 => x"73",
          4376 => x"0c",
          4377 => x"04",
          4378 => x"60",
          4379 => x"40",
          4380 => x"80",
          4381 => x"3d",
          4382 => x"78",
          4383 => x"3f",
          4384 => x"08",
          4385 => x"c8",
          4386 => x"91",
          4387 => x"74",
          4388 => x"38",
          4389 => x"c4",
          4390 => x"33",
          4391 => x"87",
          4392 => x"2e",
          4393 => x"95",
          4394 => x"91",
          4395 => x"56",
          4396 => x"81",
          4397 => x"34",
          4398 => x"a0",
          4399 => x"08",
          4400 => x"31",
          4401 => x"27",
          4402 => x"5c",
          4403 => x"82",
          4404 => x"19",
          4405 => x"ff",
          4406 => x"74",
          4407 => x"7e",
          4408 => x"ff",
          4409 => x"2a",
          4410 => x"79",
          4411 => x"87",
          4412 => x"08",
          4413 => x"98",
          4414 => x"78",
          4415 => x"3f",
          4416 => x"08",
          4417 => x"27",
          4418 => x"74",
          4419 => x"a3",
          4420 => x"1a",
          4421 => x"08",
          4422 => x"d4",
          4423 => x"f8",
          4424 => x"2e",
          4425 => x"81",
          4426 => x"1a",
          4427 => x"59",
          4428 => x"2e",
          4429 => x"77",
          4430 => x"11",
          4431 => x"55",
          4432 => x"85",
          4433 => x"31",
          4434 => x"76",
          4435 => x"81",
          4436 => x"ca",
          4437 => x"f8",
          4438 => x"d7",
          4439 => x"11",
          4440 => x"74",
          4441 => x"38",
          4442 => x"77",
          4443 => x"78",
          4444 => x"84",
          4445 => x"16",
          4446 => x"08",
          4447 => x"2b",
          4448 => x"cf",
          4449 => x"89",
          4450 => x"39",
          4451 => x"0c",
          4452 => x"83",
          4453 => x"80",
          4454 => x"55",
          4455 => x"83",
          4456 => x"9c",
          4457 => x"7e",
          4458 => x"3f",
          4459 => x"08",
          4460 => x"75",
          4461 => x"08",
          4462 => x"1f",
          4463 => x"7c",
          4464 => x"3f",
          4465 => x"7e",
          4466 => x"0c",
          4467 => x"1b",
          4468 => x"1c",
          4469 => x"fd",
          4470 => x"56",
          4471 => x"c8",
          4472 => x"0d",
          4473 => x"0d",
          4474 => x"64",
          4475 => x"58",
          4476 => x"90",
          4477 => x"52",
          4478 => x"d2",
          4479 => x"c8",
          4480 => x"f8",
          4481 => x"38",
          4482 => x"55",
          4483 => x"86",
          4484 => x"83",
          4485 => x"18",
          4486 => x"2a",
          4487 => x"51",
          4488 => x"56",
          4489 => x"83",
          4490 => x"39",
          4491 => x"19",
          4492 => x"83",
          4493 => x"0b",
          4494 => x"81",
          4495 => x"39",
          4496 => x"7c",
          4497 => x"74",
          4498 => x"38",
          4499 => x"7b",
          4500 => x"ec",
          4501 => x"08",
          4502 => x"06",
          4503 => x"81",
          4504 => x"8a",
          4505 => x"05",
          4506 => x"06",
          4507 => x"bf",
          4508 => x"38",
          4509 => x"55",
          4510 => x"7a",
          4511 => x"98",
          4512 => x"77",
          4513 => x"3f",
          4514 => x"08",
          4515 => x"c8",
          4516 => x"82",
          4517 => x"81",
          4518 => x"38",
          4519 => x"ff",
          4520 => x"98",
          4521 => x"18",
          4522 => x"74",
          4523 => x"7e",
          4524 => x"08",
          4525 => x"2e",
          4526 => x"8d",
          4527 => x"ce",
          4528 => x"f8",
          4529 => x"ee",
          4530 => x"08",
          4531 => x"d1",
          4532 => x"f8",
          4533 => x"2e",
          4534 => x"81",
          4535 => x"1b",
          4536 => x"5a",
          4537 => x"2e",
          4538 => x"78",
          4539 => x"11",
          4540 => x"55",
          4541 => x"85",
          4542 => x"31",
          4543 => x"76",
          4544 => x"81",
          4545 => x"c8",
          4546 => x"f8",
          4547 => x"a6",
          4548 => x"11",
          4549 => x"56",
          4550 => x"27",
          4551 => x"80",
          4552 => x"08",
          4553 => x"2b",
          4554 => x"b4",
          4555 => x"b5",
          4556 => x"80",
          4557 => x"34",
          4558 => x"56",
          4559 => x"8c",
          4560 => x"19",
          4561 => x"38",
          4562 => x"b6",
          4563 => x"c8",
          4564 => x"38",
          4565 => x"12",
          4566 => x"9c",
          4567 => x"18",
          4568 => x"06",
          4569 => x"31",
          4570 => x"76",
          4571 => x"7b",
          4572 => x"08",
          4573 => x"cd",
          4574 => x"f8",
          4575 => x"b6",
          4576 => x"7c",
          4577 => x"08",
          4578 => x"1f",
          4579 => x"cb",
          4580 => x"55",
          4581 => x"16",
          4582 => x"31",
          4583 => x"7f",
          4584 => x"94",
          4585 => x"70",
          4586 => x"8c",
          4587 => x"58",
          4588 => x"76",
          4589 => x"75",
          4590 => x"19",
          4591 => x"39",
          4592 => x"80",
          4593 => x"74",
          4594 => x"80",
          4595 => x"f8",
          4596 => x"3d",
          4597 => x"3d",
          4598 => x"3d",
          4599 => x"70",
          4600 => x"ea",
          4601 => x"c8",
          4602 => x"f8",
          4603 => x"fb",
          4604 => x"33",
          4605 => x"70",
          4606 => x"55",
          4607 => x"2e",
          4608 => x"a0",
          4609 => x"78",
          4610 => x"3f",
          4611 => x"08",
          4612 => x"c8",
          4613 => x"38",
          4614 => x"8b",
          4615 => x"07",
          4616 => x"8b",
          4617 => x"16",
          4618 => x"52",
          4619 => x"dd",
          4620 => x"16",
          4621 => x"15",
          4622 => x"3f",
          4623 => x"0a",
          4624 => x"51",
          4625 => x"76",
          4626 => x"51",
          4627 => x"78",
          4628 => x"83",
          4629 => x"51",
          4630 => x"81",
          4631 => x"90",
          4632 => x"bf",
          4633 => x"73",
          4634 => x"76",
          4635 => x"0c",
          4636 => x"04",
          4637 => x"76",
          4638 => x"fe",
          4639 => x"f8",
          4640 => x"81",
          4641 => x"9c",
          4642 => x"fc",
          4643 => x"51",
          4644 => x"81",
          4645 => x"53",
          4646 => x"08",
          4647 => x"f8",
          4648 => x"0c",
          4649 => x"c8",
          4650 => x"0d",
          4651 => x"0d",
          4652 => x"e6",
          4653 => x"52",
          4654 => x"f8",
          4655 => x"8b",
          4656 => x"c8",
          4657 => x"8c",
          4658 => x"71",
          4659 => x"0c",
          4660 => x"04",
          4661 => x"80",
          4662 => x"d0",
          4663 => x"3d",
          4664 => x"3f",
          4665 => x"08",
          4666 => x"c8",
          4667 => x"38",
          4668 => x"52",
          4669 => x"05",
          4670 => x"3f",
          4671 => x"08",
          4672 => x"c8",
          4673 => x"02",
          4674 => x"33",
          4675 => x"55",
          4676 => x"25",
          4677 => x"7a",
          4678 => x"54",
          4679 => x"a2",
          4680 => x"84",
          4681 => x"06",
          4682 => x"73",
          4683 => x"38",
          4684 => x"70",
          4685 => x"a8",
          4686 => x"c8",
          4687 => x"0c",
          4688 => x"f8",
          4689 => x"2e",
          4690 => x"83",
          4691 => x"74",
          4692 => x"0c",
          4693 => x"04",
          4694 => x"6f",
          4695 => x"80",
          4696 => x"53",
          4697 => x"b8",
          4698 => x"3d",
          4699 => x"3f",
          4700 => x"08",
          4701 => x"c8",
          4702 => x"38",
          4703 => x"7c",
          4704 => x"47",
          4705 => x"54",
          4706 => x"81",
          4707 => x"52",
          4708 => x"52",
          4709 => x"3f",
          4710 => x"08",
          4711 => x"c8",
          4712 => x"38",
          4713 => x"51",
          4714 => x"81",
          4715 => x"57",
          4716 => x"08",
          4717 => x"69",
          4718 => x"da",
          4719 => x"f8",
          4720 => x"76",
          4721 => x"d5",
          4722 => x"f8",
          4723 => x"81",
          4724 => x"82",
          4725 => x"52",
          4726 => x"eb",
          4727 => x"c8",
          4728 => x"f8",
          4729 => x"38",
          4730 => x"51",
          4731 => x"73",
          4732 => x"08",
          4733 => x"76",
          4734 => x"d6",
          4735 => x"f8",
          4736 => x"81",
          4737 => x"80",
          4738 => x"76",
          4739 => x"81",
          4740 => x"82",
          4741 => x"39",
          4742 => x"38",
          4743 => x"bc",
          4744 => x"51",
          4745 => x"76",
          4746 => x"11",
          4747 => x"51",
          4748 => x"73",
          4749 => x"38",
          4750 => x"55",
          4751 => x"16",
          4752 => x"56",
          4753 => x"38",
          4754 => x"73",
          4755 => x"90",
          4756 => x"2e",
          4757 => x"16",
          4758 => x"ff",
          4759 => x"ff",
          4760 => x"58",
          4761 => x"74",
          4762 => x"75",
          4763 => x"18",
          4764 => x"58",
          4765 => x"fe",
          4766 => x"7b",
          4767 => x"06",
          4768 => x"18",
          4769 => x"58",
          4770 => x"80",
          4771 => x"8c",
          4772 => x"29",
          4773 => x"05",
          4774 => x"33",
          4775 => x"56",
          4776 => x"2e",
          4777 => x"16",
          4778 => x"33",
          4779 => x"73",
          4780 => x"16",
          4781 => x"26",
          4782 => x"55",
          4783 => x"91",
          4784 => x"54",
          4785 => x"70",
          4786 => x"34",
          4787 => x"ec",
          4788 => x"70",
          4789 => x"34",
          4790 => x"09",
          4791 => x"38",
          4792 => x"39",
          4793 => x"19",
          4794 => x"33",
          4795 => x"05",
          4796 => x"78",
          4797 => x"80",
          4798 => x"81",
          4799 => x"9e",
          4800 => x"f7",
          4801 => x"7d",
          4802 => x"05",
          4803 => x"57",
          4804 => x"3f",
          4805 => x"08",
          4806 => x"c8",
          4807 => x"38",
          4808 => x"53",
          4809 => x"38",
          4810 => x"54",
          4811 => x"92",
          4812 => x"33",
          4813 => x"70",
          4814 => x"54",
          4815 => x"38",
          4816 => x"15",
          4817 => x"70",
          4818 => x"58",
          4819 => x"82",
          4820 => x"8a",
          4821 => x"89",
          4822 => x"53",
          4823 => x"b7",
          4824 => x"ff",
          4825 => x"fc",
          4826 => x"f8",
          4827 => x"15",
          4828 => x"53",
          4829 => x"fc",
          4830 => x"f8",
          4831 => x"26",
          4832 => x"30",
          4833 => x"70",
          4834 => x"77",
          4835 => x"18",
          4836 => x"51",
          4837 => x"88",
          4838 => x"73",
          4839 => x"52",
          4840 => x"ca",
          4841 => x"c8",
          4842 => x"f8",
          4843 => x"2e",
          4844 => x"81",
          4845 => x"ff",
          4846 => x"38",
          4847 => x"08",
          4848 => x"73",
          4849 => x"73",
          4850 => x"9c",
          4851 => x"27",
          4852 => x"75",
          4853 => x"16",
          4854 => x"17",
          4855 => x"33",
          4856 => x"70",
          4857 => x"55",
          4858 => x"80",
          4859 => x"73",
          4860 => x"cc",
          4861 => x"f8",
          4862 => x"81",
          4863 => x"94",
          4864 => x"c8",
          4865 => x"39",
          4866 => x"51",
          4867 => x"81",
          4868 => x"54",
          4869 => x"be",
          4870 => x"27",
          4871 => x"53",
          4872 => x"08",
          4873 => x"73",
          4874 => x"ff",
          4875 => x"15",
          4876 => x"16",
          4877 => x"ff",
          4878 => x"80",
          4879 => x"73",
          4880 => x"c6",
          4881 => x"f8",
          4882 => x"38",
          4883 => x"16",
          4884 => x"80",
          4885 => x"0b",
          4886 => x"81",
          4887 => x"75",
          4888 => x"f8",
          4889 => x"58",
          4890 => x"54",
          4891 => x"74",
          4892 => x"73",
          4893 => x"90",
          4894 => x"c0",
          4895 => x"90",
          4896 => x"83",
          4897 => x"72",
          4898 => x"38",
          4899 => x"08",
          4900 => x"77",
          4901 => x"80",
          4902 => x"f8",
          4903 => x"3d",
          4904 => x"3d",
          4905 => x"89",
          4906 => x"2e",
          4907 => x"80",
          4908 => x"fc",
          4909 => x"3d",
          4910 => x"e1",
          4911 => x"f8",
          4912 => x"81",
          4913 => x"80",
          4914 => x"76",
          4915 => x"75",
          4916 => x"3f",
          4917 => x"08",
          4918 => x"c8",
          4919 => x"38",
          4920 => x"70",
          4921 => x"57",
          4922 => x"a2",
          4923 => x"33",
          4924 => x"70",
          4925 => x"55",
          4926 => x"2e",
          4927 => x"16",
          4928 => x"51",
          4929 => x"81",
          4930 => x"88",
          4931 => x"54",
          4932 => x"84",
          4933 => x"52",
          4934 => x"e5",
          4935 => x"c8",
          4936 => x"84",
          4937 => x"06",
          4938 => x"55",
          4939 => x"80",
          4940 => x"80",
          4941 => x"54",
          4942 => x"c8",
          4943 => x"0d",
          4944 => x"0d",
          4945 => x"fc",
          4946 => x"52",
          4947 => x"3f",
          4948 => x"08",
          4949 => x"f8",
          4950 => x"0c",
          4951 => x"04",
          4952 => x"77",
          4953 => x"fc",
          4954 => x"53",
          4955 => x"de",
          4956 => x"c8",
          4957 => x"f8",
          4958 => x"df",
          4959 => x"38",
          4960 => x"08",
          4961 => x"cd",
          4962 => x"f8",
          4963 => x"80",
          4964 => x"f8",
          4965 => x"73",
          4966 => x"3f",
          4967 => x"08",
          4968 => x"c8",
          4969 => x"09",
          4970 => x"38",
          4971 => x"39",
          4972 => x"08",
          4973 => x"52",
          4974 => x"b3",
          4975 => x"73",
          4976 => x"3f",
          4977 => x"08",
          4978 => x"30",
          4979 => x"9f",
          4980 => x"f8",
          4981 => x"51",
          4982 => x"72",
          4983 => x"0c",
          4984 => x"04",
          4985 => x"65",
          4986 => x"89",
          4987 => x"96",
          4988 => x"df",
          4989 => x"f8",
          4990 => x"81",
          4991 => x"b2",
          4992 => x"75",
          4993 => x"3f",
          4994 => x"08",
          4995 => x"c8",
          4996 => x"02",
          4997 => x"33",
          4998 => x"55",
          4999 => x"25",
          5000 => x"55",
          5001 => x"80",
          5002 => x"76",
          5003 => x"d4",
          5004 => x"81",
          5005 => x"94",
          5006 => x"f0",
          5007 => x"65",
          5008 => x"53",
          5009 => x"05",
          5010 => x"51",
          5011 => x"81",
          5012 => x"5b",
          5013 => x"08",
          5014 => x"7c",
          5015 => x"08",
          5016 => x"fe",
          5017 => x"08",
          5018 => x"55",
          5019 => x"91",
          5020 => x"0c",
          5021 => x"81",
          5022 => x"39",
          5023 => x"c7",
          5024 => x"c8",
          5025 => x"55",
          5026 => x"2e",
          5027 => x"bf",
          5028 => x"5f",
          5029 => x"92",
          5030 => x"51",
          5031 => x"81",
          5032 => x"ff",
          5033 => x"81",
          5034 => x"81",
          5035 => x"81",
          5036 => x"30",
          5037 => x"c8",
          5038 => x"25",
          5039 => x"19",
          5040 => x"5a",
          5041 => x"08",
          5042 => x"38",
          5043 => x"a4",
          5044 => x"f8",
          5045 => x"58",
          5046 => x"77",
          5047 => x"7d",
          5048 => x"bf",
          5049 => x"f8",
          5050 => x"81",
          5051 => x"80",
          5052 => x"70",
          5053 => x"ff",
          5054 => x"56",
          5055 => x"2e",
          5056 => x"9e",
          5057 => x"51",
          5058 => x"3f",
          5059 => x"08",
          5060 => x"06",
          5061 => x"80",
          5062 => x"19",
          5063 => x"54",
          5064 => x"14",
          5065 => x"c5",
          5066 => x"c8",
          5067 => x"06",
          5068 => x"80",
          5069 => x"19",
          5070 => x"54",
          5071 => x"06",
          5072 => x"79",
          5073 => x"78",
          5074 => x"79",
          5075 => x"84",
          5076 => x"07",
          5077 => x"84",
          5078 => x"81",
          5079 => x"92",
          5080 => x"f9",
          5081 => x"8a",
          5082 => x"53",
          5083 => x"e3",
          5084 => x"f8",
          5085 => x"81",
          5086 => x"81",
          5087 => x"17",
          5088 => x"81",
          5089 => x"17",
          5090 => x"2a",
          5091 => x"51",
          5092 => x"55",
          5093 => x"81",
          5094 => x"17",
          5095 => x"8c",
          5096 => x"81",
          5097 => x"9b",
          5098 => x"c8",
          5099 => x"17",
          5100 => x"51",
          5101 => x"81",
          5102 => x"74",
          5103 => x"56",
          5104 => x"98",
          5105 => x"76",
          5106 => x"c6",
          5107 => x"c8",
          5108 => x"09",
          5109 => x"38",
          5110 => x"f8",
          5111 => x"2e",
          5112 => x"85",
          5113 => x"a3",
          5114 => x"38",
          5115 => x"f8",
          5116 => x"15",
          5117 => x"38",
          5118 => x"53",
          5119 => x"08",
          5120 => x"c3",
          5121 => x"f8",
          5122 => x"94",
          5123 => x"18",
          5124 => x"33",
          5125 => x"54",
          5126 => x"34",
          5127 => x"85",
          5128 => x"18",
          5129 => x"74",
          5130 => x"0c",
          5131 => x"04",
          5132 => x"82",
          5133 => x"ff",
          5134 => x"a1",
          5135 => x"e4",
          5136 => x"c8",
          5137 => x"f8",
          5138 => x"f5",
          5139 => x"a1",
          5140 => x"95",
          5141 => x"58",
          5142 => x"81",
          5143 => x"55",
          5144 => x"08",
          5145 => x"02",
          5146 => x"33",
          5147 => x"70",
          5148 => x"55",
          5149 => x"73",
          5150 => x"75",
          5151 => x"80",
          5152 => x"bd",
          5153 => x"d6",
          5154 => x"81",
          5155 => x"87",
          5156 => x"ad",
          5157 => x"78",
          5158 => x"3f",
          5159 => x"08",
          5160 => x"70",
          5161 => x"55",
          5162 => x"2e",
          5163 => x"78",
          5164 => x"c8",
          5165 => x"08",
          5166 => x"38",
          5167 => x"f8",
          5168 => x"76",
          5169 => x"70",
          5170 => x"b5",
          5171 => x"c8",
          5172 => x"f8",
          5173 => x"e9",
          5174 => x"c8",
          5175 => x"51",
          5176 => x"81",
          5177 => x"55",
          5178 => x"08",
          5179 => x"55",
          5180 => x"81",
          5181 => x"84",
          5182 => x"81",
          5183 => x"80",
          5184 => x"51",
          5185 => x"81",
          5186 => x"81",
          5187 => x"30",
          5188 => x"c8",
          5189 => x"25",
          5190 => x"75",
          5191 => x"38",
          5192 => x"8f",
          5193 => x"75",
          5194 => x"c1",
          5195 => x"f8",
          5196 => x"74",
          5197 => x"51",
          5198 => x"3f",
          5199 => x"08",
          5200 => x"f8",
          5201 => x"3d",
          5202 => x"3d",
          5203 => x"99",
          5204 => x"52",
          5205 => x"d8",
          5206 => x"f8",
          5207 => x"81",
          5208 => x"82",
          5209 => x"5e",
          5210 => x"3d",
          5211 => x"cf",
          5212 => x"f8",
          5213 => x"81",
          5214 => x"86",
          5215 => x"82",
          5216 => x"f8",
          5217 => x"2e",
          5218 => x"82",
          5219 => x"80",
          5220 => x"70",
          5221 => x"06",
          5222 => x"54",
          5223 => x"38",
          5224 => x"52",
          5225 => x"52",
          5226 => x"3f",
          5227 => x"08",
          5228 => x"81",
          5229 => x"83",
          5230 => x"81",
          5231 => x"81",
          5232 => x"06",
          5233 => x"54",
          5234 => x"08",
          5235 => x"81",
          5236 => x"81",
          5237 => x"39",
          5238 => x"38",
          5239 => x"08",
          5240 => x"c4",
          5241 => x"f8",
          5242 => x"81",
          5243 => x"81",
          5244 => x"53",
          5245 => x"19",
          5246 => x"8c",
          5247 => x"ae",
          5248 => x"34",
          5249 => x"0b",
          5250 => x"82",
          5251 => x"52",
          5252 => x"51",
          5253 => x"3f",
          5254 => x"b4",
          5255 => x"c9",
          5256 => x"53",
          5257 => x"53",
          5258 => x"51",
          5259 => x"3f",
          5260 => x"0b",
          5261 => x"34",
          5262 => x"80",
          5263 => x"51",
          5264 => x"78",
          5265 => x"83",
          5266 => x"51",
          5267 => x"81",
          5268 => x"54",
          5269 => x"08",
          5270 => x"88",
          5271 => x"64",
          5272 => x"ff",
          5273 => x"75",
          5274 => x"78",
          5275 => x"3f",
          5276 => x"0b",
          5277 => x"78",
          5278 => x"83",
          5279 => x"51",
          5280 => x"3f",
          5281 => x"08",
          5282 => x"80",
          5283 => x"76",
          5284 => x"ae",
          5285 => x"f8",
          5286 => x"3d",
          5287 => x"3d",
          5288 => x"84",
          5289 => x"f1",
          5290 => x"a8",
          5291 => x"05",
          5292 => x"51",
          5293 => x"81",
          5294 => x"55",
          5295 => x"08",
          5296 => x"78",
          5297 => x"08",
          5298 => x"70",
          5299 => x"b8",
          5300 => x"c8",
          5301 => x"f8",
          5302 => x"b9",
          5303 => x"9b",
          5304 => x"a0",
          5305 => x"55",
          5306 => x"38",
          5307 => x"3d",
          5308 => x"3d",
          5309 => x"51",
          5310 => x"3f",
          5311 => x"52",
          5312 => x"52",
          5313 => x"dd",
          5314 => x"08",
          5315 => x"cb",
          5316 => x"f8",
          5317 => x"81",
          5318 => x"95",
          5319 => x"2e",
          5320 => x"88",
          5321 => x"3d",
          5322 => x"38",
          5323 => x"e5",
          5324 => x"c8",
          5325 => x"09",
          5326 => x"b8",
          5327 => x"c9",
          5328 => x"f8",
          5329 => x"81",
          5330 => x"81",
          5331 => x"56",
          5332 => x"3d",
          5333 => x"52",
          5334 => x"ff",
          5335 => x"02",
          5336 => x"8b",
          5337 => x"16",
          5338 => x"2a",
          5339 => x"51",
          5340 => x"89",
          5341 => x"07",
          5342 => x"17",
          5343 => x"81",
          5344 => x"34",
          5345 => x"70",
          5346 => x"81",
          5347 => x"55",
          5348 => x"80",
          5349 => x"64",
          5350 => x"38",
          5351 => x"51",
          5352 => x"81",
          5353 => x"52",
          5354 => x"b7",
          5355 => x"55",
          5356 => x"08",
          5357 => x"dd",
          5358 => x"c8",
          5359 => x"51",
          5360 => x"3f",
          5361 => x"08",
          5362 => x"11",
          5363 => x"81",
          5364 => x"80",
          5365 => x"16",
          5366 => x"ae",
          5367 => x"06",
          5368 => x"53",
          5369 => x"51",
          5370 => x"78",
          5371 => x"83",
          5372 => x"39",
          5373 => x"08",
          5374 => x"51",
          5375 => x"81",
          5376 => x"55",
          5377 => x"08",
          5378 => x"51",
          5379 => x"3f",
          5380 => x"08",
          5381 => x"f8",
          5382 => x"3d",
          5383 => x"3d",
          5384 => x"db",
          5385 => x"84",
          5386 => x"05",
          5387 => x"82",
          5388 => x"d0",
          5389 => x"3d",
          5390 => x"3f",
          5391 => x"08",
          5392 => x"c8",
          5393 => x"38",
          5394 => x"52",
          5395 => x"05",
          5396 => x"3f",
          5397 => x"08",
          5398 => x"c8",
          5399 => x"02",
          5400 => x"33",
          5401 => x"54",
          5402 => x"aa",
          5403 => x"06",
          5404 => x"8b",
          5405 => x"06",
          5406 => x"07",
          5407 => x"56",
          5408 => x"34",
          5409 => x"0b",
          5410 => x"78",
          5411 => x"a9",
          5412 => x"c8",
          5413 => x"81",
          5414 => x"95",
          5415 => x"ef",
          5416 => x"56",
          5417 => x"3d",
          5418 => x"94",
          5419 => x"f4",
          5420 => x"c8",
          5421 => x"f8",
          5422 => x"cb",
          5423 => x"63",
          5424 => x"d4",
          5425 => x"c0",
          5426 => x"c8",
          5427 => x"f8",
          5428 => x"38",
          5429 => x"05",
          5430 => x"06",
          5431 => x"73",
          5432 => x"16",
          5433 => x"22",
          5434 => x"07",
          5435 => x"1f",
          5436 => x"c2",
          5437 => x"81",
          5438 => x"34",
          5439 => x"b3",
          5440 => x"f8",
          5441 => x"74",
          5442 => x"0c",
          5443 => x"04",
          5444 => x"69",
          5445 => x"80",
          5446 => x"d0",
          5447 => x"3d",
          5448 => x"3f",
          5449 => x"08",
          5450 => x"08",
          5451 => x"f8",
          5452 => x"80",
          5453 => x"57",
          5454 => x"81",
          5455 => x"70",
          5456 => x"55",
          5457 => x"80",
          5458 => x"5d",
          5459 => x"52",
          5460 => x"52",
          5461 => x"a9",
          5462 => x"c8",
          5463 => x"f8",
          5464 => x"d1",
          5465 => x"73",
          5466 => x"3f",
          5467 => x"08",
          5468 => x"c8",
          5469 => x"81",
          5470 => x"81",
          5471 => x"65",
          5472 => x"78",
          5473 => x"7b",
          5474 => x"55",
          5475 => x"34",
          5476 => x"8a",
          5477 => x"38",
          5478 => x"1a",
          5479 => x"34",
          5480 => x"9e",
          5481 => x"70",
          5482 => x"51",
          5483 => x"a0",
          5484 => x"8e",
          5485 => x"2e",
          5486 => x"86",
          5487 => x"34",
          5488 => x"30",
          5489 => x"80",
          5490 => x"7a",
          5491 => x"c1",
          5492 => x"2e",
          5493 => x"a0",
          5494 => x"51",
          5495 => x"3f",
          5496 => x"08",
          5497 => x"c8",
          5498 => x"7b",
          5499 => x"55",
          5500 => x"73",
          5501 => x"38",
          5502 => x"73",
          5503 => x"38",
          5504 => x"15",
          5505 => x"ff",
          5506 => x"81",
          5507 => x"7b",
          5508 => x"f8",
          5509 => x"3d",
          5510 => x"3d",
          5511 => x"9c",
          5512 => x"05",
          5513 => x"51",
          5514 => x"81",
          5515 => x"81",
          5516 => x"56",
          5517 => x"c8",
          5518 => x"38",
          5519 => x"52",
          5520 => x"52",
          5521 => x"c0",
          5522 => x"70",
          5523 => x"ff",
          5524 => x"55",
          5525 => x"27",
          5526 => x"78",
          5527 => x"ff",
          5528 => x"05",
          5529 => x"55",
          5530 => x"3f",
          5531 => x"08",
          5532 => x"38",
          5533 => x"70",
          5534 => x"ff",
          5535 => x"81",
          5536 => x"80",
          5537 => x"74",
          5538 => x"07",
          5539 => x"4e",
          5540 => x"81",
          5541 => x"55",
          5542 => x"70",
          5543 => x"06",
          5544 => x"99",
          5545 => x"e0",
          5546 => x"ff",
          5547 => x"54",
          5548 => x"27",
          5549 => x"e5",
          5550 => x"55",
          5551 => x"a3",
          5552 => x"81",
          5553 => x"ff",
          5554 => x"81",
          5555 => x"93",
          5556 => x"75",
          5557 => x"76",
          5558 => x"38",
          5559 => x"77",
          5560 => x"86",
          5561 => x"39",
          5562 => x"27",
          5563 => x"88",
          5564 => x"78",
          5565 => x"5a",
          5566 => x"57",
          5567 => x"81",
          5568 => x"81",
          5569 => x"33",
          5570 => x"06",
          5571 => x"57",
          5572 => x"fe",
          5573 => x"3d",
          5574 => x"55",
          5575 => x"2e",
          5576 => x"76",
          5577 => x"38",
          5578 => x"55",
          5579 => x"33",
          5580 => x"a0",
          5581 => x"06",
          5582 => x"17",
          5583 => x"38",
          5584 => x"43",
          5585 => x"3d",
          5586 => x"ff",
          5587 => x"81",
          5588 => x"54",
          5589 => x"08",
          5590 => x"81",
          5591 => x"ff",
          5592 => x"81",
          5593 => x"54",
          5594 => x"08",
          5595 => x"80",
          5596 => x"54",
          5597 => x"80",
          5598 => x"f8",
          5599 => x"2e",
          5600 => x"80",
          5601 => x"54",
          5602 => x"80",
          5603 => x"52",
          5604 => x"bd",
          5605 => x"f8",
          5606 => x"81",
          5607 => x"b1",
          5608 => x"81",
          5609 => x"52",
          5610 => x"ab",
          5611 => x"54",
          5612 => x"15",
          5613 => x"78",
          5614 => x"ff",
          5615 => x"79",
          5616 => x"83",
          5617 => x"51",
          5618 => x"3f",
          5619 => x"08",
          5620 => x"74",
          5621 => x"0c",
          5622 => x"04",
          5623 => x"60",
          5624 => x"05",
          5625 => x"33",
          5626 => x"05",
          5627 => x"40",
          5628 => x"da",
          5629 => x"c8",
          5630 => x"f8",
          5631 => x"bd",
          5632 => x"33",
          5633 => x"b5",
          5634 => x"2e",
          5635 => x"1a",
          5636 => x"90",
          5637 => x"33",
          5638 => x"70",
          5639 => x"55",
          5640 => x"38",
          5641 => x"97",
          5642 => x"82",
          5643 => x"58",
          5644 => x"7e",
          5645 => x"70",
          5646 => x"55",
          5647 => x"56",
          5648 => x"e8",
          5649 => x"7d",
          5650 => x"70",
          5651 => x"2a",
          5652 => x"08",
          5653 => x"08",
          5654 => x"5d",
          5655 => x"77",
          5656 => x"98",
          5657 => x"26",
          5658 => x"57",
          5659 => x"59",
          5660 => x"52",
          5661 => x"ae",
          5662 => x"15",
          5663 => x"98",
          5664 => x"26",
          5665 => x"55",
          5666 => x"08",
          5667 => x"99",
          5668 => x"c8",
          5669 => x"ff",
          5670 => x"f8",
          5671 => x"38",
          5672 => x"75",
          5673 => x"81",
          5674 => x"93",
          5675 => x"80",
          5676 => x"2e",
          5677 => x"ff",
          5678 => x"58",
          5679 => x"7d",
          5680 => x"38",
          5681 => x"55",
          5682 => x"b4",
          5683 => x"56",
          5684 => x"09",
          5685 => x"38",
          5686 => x"53",
          5687 => x"51",
          5688 => x"3f",
          5689 => x"08",
          5690 => x"c8",
          5691 => x"38",
          5692 => x"ff",
          5693 => x"5c",
          5694 => x"84",
          5695 => x"5c",
          5696 => x"12",
          5697 => x"80",
          5698 => x"78",
          5699 => x"7c",
          5700 => x"90",
          5701 => x"c0",
          5702 => x"90",
          5703 => x"15",
          5704 => x"90",
          5705 => x"54",
          5706 => x"91",
          5707 => x"31",
          5708 => x"84",
          5709 => x"07",
          5710 => x"16",
          5711 => x"73",
          5712 => x"0c",
          5713 => x"04",
          5714 => x"6b",
          5715 => x"05",
          5716 => x"33",
          5717 => x"5a",
          5718 => x"bd",
          5719 => x"80",
          5720 => x"c8",
          5721 => x"f8",
          5722 => x"c8",
          5723 => x"81",
          5724 => x"70",
          5725 => x"74",
          5726 => x"38",
          5727 => x"81",
          5728 => x"81",
          5729 => x"81",
          5730 => x"ff",
          5731 => x"81",
          5732 => x"81",
          5733 => x"81",
          5734 => x"83",
          5735 => x"c0",
          5736 => x"2a",
          5737 => x"51",
          5738 => x"74",
          5739 => x"99",
          5740 => x"53",
          5741 => x"51",
          5742 => x"3f",
          5743 => x"08",
          5744 => x"55",
          5745 => x"92",
          5746 => x"80",
          5747 => x"38",
          5748 => x"06",
          5749 => x"2e",
          5750 => x"48",
          5751 => x"87",
          5752 => x"79",
          5753 => x"78",
          5754 => x"26",
          5755 => x"19",
          5756 => x"74",
          5757 => x"38",
          5758 => x"e4",
          5759 => x"2a",
          5760 => x"70",
          5761 => x"59",
          5762 => x"7a",
          5763 => x"56",
          5764 => x"80",
          5765 => x"51",
          5766 => x"74",
          5767 => x"99",
          5768 => x"53",
          5769 => x"51",
          5770 => x"3f",
          5771 => x"f8",
          5772 => x"ac",
          5773 => x"2a",
          5774 => x"81",
          5775 => x"43",
          5776 => x"83",
          5777 => x"66",
          5778 => x"60",
          5779 => x"90",
          5780 => x"31",
          5781 => x"80",
          5782 => x"8a",
          5783 => x"56",
          5784 => x"26",
          5785 => x"77",
          5786 => x"81",
          5787 => x"74",
          5788 => x"38",
          5789 => x"55",
          5790 => x"83",
          5791 => x"81",
          5792 => x"80",
          5793 => x"38",
          5794 => x"55",
          5795 => x"5e",
          5796 => x"89",
          5797 => x"5a",
          5798 => x"09",
          5799 => x"e1",
          5800 => x"38",
          5801 => x"57",
          5802 => x"e7",
          5803 => x"5a",
          5804 => x"9d",
          5805 => x"26",
          5806 => x"e7",
          5807 => x"10",
          5808 => x"22",
          5809 => x"74",
          5810 => x"38",
          5811 => x"ee",
          5812 => x"66",
          5813 => x"d4",
          5814 => x"c8",
          5815 => x"84",
          5816 => x"89",
          5817 => x"a0",
          5818 => x"81",
          5819 => x"fc",
          5820 => x"56",
          5821 => x"f0",
          5822 => x"80",
          5823 => x"d3",
          5824 => x"38",
          5825 => x"57",
          5826 => x"e7",
          5827 => x"5a",
          5828 => x"9d",
          5829 => x"26",
          5830 => x"e7",
          5831 => x"10",
          5832 => x"22",
          5833 => x"74",
          5834 => x"38",
          5835 => x"ee",
          5836 => x"66",
          5837 => x"f4",
          5838 => x"c8",
          5839 => x"05",
          5840 => x"c8",
          5841 => x"26",
          5842 => x"0b",
          5843 => x"08",
          5844 => x"c8",
          5845 => x"11",
          5846 => x"05",
          5847 => x"83",
          5848 => x"2a",
          5849 => x"a0",
          5850 => x"7d",
          5851 => x"69",
          5852 => x"05",
          5853 => x"72",
          5854 => x"5c",
          5855 => x"59",
          5856 => x"2e",
          5857 => x"89",
          5858 => x"60",
          5859 => x"84",
          5860 => x"5d",
          5861 => x"18",
          5862 => x"68",
          5863 => x"74",
          5864 => x"af",
          5865 => x"31",
          5866 => x"53",
          5867 => x"52",
          5868 => x"f8",
          5869 => x"c8",
          5870 => x"83",
          5871 => x"06",
          5872 => x"f8",
          5873 => x"ff",
          5874 => x"dd",
          5875 => x"83",
          5876 => x"2a",
          5877 => x"be",
          5878 => x"39",
          5879 => x"09",
          5880 => x"c5",
          5881 => x"f5",
          5882 => x"c8",
          5883 => x"38",
          5884 => x"79",
          5885 => x"80",
          5886 => x"38",
          5887 => x"96",
          5888 => x"06",
          5889 => x"2e",
          5890 => x"5e",
          5891 => x"81",
          5892 => x"9f",
          5893 => x"38",
          5894 => x"38",
          5895 => x"81",
          5896 => x"fc",
          5897 => x"ab",
          5898 => x"7d",
          5899 => x"81",
          5900 => x"7d",
          5901 => x"78",
          5902 => x"74",
          5903 => x"8e",
          5904 => x"9c",
          5905 => x"53",
          5906 => x"51",
          5907 => x"3f",
          5908 => x"e6",
          5909 => x"51",
          5910 => x"3f",
          5911 => x"8b",
          5912 => x"a1",
          5913 => x"8d",
          5914 => x"83",
          5915 => x"52",
          5916 => x"ff",
          5917 => x"81",
          5918 => x"34",
          5919 => x"70",
          5920 => x"2a",
          5921 => x"54",
          5922 => x"1b",
          5923 => x"88",
          5924 => x"74",
          5925 => x"26",
          5926 => x"83",
          5927 => x"52",
          5928 => x"ff",
          5929 => x"8a",
          5930 => x"a0",
          5931 => x"a1",
          5932 => x"0b",
          5933 => x"bf",
          5934 => x"51",
          5935 => x"3f",
          5936 => x"9a",
          5937 => x"a0",
          5938 => x"52",
          5939 => x"ff",
          5940 => x"7d",
          5941 => x"81",
          5942 => x"38",
          5943 => x"0a",
          5944 => x"1b",
          5945 => x"ce",
          5946 => x"a4",
          5947 => x"a0",
          5948 => x"52",
          5949 => x"ff",
          5950 => x"81",
          5951 => x"51",
          5952 => x"3f",
          5953 => x"1b",
          5954 => x"8c",
          5955 => x"0b",
          5956 => x"34",
          5957 => x"c2",
          5958 => x"53",
          5959 => x"52",
          5960 => x"51",
          5961 => x"88",
          5962 => x"a7",
          5963 => x"a0",
          5964 => x"83",
          5965 => x"52",
          5966 => x"ff",
          5967 => x"ff",
          5968 => x"1c",
          5969 => x"a6",
          5970 => x"53",
          5971 => x"52",
          5972 => x"ff",
          5973 => x"82",
          5974 => x"83",
          5975 => x"52",
          5976 => x"b4",
          5977 => x"60",
          5978 => x"7e",
          5979 => x"d7",
          5980 => x"81",
          5981 => x"83",
          5982 => x"83",
          5983 => x"06",
          5984 => x"75",
          5985 => x"05",
          5986 => x"7e",
          5987 => x"b7",
          5988 => x"53",
          5989 => x"51",
          5990 => x"3f",
          5991 => x"a4",
          5992 => x"51",
          5993 => x"3f",
          5994 => x"e4",
          5995 => x"e4",
          5996 => x"9f",
          5997 => x"18",
          5998 => x"1b",
          5999 => x"f6",
          6000 => x"83",
          6001 => x"ff",
          6002 => x"82",
          6003 => x"78",
          6004 => x"c4",
          6005 => x"60",
          6006 => x"7a",
          6007 => x"ff",
          6008 => x"75",
          6009 => x"53",
          6010 => x"51",
          6011 => x"3f",
          6012 => x"52",
          6013 => x"9f",
          6014 => x"56",
          6015 => x"83",
          6016 => x"06",
          6017 => x"52",
          6018 => x"9e",
          6019 => x"52",
          6020 => x"ff",
          6021 => x"f0",
          6022 => x"1b",
          6023 => x"87",
          6024 => x"55",
          6025 => x"83",
          6026 => x"74",
          6027 => x"ff",
          6028 => x"7c",
          6029 => x"74",
          6030 => x"38",
          6031 => x"54",
          6032 => x"52",
          6033 => x"99",
          6034 => x"f8",
          6035 => x"87",
          6036 => x"53",
          6037 => x"08",
          6038 => x"ff",
          6039 => x"76",
          6040 => x"31",
          6041 => x"cd",
          6042 => x"58",
          6043 => x"ff",
          6044 => x"55",
          6045 => x"83",
          6046 => x"61",
          6047 => x"26",
          6048 => x"57",
          6049 => x"53",
          6050 => x"51",
          6051 => x"3f",
          6052 => x"08",
          6053 => x"76",
          6054 => x"31",
          6055 => x"db",
          6056 => x"7d",
          6057 => x"38",
          6058 => x"83",
          6059 => x"8a",
          6060 => x"7d",
          6061 => x"38",
          6062 => x"81",
          6063 => x"80",
          6064 => x"80",
          6065 => x"7a",
          6066 => x"bc",
          6067 => x"d5",
          6068 => x"ff",
          6069 => x"83",
          6070 => x"77",
          6071 => x"0b",
          6072 => x"81",
          6073 => x"34",
          6074 => x"34",
          6075 => x"34",
          6076 => x"56",
          6077 => x"52",
          6078 => x"d5",
          6079 => x"0b",
          6080 => x"81",
          6081 => x"82",
          6082 => x"56",
          6083 => x"34",
          6084 => x"08",
          6085 => x"60",
          6086 => x"1b",
          6087 => x"96",
          6088 => x"83",
          6089 => x"ff",
          6090 => x"81",
          6091 => x"7a",
          6092 => x"ff",
          6093 => x"81",
          6094 => x"c8",
          6095 => x"80",
          6096 => x"7e",
          6097 => x"e3",
          6098 => x"81",
          6099 => x"90",
          6100 => x"8e",
          6101 => x"81",
          6102 => x"81",
          6103 => x"56",
          6104 => x"c8",
          6105 => x"0d",
          6106 => x"0d",
          6107 => x"59",
          6108 => x"ff",
          6109 => x"57",
          6110 => x"b4",
          6111 => x"f8",
          6112 => x"81",
          6113 => x"52",
          6114 => x"dc",
          6115 => x"2e",
          6116 => x"9c",
          6117 => x"33",
          6118 => x"2e",
          6119 => x"76",
          6120 => x"58",
          6121 => x"57",
          6122 => x"09",
          6123 => x"38",
          6124 => x"78",
          6125 => x"38",
          6126 => x"81",
          6127 => x"8d",
          6128 => x"f7",
          6129 => x"02",
          6130 => x"05",
          6131 => x"77",
          6132 => x"81",
          6133 => x"8d",
          6134 => x"e7",
          6135 => x"08",
          6136 => x"24",
          6137 => x"17",
          6138 => x"8c",
          6139 => x"77",
          6140 => x"16",
          6141 => x"25",
          6142 => x"3d",
          6143 => x"75",
          6144 => x"52",
          6145 => x"cb",
          6146 => x"76",
          6147 => x"70",
          6148 => x"2a",
          6149 => x"51",
          6150 => x"84",
          6151 => x"19",
          6152 => x"8b",
          6153 => x"f9",
          6154 => x"84",
          6155 => x"56",
          6156 => x"a7",
          6157 => x"fc",
          6158 => x"53",
          6159 => x"75",
          6160 => x"a1",
          6161 => x"c8",
          6162 => x"84",
          6163 => x"2e",
          6164 => x"87",
          6165 => x"08",
          6166 => x"ff",
          6167 => x"f8",
          6168 => x"3d",
          6169 => x"3d",
          6170 => x"80",
          6171 => x"52",
          6172 => x"9a",
          6173 => x"74",
          6174 => x"0d",
          6175 => x"0d",
          6176 => x"05",
          6177 => x"86",
          6178 => x"54",
          6179 => x"73",
          6180 => x"fe",
          6181 => x"51",
          6182 => x"98",
          6183 => x"f8",
          6184 => x"70",
          6185 => x"56",
          6186 => x"2e",
          6187 => x"8c",
          6188 => x"79",
          6189 => x"33",
          6190 => x"39",
          6191 => x"73",
          6192 => x"81",
          6193 => x"81",
          6194 => x"39",
          6195 => x"90",
          6196 => x"b8",
          6197 => x"52",
          6198 => x"f2",
          6199 => x"c8",
          6200 => x"c8",
          6201 => x"53",
          6202 => x"58",
          6203 => x"3f",
          6204 => x"08",
          6205 => x"16",
          6206 => x"81",
          6207 => x"38",
          6208 => x"81",
          6209 => x"54",
          6210 => x"c2",
          6211 => x"73",
          6212 => x"0c",
          6213 => x"04",
          6214 => x"73",
          6215 => x"26",
          6216 => x"71",
          6217 => x"dd",
          6218 => x"71",
          6219 => x"e9",
          6220 => x"80",
          6221 => x"c0",
          6222 => x"39",
          6223 => x"51",
          6224 => x"81",
          6225 => x"80",
          6226 => x"e9",
          6227 => x"e4",
          6228 => x"88",
          6229 => x"39",
          6230 => x"51",
          6231 => x"81",
          6232 => x"80",
          6233 => x"ea",
          6234 => x"c8",
          6235 => x"dc",
          6236 => x"39",
          6237 => x"51",
          6238 => x"eb",
          6239 => x"39",
          6240 => x"51",
          6241 => x"eb",
          6242 => x"39",
          6243 => x"51",
          6244 => x"ec",
          6245 => x"39",
          6246 => x"51",
          6247 => x"ec",
          6248 => x"39",
          6249 => x"51",
          6250 => x"ec",
          6251 => x"39",
          6252 => x"51",
          6253 => x"3f",
          6254 => x"04",
          6255 => x"77",
          6256 => x"74",
          6257 => x"8a",
          6258 => x"75",
          6259 => x"51",
          6260 => x"e8",
          6261 => x"fe",
          6262 => x"81",
          6263 => x"52",
          6264 => x"cf",
          6265 => x"f8",
          6266 => x"79",
          6267 => x"81",
          6268 => x"fe",
          6269 => x"87",
          6270 => x"ec",
          6271 => x"02",
          6272 => x"e3",
          6273 => x"57",
          6274 => x"30",
          6275 => x"73",
          6276 => x"59",
          6277 => x"77",
          6278 => x"83",
          6279 => x"74",
          6280 => x"81",
          6281 => x"55",
          6282 => x"81",
          6283 => x"53",
          6284 => x"3d",
          6285 => x"ff",
          6286 => x"81",
          6287 => x"57",
          6288 => x"08",
          6289 => x"f8",
          6290 => x"c0",
          6291 => x"81",
          6292 => x"59",
          6293 => x"05",
          6294 => x"53",
          6295 => x"51",
          6296 => x"81",
          6297 => x"57",
          6298 => x"08",
          6299 => x"55",
          6300 => x"89",
          6301 => x"75",
          6302 => x"d8",
          6303 => x"d8",
          6304 => x"f0",
          6305 => x"70",
          6306 => x"25",
          6307 => x"9f",
          6308 => x"51",
          6309 => x"74",
          6310 => x"38",
          6311 => x"53",
          6312 => x"88",
          6313 => x"51",
          6314 => x"76",
          6315 => x"f8",
          6316 => x"3d",
          6317 => x"3d",
          6318 => x"84",
          6319 => x"33",
          6320 => x"57",
          6321 => x"52",
          6322 => x"af",
          6323 => x"c8",
          6324 => x"75",
          6325 => x"38",
          6326 => x"98",
          6327 => x"60",
          6328 => x"81",
          6329 => x"7e",
          6330 => x"77",
          6331 => x"c8",
          6332 => x"39",
          6333 => x"81",
          6334 => x"89",
          6335 => x"f3",
          6336 => x"61",
          6337 => x"05",
          6338 => x"33",
          6339 => x"68",
          6340 => x"5c",
          6341 => x"7a",
          6342 => x"a8",
          6343 => x"a9",
          6344 => x"b0",
          6345 => x"bd",
          6346 => x"74",
          6347 => x"fc",
          6348 => x"2e",
          6349 => x"a0",
          6350 => x"80",
          6351 => x"18",
          6352 => x"27",
          6353 => x"22",
          6354 => x"b4",
          6355 => x"f9",
          6356 => x"81",
          6357 => x"fe",
          6358 => x"82",
          6359 => x"c3",
          6360 => x"53",
          6361 => x"8e",
          6362 => x"52",
          6363 => x"51",
          6364 => x"3f",
          6365 => x"ed",
          6366 => x"ee",
          6367 => x"15",
          6368 => x"74",
          6369 => x"7a",
          6370 => x"72",
          6371 => x"ed",
          6372 => x"f4",
          6373 => x"39",
          6374 => x"51",
          6375 => x"3f",
          6376 => x"a0",
          6377 => x"e0",
          6378 => x"39",
          6379 => x"51",
          6380 => x"3f",
          6381 => x"79",
          6382 => x"74",
          6383 => x"55",
          6384 => x"72",
          6385 => x"38",
          6386 => x"53",
          6387 => x"83",
          6388 => x"75",
          6389 => x"81",
          6390 => x"53",
          6391 => x"8b",
          6392 => x"fe",
          6393 => x"73",
          6394 => x"a0",
          6395 => x"98",
          6396 => x"55",
          6397 => x"ed",
          6398 => x"ed",
          6399 => x"18",
          6400 => x"58",
          6401 => x"3f",
          6402 => x"08",
          6403 => x"98",
          6404 => x"76",
          6405 => x"81",
          6406 => x"fe",
          6407 => x"81",
          6408 => x"98",
          6409 => x"2c",
          6410 => x"70",
          6411 => x"32",
          6412 => x"72",
          6413 => x"07",
          6414 => x"58",
          6415 => x"57",
          6416 => x"d7",
          6417 => x"2e",
          6418 => x"85",
          6419 => x"8c",
          6420 => x"53",
          6421 => x"fd",
          6422 => x"53",
          6423 => x"c8",
          6424 => x"0d",
          6425 => x"0d",
          6426 => x"33",
          6427 => x"53",
          6428 => x"52",
          6429 => x"d1",
          6430 => x"f8",
          6431 => x"e7",
          6432 => x"ed",
          6433 => x"ed",
          6434 => x"f3",
          6435 => x"81",
          6436 => x"fe",
          6437 => x"74",
          6438 => x"38",
          6439 => x"3f",
          6440 => x"04",
          6441 => x"87",
          6442 => x"08",
          6443 => x"b1",
          6444 => x"fe",
          6445 => x"81",
          6446 => x"fe",
          6447 => x"80",
          6448 => x"ae",
          6449 => x"2a",
          6450 => x"51",
          6451 => x"2e",
          6452 => x"51",
          6453 => x"3f",
          6454 => x"51",
          6455 => x"3f",
          6456 => x"d9",
          6457 => x"82",
          6458 => x"06",
          6459 => x"80",
          6460 => x"81",
          6461 => x"fa",
          6462 => x"c8",
          6463 => x"f2",
          6464 => x"fe",
          6465 => x"72",
          6466 => x"81",
          6467 => x"71",
          6468 => x"38",
          6469 => x"d8",
          6470 => x"ee",
          6471 => x"da",
          6472 => x"51",
          6473 => x"3f",
          6474 => x"70",
          6475 => x"52",
          6476 => x"95",
          6477 => x"fe",
          6478 => x"81",
          6479 => x"fe",
          6480 => x"80",
          6481 => x"aa",
          6482 => x"2a",
          6483 => x"51",
          6484 => x"2e",
          6485 => x"51",
          6486 => x"3f",
          6487 => x"51",
          6488 => x"3f",
          6489 => x"d8",
          6490 => x"86",
          6491 => x"06",
          6492 => x"80",
          6493 => x"81",
          6494 => x"f6",
          6495 => x"94",
          6496 => x"ee",
          6497 => x"fe",
          6498 => x"72",
          6499 => x"81",
          6500 => x"71",
          6501 => x"38",
          6502 => x"d7",
          6503 => x"ef",
          6504 => x"d9",
          6505 => x"51",
          6506 => x"3f",
          6507 => x"70",
          6508 => x"52",
          6509 => x"95",
          6510 => x"fe",
          6511 => x"81",
          6512 => x"fe",
          6513 => x"80",
          6514 => x"a6",
          6515 => x"99",
          6516 => x"0d",
          6517 => x"0d",
          6518 => x"05",
          6519 => x"70",
          6520 => x"80",
          6521 => x"fe",
          6522 => x"81",
          6523 => x"54",
          6524 => x"81",
          6525 => x"fc",
          6526 => x"e0",
          6527 => x"83",
          6528 => x"c8",
          6529 => x"81",
          6530 => x"07",
          6531 => x"71",
          6532 => x"54",
          6533 => x"b4",
          6534 => x"b4",
          6535 => x"81",
          6536 => x"06",
          6537 => x"8f",
          6538 => x"52",
          6539 => x"b9",
          6540 => x"c8",
          6541 => x"8c",
          6542 => x"c8",
          6543 => x"e9",
          6544 => x"39",
          6545 => x"51",
          6546 => x"82",
          6547 => x"b4",
          6548 => x"b4",
          6549 => x"82",
          6550 => x"06",
          6551 => x"52",
          6552 => x"fa",
          6553 => x"0b",
          6554 => x"0c",
          6555 => x"04",
          6556 => x"80",
          6557 => x"8f",
          6558 => x"5d",
          6559 => x"51",
          6560 => x"3f",
          6561 => x"08",
          6562 => x"59",
          6563 => x"09",
          6564 => x"38",
          6565 => x"52",
          6566 => x"52",
          6567 => x"bf",
          6568 => x"78",
          6569 => x"8c",
          6570 => x"f6",
          6571 => x"c8",
          6572 => x"88",
          6573 => x"90",
          6574 => x"39",
          6575 => x"5d",
          6576 => x"51",
          6577 => x"3f",
          6578 => x"46",
          6579 => x"52",
          6580 => x"81",
          6581 => x"ff",
          6582 => x"f3",
          6583 => x"f8",
          6584 => x"2b",
          6585 => x"51",
          6586 => x"c2",
          6587 => x"38",
          6588 => x"24",
          6589 => x"bd",
          6590 => x"38",
          6591 => x"90",
          6592 => x"2e",
          6593 => x"78",
          6594 => x"da",
          6595 => x"39",
          6596 => x"2e",
          6597 => x"78",
          6598 => x"85",
          6599 => x"bf",
          6600 => x"38",
          6601 => x"78",
          6602 => x"89",
          6603 => x"80",
          6604 => x"38",
          6605 => x"2e",
          6606 => x"78",
          6607 => x"89",
          6608 => x"b4",
          6609 => x"83",
          6610 => x"38",
          6611 => x"24",
          6612 => x"81",
          6613 => x"fd",
          6614 => x"39",
          6615 => x"2e",
          6616 => x"8a",
          6617 => x"3d",
          6618 => x"53",
          6619 => x"51",
          6620 => x"3f",
          6621 => x"08",
          6622 => x"c4",
          6623 => x"fe",
          6624 => x"ff",
          6625 => x"fe",
          6626 => x"81",
          6627 => x"80",
          6628 => x"38",
          6629 => x"f8",
          6630 => x"84",
          6631 => x"ee",
          6632 => x"f8",
          6633 => x"38",
          6634 => x"08",
          6635 => x"cc",
          6636 => x"b1",
          6637 => x"5c",
          6638 => x"27",
          6639 => x"61",
          6640 => x"70",
          6641 => x"0c",
          6642 => x"f5",
          6643 => x"39",
          6644 => x"80",
          6645 => x"84",
          6646 => x"ed",
          6647 => x"f8",
          6648 => x"2e",
          6649 => x"b4",
          6650 => x"11",
          6651 => x"05",
          6652 => x"ca",
          6653 => x"c8",
          6654 => x"fd",
          6655 => x"3d",
          6656 => x"53",
          6657 => x"51",
          6658 => x"3f",
          6659 => x"08",
          6660 => x"ac",
          6661 => x"dc",
          6662 => x"c9",
          6663 => x"79",
          6664 => x"8c",
          6665 => x"79",
          6666 => x"5b",
          6667 => x"61",
          6668 => x"eb",
          6669 => x"ff",
          6670 => x"ff",
          6671 => x"fe",
          6672 => x"81",
          6673 => x"80",
          6674 => x"38",
          6675 => x"fc",
          6676 => x"84",
          6677 => x"ec",
          6678 => x"f8",
          6679 => x"2e",
          6680 => x"b4",
          6681 => x"11",
          6682 => x"05",
          6683 => x"ce",
          6684 => x"c8",
          6685 => x"fc",
          6686 => x"f0",
          6687 => x"e4",
          6688 => x"5a",
          6689 => x"a8",
          6690 => x"33",
          6691 => x"5a",
          6692 => x"2e",
          6693 => x"55",
          6694 => x"33",
          6695 => x"81",
          6696 => x"fe",
          6697 => x"81",
          6698 => x"05",
          6699 => x"39",
          6700 => x"51",
          6701 => x"b4",
          6702 => x"11",
          6703 => x"05",
          6704 => x"fa",
          6705 => x"c8",
          6706 => x"38",
          6707 => x"33",
          6708 => x"2e",
          6709 => x"f3",
          6710 => x"80",
          6711 => x"f4",
          6712 => x"78",
          6713 => x"38",
          6714 => x"08",
          6715 => x"81",
          6716 => x"59",
          6717 => x"88",
          6718 => x"d4",
          6719 => x"39",
          6720 => x"33",
          6721 => x"2e",
          6722 => x"f3",
          6723 => x"9a",
          6724 => x"8a",
          6725 => x"80",
          6726 => x"81",
          6727 => x"44",
          6728 => x"f3",
          6729 => x"80",
          6730 => x"3d",
          6731 => x"53",
          6732 => x"51",
          6733 => x"3f",
          6734 => x"08",
          6735 => x"81",
          6736 => x"59",
          6737 => x"89",
          6738 => x"c8",
          6739 => x"cc",
          6740 => x"8d",
          6741 => x"80",
          6742 => x"81",
          6743 => x"43",
          6744 => x"f4",
          6745 => x"78",
          6746 => x"38",
          6747 => x"08",
          6748 => x"81",
          6749 => x"59",
          6750 => x"88",
          6751 => x"e0",
          6752 => x"39",
          6753 => x"33",
          6754 => x"2e",
          6755 => x"f3",
          6756 => x"88",
          6757 => x"f4",
          6758 => x"43",
          6759 => x"f8",
          6760 => x"84",
          6761 => x"ea",
          6762 => x"f8",
          6763 => x"2e",
          6764 => x"62",
          6765 => x"88",
          6766 => x"81",
          6767 => x"32",
          6768 => x"72",
          6769 => x"70",
          6770 => x"51",
          6771 => x"80",
          6772 => x"7a",
          6773 => x"38",
          6774 => x"f1",
          6775 => x"e2",
          6776 => x"55",
          6777 => x"53",
          6778 => x"51",
          6779 => x"81",
          6780 => x"fe",
          6781 => x"f9",
          6782 => x"3d",
          6783 => x"53",
          6784 => x"51",
          6785 => x"3f",
          6786 => x"08",
          6787 => x"b0",
          6788 => x"fe",
          6789 => x"ff",
          6790 => x"fe",
          6791 => x"81",
          6792 => x"80",
          6793 => x"63",
          6794 => x"cb",
          6795 => x"34",
          6796 => x"44",
          6797 => x"fc",
          6798 => x"84",
          6799 => x"e8",
          6800 => x"f8",
          6801 => x"38",
          6802 => x"63",
          6803 => x"52",
          6804 => x"51",
          6805 => x"3f",
          6806 => x"79",
          6807 => x"c3",
          6808 => x"79",
          6809 => x"ae",
          6810 => x"38",
          6811 => x"a0",
          6812 => x"fe",
          6813 => x"ff",
          6814 => x"fe",
          6815 => x"81",
          6816 => x"80",
          6817 => x"63",
          6818 => x"cb",
          6819 => x"34",
          6820 => x"44",
          6821 => x"81",
          6822 => x"fe",
          6823 => x"ff",
          6824 => x"3d",
          6825 => x"53",
          6826 => x"51",
          6827 => x"3f",
          6828 => x"08",
          6829 => x"88",
          6830 => x"fe",
          6831 => x"ff",
          6832 => x"fe",
          6833 => x"81",
          6834 => x"80",
          6835 => x"60",
          6836 => x"05",
          6837 => x"82",
          6838 => x"78",
          6839 => x"fe",
          6840 => x"ff",
          6841 => x"fe",
          6842 => x"81",
          6843 => x"df",
          6844 => x"39",
          6845 => x"54",
          6846 => x"c4",
          6847 => x"c9",
          6848 => x"52",
          6849 => x"e6",
          6850 => x"45",
          6851 => x"78",
          6852 => x"ac",
          6853 => x"26",
          6854 => x"82",
          6855 => x"39",
          6856 => x"f0",
          6857 => x"84",
          6858 => x"e9",
          6859 => x"f8",
          6860 => x"2e",
          6861 => x"59",
          6862 => x"22",
          6863 => x"05",
          6864 => x"41",
          6865 => x"81",
          6866 => x"fe",
          6867 => x"ff",
          6868 => x"3d",
          6869 => x"53",
          6870 => x"51",
          6871 => x"3f",
          6872 => x"08",
          6873 => x"d8",
          6874 => x"fe",
          6875 => x"ff",
          6876 => x"fe",
          6877 => x"81",
          6878 => x"80",
          6879 => x"60",
          6880 => x"59",
          6881 => x"41",
          6882 => x"f0",
          6883 => x"84",
          6884 => x"e8",
          6885 => x"f8",
          6886 => x"38",
          6887 => x"60",
          6888 => x"52",
          6889 => x"51",
          6890 => x"3f",
          6891 => x"79",
          6892 => x"ef",
          6893 => x"79",
          6894 => x"ae",
          6895 => x"38",
          6896 => x"9c",
          6897 => x"fe",
          6898 => x"ff",
          6899 => x"fe",
          6900 => x"81",
          6901 => x"80",
          6902 => x"60",
          6903 => x"59",
          6904 => x"41",
          6905 => x"81",
          6906 => x"fe",
          6907 => x"ff",
          6908 => x"3d",
          6909 => x"53",
          6910 => x"51",
          6911 => x"3f",
          6912 => x"08",
          6913 => x"b8",
          6914 => x"81",
          6915 => x"fe",
          6916 => x"63",
          6917 => x"b4",
          6918 => x"11",
          6919 => x"05",
          6920 => x"9a",
          6921 => x"c8",
          6922 => x"f5",
          6923 => x"52",
          6924 => x"51",
          6925 => x"3f",
          6926 => x"2d",
          6927 => x"08",
          6928 => x"fc",
          6929 => x"c8",
          6930 => x"f2",
          6931 => x"e2",
          6932 => x"ec",
          6933 => x"b0",
          6934 => x"89",
          6935 => x"ad",
          6936 => x"39",
          6937 => x"51",
          6938 => x"3f",
          6939 => x"a5",
          6940 => x"8e",
          6941 => x"39",
          6942 => x"33",
          6943 => x"2e",
          6944 => x"7d",
          6945 => x"78",
          6946 => x"d3",
          6947 => x"ff",
          6948 => x"fe",
          6949 => x"81",
          6950 => x"5c",
          6951 => x"82",
          6952 => x"7a",
          6953 => x"38",
          6954 => x"8c",
          6955 => x"39",
          6956 => x"b0",
          6957 => x"39",
          6958 => x"56",
          6959 => x"f2",
          6960 => x"53",
          6961 => x"52",
          6962 => x"b0",
          6963 => x"e2",
          6964 => x"39",
          6965 => x"52",
          6966 => x"b0",
          6967 => x"e1",
          6968 => x"39",
          6969 => x"f2",
          6970 => x"53",
          6971 => x"52",
          6972 => x"b0",
          6973 => x"e1",
          6974 => x"39",
          6975 => x"53",
          6976 => x"52",
          6977 => x"b0",
          6978 => x"e1",
          6979 => x"f3",
          6980 => x"f9",
          6981 => x"56",
          6982 => x"54",
          6983 => x"53",
          6984 => x"52",
          6985 => x"b0",
          6986 => x"8a",
          6987 => x"c8",
          6988 => x"c8",
          6989 => x"30",
          6990 => x"80",
          6991 => x"5b",
          6992 => x"7a",
          6993 => x"38",
          6994 => x"7a",
          6995 => x"80",
          6996 => x"81",
          6997 => x"ff",
          6998 => x"7a",
          6999 => x"7d",
          7000 => x"81",
          7001 => x"78",
          7002 => x"ff",
          7003 => x"06",
          7004 => x"81",
          7005 => x"fe",
          7006 => x"f2",
          7007 => x"3d",
          7008 => x"81",
          7009 => x"87",
          7010 => x"70",
          7011 => x"87",
          7012 => x"72",
          7013 => x"94",
          7014 => x"c8",
          7015 => x"75",
          7016 => x"87",
          7017 => x"73",
          7018 => x"80",
          7019 => x"f8",
          7020 => x"75",
          7021 => x"94",
          7022 => x"54",
          7023 => x"80",
          7024 => x"fe",
          7025 => x"81",
          7026 => x"90",
          7027 => x"55",
          7028 => x"80",
          7029 => x"fe",
          7030 => x"72",
          7031 => x"08",
          7032 => x"8c",
          7033 => x"87",
          7034 => x"0c",
          7035 => x"0b",
          7036 => x"94",
          7037 => x"0b",
          7038 => x"0c",
          7039 => x"81",
          7040 => x"fe",
          7041 => x"fe",
          7042 => x"81",
          7043 => x"fe",
          7044 => x"81",
          7045 => x"fe",
          7046 => x"81",
          7047 => x"fe",
          7048 => x"81",
          7049 => x"3f",
          7050 => x"80",
          7051 => x"ff",
          7052 => x"ff",
          7053 => x"00",
          7054 => x"ff",
          7055 => x"18",
          7056 => x"18",
          7057 => x"18",
          7058 => x"18",
          7059 => x"18",
          7060 => x"25",
          7061 => x"26",
          7062 => x"27",
          7063 => x"27",
          7064 => x"27",
          7065 => x"28",
          7066 => x"24",
          7067 => x"24",
          7068 => x"28",
          7069 => x"28",
          7070 => x"29",
          7071 => x"29",
          7072 => x"61",
          7073 => x"61",
          7074 => x"61",
          7075 => x"61",
          7076 => x"61",
          7077 => x"61",
          7078 => x"61",
          7079 => x"61",
          7080 => x"61",
          7081 => x"61",
          7082 => x"61",
          7083 => x"61",
          7084 => x"61",
          7085 => x"61",
          7086 => x"61",
          7087 => x"61",
          7088 => x"61",
          7089 => x"61",
          7090 => x"61",
          7091 => x"61",
          7092 => x"2f",
          7093 => x"25",
          7094 => x"64",
          7095 => x"3a",
          7096 => x"25",
          7097 => x"0a",
          7098 => x"43",
          7099 => x"6e",
          7100 => x"75",
          7101 => x"69",
          7102 => x"00",
          7103 => x"66",
          7104 => x"20",
          7105 => x"20",
          7106 => x"66",
          7107 => x"00",
          7108 => x"44",
          7109 => x"63",
          7110 => x"69",
          7111 => x"65",
          7112 => x"74",
          7113 => x"0a",
          7114 => x"20",
          7115 => x"20",
          7116 => x"41",
          7117 => x"28",
          7118 => x"58",
          7119 => x"38",
          7120 => x"0a",
          7121 => x"20",
          7122 => x"52",
          7123 => x"20",
          7124 => x"28",
          7125 => x"58",
          7126 => x"38",
          7127 => x"0a",
          7128 => x"20",
          7129 => x"53",
          7130 => x"52",
          7131 => x"28",
          7132 => x"58",
          7133 => x"38",
          7134 => x"0a",
          7135 => x"20",
          7136 => x"41",
          7137 => x"20",
          7138 => x"28",
          7139 => x"58",
          7140 => x"38",
          7141 => x"0a",
          7142 => x"20",
          7143 => x"4d",
          7144 => x"20",
          7145 => x"28",
          7146 => x"58",
          7147 => x"38",
          7148 => x"0a",
          7149 => x"20",
          7150 => x"20",
          7151 => x"44",
          7152 => x"28",
          7153 => x"69",
          7154 => x"20",
          7155 => x"32",
          7156 => x"0a",
          7157 => x"20",
          7158 => x"4d",
          7159 => x"20",
          7160 => x"28",
          7161 => x"65",
          7162 => x"20",
          7163 => x"32",
          7164 => x"0a",
          7165 => x"20",
          7166 => x"54",
          7167 => x"54",
          7168 => x"28",
          7169 => x"6e",
          7170 => x"73",
          7171 => x"32",
          7172 => x"0a",
          7173 => x"20",
          7174 => x"53",
          7175 => x"4e",
          7176 => x"55",
          7177 => x"00",
          7178 => x"20",
          7179 => x"20",
          7180 => x"0a",
          7181 => x"20",
          7182 => x"43",
          7183 => x"00",
          7184 => x"20",
          7185 => x"32",
          7186 => x"00",
          7187 => x"20",
          7188 => x"49",
          7189 => x"00",
          7190 => x"64",
          7191 => x"73",
          7192 => x"0a",
          7193 => x"20",
          7194 => x"55",
          7195 => x"73",
          7196 => x"56",
          7197 => x"6f",
          7198 => x"64",
          7199 => x"73",
          7200 => x"20",
          7201 => x"58",
          7202 => x"00",
          7203 => x"20",
          7204 => x"55",
          7205 => x"6d",
          7206 => x"20",
          7207 => x"72",
          7208 => x"64",
          7209 => x"73",
          7210 => x"20",
          7211 => x"58",
          7212 => x"00",
          7213 => x"20",
          7214 => x"61",
          7215 => x"53",
          7216 => x"74",
          7217 => x"64",
          7218 => x"73",
          7219 => x"20",
          7220 => x"20",
          7221 => x"58",
          7222 => x"00",
          7223 => x"73",
          7224 => x"00",
          7225 => x"20",
          7226 => x"55",
          7227 => x"20",
          7228 => x"20",
          7229 => x"20",
          7230 => x"20",
          7231 => x"20",
          7232 => x"20",
          7233 => x"58",
          7234 => x"00",
          7235 => x"20",
          7236 => x"73",
          7237 => x"20",
          7238 => x"63",
          7239 => x"72",
          7240 => x"20",
          7241 => x"20",
          7242 => x"20",
          7243 => x"25",
          7244 => x"4d",
          7245 => x"00",
          7246 => x"20",
          7247 => x"52",
          7248 => x"43",
          7249 => x"6b",
          7250 => x"65",
          7251 => x"20",
          7252 => x"20",
          7253 => x"20",
          7254 => x"25",
          7255 => x"4d",
          7256 => x"00",
          7257 => x"20",
          7258 => x"73",
          7259 => x"6e",
          7260 => x"44",
          7261 => x"20",
          7262 => x"63",
          7263 => x"72",
          7264 => x"20",
          7265 => x"25",
          7266 => x"4d",
          7267 => x"00",
          7268 => x"61",
          7269 => x"00",
          7270 => x"64",
          7271 => x"00",
          7272 => x"65",
          7273 => x"00",
          7274 => x"4f",
          7275 => x"4f",
          7276 => x"00",
          7277 => x"6b",
          7278 => x"6e",
          7279 => x"73",
          7280 => x"79",
          7281 => x"74",
          7282 => x"73",
          7283 => x"79",
          7284 => x"73",
          7285 => x"00",
          7286 => x"00",
          7287 => x"34",
          7288 => x"25",
          7289 => x"00",
          7290 => x"69",
          7291 => x"20",
          7292 => x"72",
          7293 => x"74",
          7294 => x"65",
          7295 => x"73",
          7296 => x"79",
          7297 => x"6c",
          7298 => x"6f",
          7299 => x"46",
          7300 => x"00",
          7301 => x"6e",
          7302 => x"20",
          7303 => x"6e",
          7304 => x"65",
          7305 => x"20",
          7306 => x"74",
          7307 => x"20",
          7308 => x"65",
          7309 => x"69",
          7310 => x"6c",
          7311 => x"2e",
          7312 => x"00",
          7313 => x"72",
          7314 => x"00",
          7315 => x"00",
          7316 => x"72",
          7317 => x"00",
          7318 => x"00",
          7319 => x"72",
          7320 => x"00",
          7321 => x"00",
          7322 => x"72",
          7323 => x"00",
          7324 => x"00",
          7325 => x"72",
          7326 => x"00",
          7327 => x"00",
          7328 => x"72",
          7329 => x"00",
          7330 => x"00",
          7331 => x"72",
          7332 => x"00",
          7333 => x"00",
          7334 => x"72",
          7335 => x"00",
          7336 => x"00",
          7337 => x"72",
          7338 => x"00",
          7339 => x"00",
          7340 => x"72",
          7341 => x"00",
          7342 => x"00",
          7343 => x"72",
          7344 => x"00",
          7345 => x"00",
          7346 => x"44",
          7347 => x"43",
          7348 => x"42",
          7349 => x"41",
          7350 => x"36",
          7351 => x"35",
          7352 => x"34",
          7353 => x"33",
          7354 => x"31",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"2b",
          7359 => x"3c",
          7360 => x"5b",
          7361 => x"00",
          7362 => x"54",
          7363 => x"54",
          7364 => x"00",
          7365 => x"90",
          7366 => x"4f",
          7367 => x"30",
          7368 => x"20",
          7369 => x"45",
          7370 => x"20",
          7371 => x"33",
          7372 => x"20",
          7373 => x"20",
          7374 => x"45",
          7375 => x"20",
          7376 => x"20",
          7377 => x"20",
          7378 => x"72",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"45",
          7383 => x"8f",
          7384 => x"45",
          7385 => x"8e",
          7386 => x"92",
          7387 => x"55",
          7388 => x"9a",
          7389 => x"9e",
          7390 => x"4f",
          7391 => x"a6",
          7392 => x"aa",
          7393 => x"ae",
          7394 => x"b2",
          7395 => x"b6",
          7396 => x"ba",
          7397 => x"be",
          7398 => x"c2",
          7399 => x"c6",
          7400 => x"ca",
          7401 => x"ce",
          7402 => x"d2",
          7403 => x"d6",
          7404 => x"da",
          7405 => x"de",
          7406 => x"e2",
          7407 => x"e6",
          7408 => x"ea",
          7409 => x"ee",
          7410 => x"f2",
          7411 => x"f6",
          7412 => x"fa",
          7413 => x"fe",
          7414 => x"2c",
          7415 => x"5d",
          7416 => x"2a",
          7417 => x"3f",
          7418 => x"00",
          7419 => x"00",
          7420 => x"00",
          7421 => x"02",
          7422 => x"00",
          7423 => x"00",
          7424 => x"00",
          7425 => x"00",
          7426 => x"00",
          7427 => x"6e",
          7428 => x"00",
          7429 => x"6f",
          7430 => x"00",
          7431 => x"6e",
          7432 => x"00",
          7433 => x"6f",
          7434 => x"00",
          7435 => x"78",
          7436 => x"00",
          7437 => x"6c",
          7438 => x"00",
          7439 => x"6f",
          7440 => x"00",
          7441 => x"69",
          7442 => x"00",
          7443 => x"75",
          7444 => x"00",
          7445 => x"62",
          7446 => x"68",
          7447 => x"77",
          7448 => x"64",
          7449 => x"65",
          7450 => x"64",
          7451 => x"65",
          7452 => x"6c",
          7453 => x"00",
          7454 => x"70",
          7455 => x"73",
          7456 => x"74",
          7457 => x"73",
          7458 => x"00",
          7459 => x"66",
          7460 => x"00",
          7461 => x"73",
          7462 => x"00",
          7463 => x"61",
          7464 => x"00",
          7465 => x"61",
          7466 => x"00",
          7467 => x"6c",
          7468 => x"00",
          7469 => x"73",
          7470 => x"72",
          7471 => x"0a",
          7472 => x"74",
          7473 => x"61",
          7474 => x"72",
          7475 => x"2e",
          7476 => x"00",
          7477 => x"73",
          7478 => x"6f",
          7479 => x"65",
          7480 => x"2e",
          7481 => x"00",
          7482 => x"20",
          7483 => x"65",
          7484 => x"75",
          7485 => x"0a",
          7486 => x"20",
          7487 => x"68",
          7488 => x"75",
          7489 => x"0a",
          7490 => x"76",
          7491 => x"64",
          7492 => x"6c",
          7493 => x"6d",
          7494 => x"00",
          7495 => x"63",
          7496 => x"20",
          7497 => x"69",
          7498 => x"0a",
          7499 => x"6c",
          7500 => x"6c",
          7501 => x"64",
          7502 => x"78",
          7503 => x"73",
          7504 => x"00",
          7505 => x"6c",
          7506 => x"61",
          7507 => x"65",
          7508 => x"76",
          7509 => x"64",
          7510 => x"00",
          7511 => x"20",
          7512 => x"77",
          7513 => x"65",
          7514 => x"6f",
          7515 => x"74",
          7516 => x"0a",
          7517 => x"69",
          7518 => x"6e",
          7519 => x"65",
          7520 => x"73",
          7521 => x"76",
          7522 => x"64",
          7523 => x"00",
          7524 => x"73",
          7525 => x"6f",
          7526 => x"6e",
          7527 => x"65",
          7528 => x"00",
          7529 => x"20",
          7530 => x"70",
          7531 => x"62",
          7532 => x"66",
          7533 => x"73",
          7534 => x"65",
          7535 => x"6f",
          7536 => x"20",
          7537 => x"64",
          7538 => x"2e",
          7539 => x"00",
          7540 => x"72",
          7541 => x"20",
          7542 => x"72",
          7543 => x"2e",
          7544 => x"00",
          7545 => x"6d",
          7546 => x"74",
          7547 => x"70",
          7548 => x"74",
          7549 => x"20",
          7550 => x"63",
          7551 => x"65",
          7552 => x"00",
          7553 => x"6c",
          7554 => x"73",
          7555 => x"63",
          7556 => x"2e",
          7557 => x"00",
          7558 => x"73",
          7559 => x"69",
          7560 => x"6e",
          7561 => x"65",
          7562 => x"79",
          7563 => x"00",
          7564 => x"6f",
          7565 => x"6e",
          7566 => x"70",
          7567 => x"66",
          7568 => x"73",
          7569 => x"00",
          7570 => x"72",
          7571 => x"74",
          7572 => x"20",
          7573 => x"6f",
          7574 => x"63",
          7575 => x"00",
          7576 => x"63",
          7577 => x"73",
          7578 => x"00",
          7579 => x"6b",
          7580 => x"6e",
          7581 => x"72",
          7582 => x"0a",
          7583 => x"6c",
          7584 => x"79",
          7585 => x"20",
          7586 => x"61",
          7587 => x"6c",
          7588 => x"79",
          7589 => x"2f",
          7590 => x"2e",
          7591 => x"00",
          7592 => x"61",
          7593 => x"00",
          7594 => x"38",
          7595 => x"00",
          7596 => x"20",
          7597 => x"34",
          7598 => x"00",
          7599 => x"20",
          7600 => x"20",
          7601 => x"00",
          7602 => x"32",
          7603 => x"00",
          7604 => x"00",
          7605 => x"00",
          7606 => x"0a",
          7607 => x"53",
          7608 => x"2a",
          7609 => x"20",
          7610 => x"00",
          7611 => x"2f",
          7612 => x"32",
          7613 => x"00",
          7614 => x"2e",
          7615 => x"00",
          7616 => x"50",
          7617 => x"72",
          7618 => x"25",
          7619 => x"29",
          7620 => x"20",
          7621 => x"2a",
          7622 => x"00",
          7623 => x"55",
          7624 => x"74",
          7625 => x"75",
          7626 => x"48",
          7627 => x"6c",
          7628 => x"00",
          7629 => x"6d",
          7630 => x"69",
          7631 => x"72",
          7632 => x"74",
          7633 => x"00",
          7634 => x"32",
          7635 => x"74",
          7636 => x"75",
          7637 => x"00",
          7638 => x"43",
          7639 => x"52",
          7640 => x"6e",
          7641 => x"72",
          7642 => x"0a",
          7643 => x"43",
          7644 => x"57",
          7645 => x"6e",
          7646 => x"72",
          7647 => x"0a",
          7648 => x"52",
          7649 => x"52",
          7650 => x"6e",
          7651 => x"72",
          7652 => x"0a",
          7653 => x"52",
          7654 => x"54",
          7655 => x"6e",
          7656 => x"72",
          7657 => x"0a",
          7658 => x"52",
          7659 => x"52",
          7660 => x"6e",
          7661 => x"72",
          7662 => x"0a",
          7663 => x"52",
          7664 => x"54",
          7665 => x"6e",
          7666 => x"72",
          7667 => x"0a",
          7668 => x"74",
          7669 => x"67",
          7670 => x"20",
          7671 => x"65",
          7672 => x"2e",
          7673 => x"00",
          7674 => x"61",
          7675 => x"6e",
          7676 => x"69",
          7677 => x"2e",
          7678 => x"00",
          7679 => x"74",
          7680 => x"65",
          7681 => x"61",
          7682 => x"00",
          7683 => x"00",
          7684 => x"69",
          7685 => x"20",
          7686 => x"69",
          7687 => x"69",
          7688 => x"73",
          7689 => x"64",
          7690 => x"72",
          7691 => x"2c",
          7692 => x"65",
          7693 => x"20",
          7694 => x"74",
          7695 => x"6e",
          7696 => x"6c",
          7697 => x"00",
          7698 => x"00",
          7699 => x"65",
          7700 => x"6e",
          7701 => x"2e",
          7702 => x"00",
          7703 => x"70",
          7704 => x"67",
          7705 => x"00",
          7706 => x"6d",
          7707 => x"69",
          7708 => x"2e",
          7709 => x"00",
          7710 => x"38",
          7711 => x"25",
          7712 => x"29",
          7713 => x"30",
          7714 => x"28",
          7715 => x"78",
          7716 => x"00",
          7717 => x"6d",
          7718 => x"65",
          7719 => x"79",
          7720 => x"00",
          7721 => x"6f",
          7722 => x"65",
          7723 => x"0a",
          7724 => x"38",
          7725 => x"30",
          7726 => x"00",
          7727 => x"3f",
          7728 => x"00",
          7729 => x"38",
          7730 => x"30",
          7731 => x"00",
          7732 => x"38",
          7733 => x"30",
          7734 => x"00",
          7735 => x"65",
          7736 => x"69",
          7737 => x"63",
          7738 => x"20",
          7739 => x"30",
          7740 => x"2e",
          7741 => x"00",
          7742 => x"6c",
          7743 => x"67",
          7744 => x"64",
          7745 => x"20",
          7746 => x"78",
          7747 => x"2e",
          7748 => x"00",
          7749 => x"6c",
          7750 => x"65",
          7751 => x"6e",
          7752 => x"63",
          7753 => x"20",
          7754 => x"29",
          7755 => x"00",
          7756 => x"73",
          7757 => x"74",
          7758 => x"20",
          7759 => x"6c",
          7760 => x"74",
          7761 => x"2e",
          7762 => x"00",
          7763 => x"6c",
          7764 => x"65",
          7765 => x"74",
          7766 => x"2e",
          7767 => x"00",
          7768 => x"55",
          7769 => x"6e",
          7770 => x"3a",
          7771 => x"5c",
          7772 => x"25",
          7773 => x"00",
          7774 => x"3a",
          7775 => x"5c",
          7776 => x"00",
          7777 => x"3a",
          7778 => x"00",
          7779 => x"64",
          7780 => x"6d",
          7781 => x"64",
          7782 => x"00",
          7783 => x"6e",
          7784 => x"67",
          7785 => x"0a",
          7786 => x"61",
          7787 => x"6e",
          7788 => x"6e",
          7789 => x"72",
          7790 => x"73",
          7791 => x"0a",
          7792 => x"00",
          7793 => x"00",
          7794 => x"7f",
          7795 => x"00",
          7796 => x"7f",
          7797 => x"00",
          7798 => x"7f",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"ff",
          7803 => x"00",
          7804 => x"00",
          7805 => x"78",
          7806 => x"00",
          7807 => x"e1",
          7808 => x"e1",
          7809 => x"e1",
          7810 => x"00",
          7811 => x"01",
          7812 => x"01",
          7813 => x"10",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"7a",
          7819 => x"7a",
          7820 => x"7a",
          7821 => x"7a",
          7822 => x"71",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"71",
          7847 => x"00",
          7848 => x"71",
          7849 => x"00",
          7850 => x"71",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"74",
          7855 => x"01",
          7856 => x"00",
          7857 => x"00",
          7858 => x"74",
          7859 => x"01",
          7860 => x"00",
          7861 => x"00",
          7862 => x"74",
          7863 => x"03",
          7864 => x"00",
          7865 => x"00",
          7866 => x"74",
          7867 => x"03",
          7868 => x"00",
          7869 => x"00",
          7870 => x"74",
          7871 => x"03",
          7872 => x"00",
          7873 => x"00",
          7874 => x"74",
          7875 => x"04",
          7876 => x"00",
          7877 => x"00",
          7878 => x"74",
          7879 => x"04",
          7880 => x"00",
          7881 => x"00",
          7882 => x"74",
          7883 => x"04",
          7884 => x"00",
          7885 => x"00",
          7886 => x"74",
          7887 => x"04",
          7888 => x"00",
          7889 => x"00",
          7890 => x"74",
          7891 => x"04",
          7892 => x"00",
          7893 => x"00",
          7894 => x"74",
          7895 => x"04",
          7896 => x"00",
          7897 => x"00",
          7898 => x"74",
          7899 => x"04",
          7900 => x"00",
          7901 => x"00",
          7902 => x"74",
          7903 => x"05",
          7904 => x"00",
          7905 => x"00",
          7906 => x"74",
          7907 => x"05",
          7908 => x"00",
          7909 => x"00",
          7910 => x"74",
          7911 => x"05",
          7912 => x"00",
          7913 => x"00",
          7914 => x"74",
          7915 => x"05",
          7916 => x"00",
          7917 => x"00",
          7918 => x"74",
          7919 => x"07",
          7920 => x"00",
          7921 => x"00",
          7922 => x"74",
          7923 => x"07",
          7924 => x"00",
          7925 => x"00",
          7926 => x"74",
          7927 => x"08",
          7928 => x"00",
          7929 => x"00",
          7930 => x"74",
          7931 => x"08",
          7932 => x"00",
          7933 => x"00",
          7934 => x"74",
          7935 => x"08",
          7936 => x"00",
          7937 => x"00",
          7938 => x"74",
          7939 => x"08",
          7940 => x"00",
          7941 => x"00",
          7942 => x"74",
          7943 => x"09",
          7944 => x"00",
          7945 => x"00",
          7946 => x"74",
          7947 => x"09",
          7948 => x"00",
          7949 => x"00",
          7950 => x"74",
          7951 => x"09",
          7952 => x"00",
          7953 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"d8",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"81",
           386 => x"a3",
           387 => x"f8",
           388 => x"80",
           389 => x"f8",
           390 => x"87",
           391 => x"d4",
           392 => x"90",
           393 => x"d4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"81",
           399 => x"83",
           400 => x"81",
           401 => x"bc",
           402 => x"f8",
           403 => x"80",
           404 => x"f8",
           405 => x"a0",
           406 => x"d4",
           407 => x"90",
           408 => x"d4",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"81",
           414 => x"83",
           415 => x"81",
           416 => x"bf",
           417 => x"f8",
           418 => x"80",
           419 => x"f8",
           420 => x"c8",
           421 => x"d4",
           422 => x"90",
           423 => x"d4",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"81",
           429 => x"83",
           430 => x"81",
           431 => x"bc",
           432 => x"f8",
           433 => x"80",
           434 => x"f8",
           435 => x"8c",
           436 => x"d4",
           437 => x"90",
           438 => x"d4",
           439 => x"2d",
           440 => x"08",
           441 => x"04",
           442 => x"0c",
           443 => x"81",
           444 => x"83",
           445 => x"81",
           446 => x"a0",
           447 => x"f8",
           448 => x"80",
           449 => x"f8",
           450 => x"e1",
           451 => x"d4",
           452 => x"90",
           453 => x"d4",
           454 => x"82",
           455 => x"d4",
           456 => x"90",
           457 => x"d4",
           458 => x"f3",
           459 => x"d4",
           460 => x"90",
           461 => x"d4",
           462 => x"e7",
           463 => x"d4",
           464 => x"90",
           465 => x"d4",
           466 => x"e4",
           467 => x"d4",
           468 => x"90",
           469 => x"d4",
           470 => x"82",
           471 => x"d4",
           472 => x"90",
           473 => x"d4",
           474 => x"e2",
           475 => x"d4",
           476 => x"90",
           477 => x"d4",
           478 => x"d5",
           479 => x"d4",
           480 => x"90",
           481 => x"d4",
           482 => x"a1",
           483 => x"d4",
           484 => x"90",
           485 => x"d4",
           486 => x"c0",
           487 => x"d4",
           488 => x"90",
           489 => x"d4",
           490 => x"df",
           491 => x"d4",
           492 => x"90",
           493 => x"d4",
           494 => x"c9",
           495 => x"d4",
           496 => x"90",
           497 => x"d4",
           498 => x"af",
           499 => x"d4",
           500 => x"90",
           501 => x"d4",
           502 => x"9d",
           503 => x"d4",
           504 => x"90",
           505 => x"d4",
           506 => x"e3",
           507 => x"d4",
           508 => x"90",
           509 => x"d4",
           510 => x"9d",
           511 => x"d4",
           512 => x"90",
           513 => x"d4",
           514 => x"9e",
           515 => x"d4",
           516 => x"90",
           517 => x"d4",
           518 => x"d3",
           519 => x"d4",
           520 => x"90",
           521 => x"d4",
           522 => x"ac",
           523 => x"d4",
           524 => x"90",
           525 => x"d4",
           526 => x"d7",
           527 => x"d4",
           528 => x"90",
           529 => x"d4",
           530 => x"ba",
           531 => x"d4",
           532 => x"90",
           533 => x"d4",
           534 => x"8f",
           535 => x"d4",
           536 => x"90",
           537 => x"d4",
           538 => x"99",
           539 => x"d4",
           540 => x"90",
           541 => x"d4",
           542 => x"db",
           543 => x"d4",
           544 => x"90",
           545 => x"d4",
           546 => x"a1",
           547 => x"d4",
           548 => x"90",
           549 => x"d4",
           550 => x"c7",
           551 => x"d4",
           552 => x"90",
           553 => x"d4",
           554 => x"fc",
           555 => x"d4",
           556 => x"90",
           557 => x"d4",
           558 => x"e8",
           559 => x"d4",
           560 => x"90",
           561 => x"d4",
           562 => x"dc",
           563 => x"d4",
           564 => x"90",
           565 => x"d4",
           566 => x"c6",
           567 => x"d4",
           568 => x"90",
           569 => x"d4",
           570 => x"aa",
           571 => x"d4",
           572 => x"90",
           573 => x"d4",
           574 => x"2d",
           575 => x"08",
           576 => x"04",
           577 => x"0c",
           578 => x"81",
           579 => x"83",
           580 => x"81",
           581 => x"a2",
           582 => x"f8",
           583 => x"80",
           584 => x"f8",
           585 => x"c2",
           586 => x"f8",
           587 => x"80",
           588 => x"04",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"04",
           598 => x"81",
           599 => x"83",
           600 => x"05",
           601 => x"10",
           602 => x"72",
           603 => x"51",
           604 => x"72",
           605 => x"06",
           606 => x"72",
           607 => x"10",
           608 => x"10",
           609 => x"ed",
           610 => x"53",
           611 => x"f8",
           612 => x"90",
           613 => x"38",
           614 => x"84",
           615 => x"0b",
           616 => x"8f",
           617 => x"51",
           618 => x"04",
           619 => x"d4",
           620 => x"f8",
           621 => x"3d",
           622 => x"81",
           623 => x"8c",
           624 => x"81",
           625 => x"88",
           626 => x"83",
           627 => x"f8",
           628 => x"81",
           629 => x"54",
           630 => x"81",
           631 => x"04",
           632 => x"08",
           633 => x"d4",
           634 => x"0d",
           635 => x"f8",
           636 => x"05",
           637 => x"f8",
           638 => x"05",
           639 => x"a1",
           640 => x"c8",
           641 => x"f8",
           642 => x"85",
           643 => x"f8",
           644 => x"81",
           645 => x"02",
           646 => x"0c",
           647 => x"80",
           648 => x"d4",
           649 => x"0c",
           650 => x"08",
           651 => x"80",
           652 => x"81",
           653 => x"88",
           654 => x"81",
           655 => x"88",
           656 => x"0b",
           657 => x"08",
           658 => x"81",
           659 => x"fc",
           660 => x"38",
           661 => x"f8",
           662 => x"05",
           663 => x"d4",
           664 => x"08",
           665 => x"08",
           666 => x"81",
           667 => x"8c",
           668 => x"25",
           669 => x"f8",
           670 => x"05",
           671 => x"f8",
           672 => x"05",
           673 => x"81",
           674 => x"f0",
           675 => x"f8",
           676 => x"05",
           677 => x"81",
           678 => x"d4",
           679 => x"0c",
           680 => x"08",
           681 => x"81",
           682 => x"fc",
           683 => x"53",
           684 => x"08",
           685 => x"52",
           686 => x"08",
           687 => x"51",
           688 => x"81",
           689 => x"70",
           690 => x"08",
           691 => x"54",
           692 => x"08",
           693 => x"80",
           694 => x"81",
           695 => x"f8",
           696 => x"81",
           697 => x"f8",
           698 => x"f8",
           699 => x"05",
           700 => x"f8",
           701 => x"89",
           702 => x"f8",
           703 => x"81",
           704 => x"02",
           705 => x"0c",
           706 => x"80",
           707 => x"d4",
           708 => x"0c",
           709 => x"08",
           710 => x"80",
           711 => x"81",
           712 => x"88",
           713 => x"81",
           714 => x"88",
           715 => x"0b",
           716 => x"08",
           717 => x"81",
           718 => x"8c",
           719 => x"25",
           720 => x"f8",
           721 => x"05",
           722 => x"f8",
           723 => x"05",
           724 => x"81",
           725 => x"8c",
           726 => x"81",
           727 => x"88",
           728 => x"bd",
           729 => x"c8",
           730 => x"f8",
           731 => x"05",
           732 => x"f8",
           733 => x"05",
           734 => x"90",
           735 => x"d4",
           736 => x"08",
           737 => x"d4",
           738 => x"0c",
           739 => x"08",
           740 => x"70",
           741 => x"0c",
           742 => x"0d",
           743 => x"0c",
           744 => x"d4",
           745 => x"f8",
           746 => x"3d",
           747 => x"81",
           748 => x"fc",
           749 => x"0b",
           750 => x"08",
           751 => x"81",
           752 => x"8c",
           753 => x"f8",
           754 => x"05",
           755 => x"38",
           756 => x"08",
           757 => x"80",
           758 => x"80",
           759 => x"d4",
           760 => x"08",
           761 => x"81",
           762 => x"8c",
           763 => x"81",
           764 => x"8c",
           765 => x"f8",
           766 => x"05",
           767 => x"f8",
           768 => x"05",
           769 => x"39",
           770 => x"08",
           771 => x"80",
           772 => x"38",
           773 => x"08",
           774 => x"81",
           775 => x"88",
           776 => x"ad",
           777 => x"d4",
           778 => x"08",
           779 => x"08",
           780 => x"31",
           781 => x"08",
           782 => x"81",
           783 => x"f8",
           784 => x"f8",
           785 => x"05",
           786 => x"f8",
           787 => x"05",
           788 => x"d4",
           789 => x"08",
           790 => x"f8",
           791 => x"05",
           792 => x"d4",
           793 => x"08",
           794 => x"f8",
           795 => x"05",
           796 => x"39",
           797 => x"08",
           798 => x"80",
           799 => x"81",
           800 => x"88",
           801 => x"81",
           802 => x"f4",
           803 => x"91",
           804 => x"d4",
           805 => x"08",
           806 => x"d4",
           807 => x"0c",
           808 => x"d4",
           809 => x"08",
           810 => x"0c",
           811 => x"81",
           812 => x"04",
           813 => x"76",
           814 => x"55",
           815 => x"8f",
           816 => x"38",
           817 => x"83",
           818 => x"80",
           819 => x"ff",
           820 => x"ff",
           821 => x"72",
           822 => x"54",
           823 => x"81",
           824 => x"ff",
           825 => x"ff",
           826 => x"06",
           827 => x"81",
           828 => x"86",
           829 => x"74",
           830 => x"84",
           831 => x"71",
           832 => x"53",
           833 => x"84",
           834 => x"71",
           835 => x"53",
           836 => x"84",
           837 => x"71",
           838 => x"53",
           839 => x"84",
           840 => x"71",
           841 => x"53",
           842 => x"52",
           843 => x"c9",
           844 => x"27",
           845 => x"70",
           846 => x"08",
           847 => x"05",
           848 => x"12",
           849 => x"26",
           850 => x"54",
           851 => x"fc",
           852 => x"79",
           853 => x"05",
           854 => x"57",
           855 => x"83",
           856 => x"38",
           857 => x"51",
           858 => x"a4",
           859 => x"52",
           860 => x"93",
           861 => x"70",
           862 => x"34",
           863 => x"71",
           864 => x"81",
           865 => x"74",
           866 => x"0c",
           867 => x"04",
           868 => x"2b",
           869 => x"71",
           870 => x"51",
           871 => x"72",
           872 => x"72",
           873 => x"05",
           874 => x"71",
           875 => x"53",
           876 => x"70",
           877 => x"0c",
           878 => x"84",
           879 => x"f0",
           880 => x"8f",
           881 => x"83",
           882 => x"38",
           883 => x"84",
           884 => x"fc",
           885 => x"83",
           886 => x"70",
           887 => x"39",
           888 => x"76",
           889 => x"73",
           890 => x"54",
           891 => x"70",
           892 => x"71",
           893 => x"09",
           894 => x"fd",
           895 => x"70",
           896 => x"81",
           897 => x"51",
           898 => x"70",
           899 => x"14",
           900 => x"84",
           901 => x"70",
           902 => x"70",
           903 => x"ff",
           904 => x"f8",
           905 => x"80",
           906 => x"53",
           907 => x"80",
           908 => x"73",
           909 => x"81",
           910 => x"51",
           911 => x"81",
           912 => x"70",
           913 => x"81",
           914 => x"86",
           915 => x"fd",
           916 => x"70",
           917 => x"53",
           918 => x"b8",
           919 => x"08",
           920 => x"fb",
           921 => x"06",
           922 => x"82",
           923 => x"51",
           924 => x"70",
           925 => x"13",
           926 => x"09",
           927 => x"ff",
           928 => x"f8",
           929 => x"80",
           930 => x"52",
           931 => x"2e",
           932 => x"52",
           933 => x"70",
           934 => x"38",
           935 => x"33",
           936 => x"f8",
           937 => x"31",
           938 => x"0c",
           939 => x"04",
           940 => x"78",
           941 => x"54",
           942 => x"72",
           943 => x"d9",
           944 => x"07",
           945 => x"70",
           946 => x"d6",
           947 => x"53",
           948 => x"b1",
           949 => x"74",
           950 => x"74",
           951 => x"81",
           952 => x"72",
           953 => x"89",
           954 => x"ff",
           955 => x"80",
           956 => x"38",
           957 => x"15",
           958 => x"55",
           959 => x"2e",
           960 => x"d1",
           961 => x"74",
           962 => x"70",
           963 => x"75",
           964 => x"71",
           965 => x"52",
           966 => x"f8",
           967 => x"3d",
           968 => x"74",
           969 => x"73",
           970 => x"71",
           971 => x"2e",
           972 => x"76",
           973 => x"95",
           974 => x"53",
           975 => x"b1",
           976 => x"70",
           977 => x"fd",
           978 => x"70",
           979 => x"81",
           980 => x"51",
           981 => x"38",
           982 => x"17",
           983 => x"73",
           984 => x"74",
           985 => x"2e",
           986 => x"76",
           987 => x"dd",
           988 => x"81",
           989 => x"88",
           990 => x"fe",
           991 => x"52",
           992 => x"88",
           993 => x"86",
           994 => x"c8",
           995 => x"06",
           996 => x"14",
           997 => x"80",
           998 => x"71",
           999 => x"0c",
          1000 => x"04",
          1001 => x"77",
          1002 => x"53",
          1003 => x"80",
          1004 => x"38",
          1005 => x"70",
          1006 => x"81",
          1007 => x"81",
          1008 => x"39",
          1009 => x"39",
          1010 => x"80",
          1011 => x"81",
          1012 => x"55",
          1013 => x"2e",
          1014 => x"55",
          1015 => x"84",
          1016 => x"38",
          1017 => x"06",
          1018 => x"2e",
          1019 => x"88",
          1020 => x"70",
          1021 => x"34",
          1022 => x"71",
          1023 => x"f8",
          1024 => x"3d",
          1025 => x"3d",
          1026 => x"72",
          1027 => x"91",
          1028 => x"fc",
          1029 => x"51",
          1030 => x"81",
          1031 => x"85",
          1032 => x"83",
          1033 => x"72",
          1034 => x"0c",
          1035 => x"04",
          1036 => x"76",
          1037 => x"ff",
          1038 => x"81",
          1039 => x"26",
          1040 => x"83",
          1041 => x"05",
          1042 => x"70",
          1043 => x"8a",
          1044 => x"33",
          1045 => x"70",
          1046 => x"fe",
          1047 => x"33",
          1048 => x"70",
          1049 => x"f2",
          1050 => x"33",
          1051 => x"70",
          1052 => x"e6",
          1053 => x"22",
          1054 => x"74",
          1055 => x"80",
          1056 => x"13",
          1057 => x"52",
          1058 => x"26",
          1059 => x"81",
          1060 => x"98",
          1061 => x"22",
          1062 => x"bc",
          1063 => x"33",
          1064 => x"b8",
          1065 => x"33",
          1066 => x"b4",
          1067 => x"33",
          1068 => x"b0",
          1069 => x"33",
          1070 => x"ac",
          1071 => x"33",
          1072 => x"a8",
          1073 => x"c0",
          1074 => x"73",
          1075 => x"a0",
          1076 => x"87",
          1077 => x"0c",
          1078 => x"81",
          1079 => x"86",
          1080 => x"f3",
          1081 => x"5b",
          1082 => x"9c",
          1083 => x"0c",
          1084 => x"bc",
          1085 => x"7b",
          1086 => x"98",
          1087 => x"79",
          1088 => x"87",
          1089 => x"08",
          1090 => x"1c",
          1091 => x"98",
          1092 => x"79",
          1093 => x"87",
          1094 => x"08",
          1095 => x"1c",
          1096 => x"98",
          1097 => x"79",
          1098 => x"87",
          1099 => x"08",
          1100 => x"1c",
          1101 => x"98",
          1102 => x"79",
          1103 => x"80",
          1104 => x"83",
          1105 => x"59",
          1106 => x"ff",
          1107 => x"1b",
          1108 => x"1b",
          1109 => x"1b",
          1110 => x"1b",
          1111 => x"1b",
          1112 => x"83",
          1113 => x"52",
          1114 => x"51",
          1115 => x"8f",
          1116 => x"ff",
          1117 => x"8f",
          1118 => x"30",
          1119 => x"51",
          1120 => x"0b",
          1121 => x"c0",
          1122 => x"0d",
          1123 => x"0d",
          1124 => x"81",
          1125 => x"70",
          1126 => x"57",
          1127 => x"c0",
          1128 => x"74",
          1129 => x"38",
          1130 => x"94",
          1131 => x"70",
          1132 => x"81",
          1133 => x"52",
          1134 => x"8c",
          1135 => x"2a",
          1136 => x"51",
          1137 => x"38",
          1138 => x"70",
          1139 => x"51",
          1140 => x"8d",
          1141 => x"2a",
          1142 => x"51",
          1143 => x"be",
          1144 => x"ff",
          1145 => x"c0",
          1146 => x"70",
          1147 => x"38",
          1148 => x"90",
          1149 => x"0c",
          1150 => x"c8",
          1151 => x"0d",
          1152 => x"0d",
          1153 => x"33",
          1154 => x"f3",
          1155 => x"81",
          1156 => x"55",
          1157 => x"94",
          1158 => x"80",
          1159 => x"87",
          1160 => x"51",
          1161 => x"96",
          1162 => x"06",
          1163 => x"70",
          1164 => x"38",
          1165 => x"70",
          1166 => x"51",
          1167 => x"72",
          1168 => x"81",
          1169 => x"70",
          1170 => x"38",
          1171 => x"70",
          1172 => x"51",
          1173 => x"38",
          1174 => x"06",
          1175 => x"94",
          1176 => x"80",
          1177 => x"87",
          1178 => x"52",
          1179 => x"87",
          1180 => x"f9",
          1181 => x"54",
          1182 => x"70",
          1183 => x"53",
          1184 => x"77",
          1185 => x"38",
          1186 => x"06",
          1187 => x"0b",
          1188 => x"33",
          1189 => x"06",
          1190 => x"58",
          1191 => x"84",
          1192 => x"2e",
          1193 => x"c0",
          1194 => x"70",
          1195 => x"2a",
          1196 => x"53",
          1197 => x"80",
          1198 => x"71",
          1199 => x"81",
          1200 => x"70",
          1201 => x"81",
          1202 => x"06",
          1203 => x"80",
          1204 => x"71",
          1205 => x"81",
          1206 => x"70",
          1207 => x"74",
          1208 => x"51",
          1209 => x"80",
          1210 => x"2e",
          1211 => x"c0",
          1212 => x"77",
          1213 => x"17",
          1214 => x"81",
          1215 => x"53",
          1216 => x"84",
          1217 => x"f8",
          1218 => x"3d",
          1219 => x"3d",
          1220 => x"81",
          1221 => x"70",
          1222 => x"54",
          1223 => x"94",
          1224 => x"80",
          1225 => x"87",
          1226 => x"51",
          1227 => x"82",
          1228 => x"06",
          1229 => x"70",
          1230 => x"38",
          1231 => x"06",
          1232 => x"94",
          1233 => x"80",
          1234 => x"87",
          1235 => x"52",
          1236 => x"81",
          1237 => x"f8",
          1238 => x"84",
          1239 => x"fe",
          1240 => x"0b",
          1241 => x"33",
          1242 => x"06",
          1243 => x"c0",
          1244 => x"70",
          1245 => x"38",
          1246 => x"94",
          1247 => x"70",
          1248 => x"81",
          1249 => x"51",
          1250 => x"80",
          1251 => x"72",
          1252 => x"51",
          1253 => x"80",
          1254 => x"2e",
          1255 => x"c0",
          1256 => x"71",
          1257 => x"2b",
          1258 => x"51",
          1259 => x"81",
          1260 => x"84",
          1261 => x"ff",
          1262 => x"c0",
          1263 => x"70",
          1264 => x"06",
          1265 => x"80",
          1266 => x"38",
          1267 => x"a4",
          1268 => x"c4",
          1269 => x"9e",
          1270 => x"f3",
          1271 => x"c0",
          1272 => x"81",
          1273 => x"87",
          1274 => x"08",
          1275 => x"0c",
          1276 => x"9c",
          1277 => x"d4",
          1278 => x"9e",
          1279 => x"f3",
          1280 => x"c0",
          1281 => x"81",
          1282 => x"87",
          1283 => x"08",
          1284 => x"0c",
          1285 => x"b4",
          1286 => x"e4",
          1287 => x"9e",
          1288 => x"f3",
          1289 => x"c0",
          1290 => x"81",
          1291 => x"87",
          1292 => x"08",
          1293 => x"0c",
          1294 => x"c4",
          1295 => x"f4",
          1296 => x"9e",
          1297 => x"70",
          1298 => x"23",
          1299 => x"84",
          1300 => x"fc",
          1301 => x"9e",
          1302 => x"f4",
          1303 => x"c0",
          1304 => x"81",
          1305 => x"81",
          1306 => x"88",
          1307 => x"87",
          1308 => x"08",
          1309 => x"0a",
          1310 => x"52",
          1311 => x"83",
          1312 => x"71",
          1313 => x"34",
          1314 => x"c0",
          1315 => x"70",
          1316 => x"06",
          1317 => x"70",
          1318 => x"38",
          1319 => x"81",
          1320 => x"80",
          1321 => x"9e",
          1322 => x"90",
          1323 => x"51",
          1324 => x"80",
          1325 => x"81",
          1326 => x"f4",
          1327 => x"0b",
          1328 => x"90",
          1329 => x"80",
          1330 => x"52",
          1331 => x"2e",
          1332 => x"52",
          1333 => x"8c",
          1334 => x"87",
          1335 => x"08",
          1336 => x"80",
          1337 => x"52",
          1338 => x"83",
          1339 => x"71",
          1340 => x"34",
          1341 => x"c0",
          1342 => x"70",
          1343 => x"06",
          1344 => x"70",
          1345 => x"38",
          1346 => x"81",
          1347 => x"80",
          1348 => x"9e",
          1349 => x"84",
          1350 => x"51",
          1351 => x"80",
          1352 => x"81",
          1353 => x"f4",
          1354 => x"0b",
          1355 => x"90",
          1356 => x"80",
          1357 => x"52",
          1358 => x"2e",
          1359 => x"52",
          1360 => x"90",
          1361 => x"87",
          1362 => x"08",
          1363 => x"80",
          1364 => x"52",
          1365 => x"83",
          1366 => x"71",
          1367 => x"34",
          1368 => x"c0",
          1369 => x"70",
          1370 => x"06",
          1371 => x"70",
          1372 => x"38",
          1373 => x"81",
          1374 => x"80",
          1375 => x"9e",
          1376 => x"a0",
          1377 => x"52",
          1378 => x"2e",
          1379 => x"52",
          1380 => x"93",
          1381 => x"9e",
          1382 => x"98",
          1383 => x"8a",
          1384 => x"51",
          1385 => x"94",
          1386 => x"87",
          1387 => x"08",
          1388 => x"06",
          1389 => x"70",
          1390 => x"38",
          1391 => x"81",
          1392 => x"87",
          1393 => x"08",
          1394 => x"06",
          1395 => x"51",
          1396 => x"81",
          1397 => x"80",
          1398 => x"9e",
          1399 => x"88",
          1400 => x"52",
          1401 => x"83",
          1402 => x"71",
          1403 => x"34",
          1404 => x"90",
          1405 => x"06",
          1406 => x"81",
          1407 => x"83",
          1408 => x"fb",
          1409 => x"dd",
          1410 => x"da",
          1411 => x"88",
          1412 => x"80",
          1413 => x"81",
          1414 => x"89",
          1415 => x"de",
          1416 => x"c2",
          1417 => x"8a",
          1418 => x"80",
          1419 => x"81",
          1420 => x"81",
          1421 => x"11",
          1422 => x"de",
          1423 => x"8a",
          1424 => x"8f",
          1425 => x"80",
          1426 => x"81",
          1427 => x"81",
          1428 => x"11",
          1429 => x"de",
          1430 => x"ee",
          1431 => x"8c",
          1432 => x"80",
          1433 => x"81",
          1434 => x"81",
          1435 => x"11",
          1436 => x"de",
          1437 => x"d2",
          1438 => x"8d",
          1439 => x"80",
          1440 => x"81",
          1441 => x"81",
          1442 => x"11",
          1443 => x"de",
          1444 => x"b6",
          1445 => x"8e",
          1446 => x"80",
          1447 => x"81",
          1448 => x"81",
          1449 => x"11",
          1450 => x"df",
          1451 => x"9a",
          1452 => x"93",
          1453 => x"80",
          1454 => x"81",
          1455 => x"52",
          1456 => x"51",
          1457 => x"81",
          1458 => x"54",
          1459 => x"8d",
          1460 => x"98",
          1461 => x"df",
          1462 => x"ee",
          1463 => x"95",
          1464 => x"80",
          1465 => x"81",
          1466 => x"52",
          1467 => x"51",
          1468 => x"81",
          1469 => x"54",
          1470 => x"88",
          1471 => x"94",
          1472 => x"3f",
          1473 => x"33",
          1474 => x"2e",
          1475 => x"e0",
          1476 => x"d2",
          1477 => x"90",
          1478 => x"80",
          1479 => x"81",
          1480 => x"87",
          1481 => x"f4",
          1482 => x"73",
          1483 => x"38",
          1484 => x"51",
          1485 => x"81",
          1486 => x"54",
          1487 => x"88",
          1488 => x"cc",
          1489 => x"3f",
          1490 => x"51",
          1491 => x"81",
          1492 => x"52",
          1493 => x"51",
          1494 => x"81",
          1495 => x"52",
          1496 => x"51",
          1497 => x"81",
          1498 => x"52",
          1499 => x"51",
          1500 => x"81",
          1501 => x"86",
          1502 => x"f3",
          1503 => x"81",
          1504 => x"8c",
          1505 => x"f3",
          1506 => x"bd",
          1507 => x"75",
          1508 => x"3f",
          1509 => x"08",
          1510 => x"29",
          1511 => x"54",
          1512 => x"c8",
          1513 => x"e2",
          1514 => x"9e",
          1515 => x"8f",
          1516 => x"80",
          1517 => x"81",
          1518 => x"56",
          1519 => x"52",
          1520 => x"e9",
          1521 => x"c8",
          1522 => x"c0",
          1523 => x"31",
          1524 => x"f8",
          1525 => x"81",
          1526 => x"8b",
          1527 => x"f4",
          1528 => x"73",
          1529 => x"38",
          1530 => x"08",
          1531 => x"c0",
          1532 => x"e3",
          1533 => x"f8",
          1534 => x"84",
          1535 => x"71",
          1536 => x"81",
          1537 => x"52",
          1538 => x"51",
          1539 => x"81",
          1540 => x"85",
          1541 => x"3d",
          1542 => x"3d",
          1543 => x"05",
          1544 => x"52",
          1545 => x"aa",
          1546 => x"29",
          1547 => x"05",
          1548 => x"04",
          1549 => x"51",
          1550 => x"e3",
          1551 => x"39",
          1552 => x"51",
          1553 => x"e3",
          1554 => x"39",
          1555 => x"51",
          1556 => x"e3",
          1557 => x"8e",
          1558 => x"0d",
          1559 => x"80",
          1560 => x"0b",
          1561 => x"84",
          1562 => x"f4",
          1563 => x"c0",
          1564 => x"04",
          1565 => x"81",
          1566 => x"89",
          1567 => x"88",
          1568 => x"d8",
          1569 => x"d8",
          1570 => x"52",
          1571 => x"70",
          1572 => x"26",
          1573 => x"81",
          1574 => x"71",
          1575 => x"f8",
          1576 => x"3d",
          1577 => x"3d",
          1578 => x"84",
          1579 => x"12",
          1580 => x"94",
          1581 => x"16",
          1582 => x"54",
          1583 => x"70",
          1584 => x"38",
          1585 => x"14",
          1586 => x"81",
          1587 => x"76",
          1588 => x"0c",
          1589 => x"75",
          1590 => x"72",
          1591 => x"71",
          1592 => x"70",
          1593 => x"70",
          1594 => x"73",
          1595 => x"74",
          1596 => x"70",
          1597 => x"70",
          1598 => x"8c",
          1599 => x"0c",
          1600 => x"0c",
          1601 => x"0c",
          1602 => x"c8",
          1603 => x"0d",
          1604 => x"0d",
          1605 => x"08",
          1606 => x"56",
          1607 => x"08",
          1608 => x"81",
          1609 => x"84",
          1610 => x"13",
          1611 => x"73",
          1612 => x"06",
          1613 => x"13",
          1614 => x"13",
          1615 => x"13",
          1616 => x"15",
          1617 => x"9f",
          1618 => x"0c",
          1619 => x"08",
          1620 => x"81",
          1621 => x"94",
          1622 => x"81",
          1623 => x"90",
          1624 => x"94",
          1625 => x"73",
          1626 => x"09",
          1627 => x"38",
          1628 => x"70",
          1629 => x"70",
          1630 => x"81",
          1631 => x"84",
          1632 => x"84",
          1633 => x"14",
          1634 => x"08",
          1635 => x"0c",
          1636 => x"0c",
          1637 => x"88",
          1638 => x"88",
          1639 => x"8c",
          1640 => x"81",
          1641 => x"86",
          1642 => x"f9",
          1643 => x"70",
          1644 => x"80",
          1645 => x"38",
          1646 => x"06",
          1647 => x"08",
          1648 => x"08",
          1649 => x"38",
          1650 => x"77",
          1651 => x"38",
          1652 => x"56",
          1653 => x"ff",
          1654 => x"80",
          1655 => x"52",
          1656 => x"3f",
          1657 => x"08",
          1658 => x"08",
          1659 => x"f8",
          1660 => x"80",
          1661 => x"c8",
          1662 => x"30",
          1663 => x"80",
          1664 => x"53",
          1665 => x"54",
          1666 => x"72",
          1667 => x"81",
          1668 => x"38",
          1669 => x"52",
          1670 => x"c8",
          1671 => x"81",
          1672 => x"0c",
          1673 => x"c8",
          1674 => x"0c",
          1675 => x"08",
          1676 => x"82",
          1677 => x"75",
          1678 => x"38",
          1679 => x"53",
          1680 => x"13",
          1681 => x"0c",
          1682 => x"0c",
          1683 => x"0c",
          1684 => x"76",
          1685 => x"53",
          1686 => x"b5",
          1687 => x"81",
          1688 => x"51",
          1689 => x"81",
          1690 => x"54",
          1691 => x"c8",
          1692 => x"0d",
          1693 => x"0d",
          1694 => x"80",
          1695 => x"f0",
          1696 => x"8d",
          1697 => x"0d",
          1698 => x"0d",
          1699 => x"33",
          1700 => x"2e",
          1701 => x"85",
          1702 => x"ed",
          1703 => x"e4",
          1704 => x"80",
          1705 => x"72",
          1706 => x"f8",
          1707 => x"05",
          1708 => x"0c",
          1709 => x"f8",
          1710 => x"71",
          1711 => x"38",
          1712 => x"2d",
          1713 => x"04",
          1714 => x"02",
          1715 => x"81",
          1716 => x"76",
          1717 => x"0c",
          1718 => x"ad",
          1719 => x"f8",
          1720 => x"3d",
          1721 => x"3d",
          1722 => x"73",
          1723 => x"ff",
          1724 => x"71",
          1725 => x"38",
          1726 => x"06",
          1727 => x"54",
          1728 => x"e7",
          1729 => x"0d",
          1730 => x"0d",
          1731 => x"dc",
          1732 => x"f8",
          1733 => x"54",
          1734 => x"81",
          1735 => x"53",
          1736 => x"8e",
          1737 => x"ff",
          1738 => x"14",
          1739 => x"3f",
          1740 => x"81",
          1741 => x"86",
          1742 => x"ec",
          1743 => x"68",
          1744 => x"70",
          1745 => x"33",
          1746 => x"2e",
          1747 => x"75",
          1748 => x"81",
          1749 => x"38",
          1750 => x"70",
          1751 => x"33",
          1752 => x"75",
          1753 => x"81",
          1754 => x"81",
          1755 => x"75",
          1756 => x"81",
          1757 => x"82",
          1758 => x"81",
          1759 => x"56",
          1760 => x"09",
          1761 => x"38",
          1762 => x"71",
          1763 => x"81",
          1764 => x"59",
          1765 => x"9d",
          1766 => x"53",
          1767 => x"95",
          1768 => x"29",
          1769 => x"76",
          1770 => x"79",
          1771 => x"5b",
          1772 => x"e5",
          1773 => x"ec",
          1774 => x"70",
          1775 => x"25",
          1776 => x"32",
          1777 => x"72",
          1778 => x"73",
          1779 => x"58",
          1780 => x"73",
          1781 => x"38",
          1782 => x"79",
          1783 => x"5b",
          1784 => x"75",
          1785 => x"de",
          1786 => x"80",
          1787 => x"89",
          1788 => x"70",
          1789 => x"55",
          1790 => x"cf",
          1791 => x"38",
          1792 => x"24",
          1793 => x"80",
          1794 => x"8e",
          1795 => x"c3",
          1796 => x"73",
          1797 => x"81",
          1798 => x"99",
          1799 => x"c4",
          1800 => x"38",
          1801 => x"73",
          1802 => x"81",
          1803 => x"80",
          1804 => x"38",
          1805 => x"2e",
          1806 => x"f9",
          1807 => x"d8",
          1808 => x"38",
          1809 => x"77",
          1810 => x"08",
          1811 => x"80",
          1812 => x"55",
          1813 => x"8d",
          1814 => x"70",
          1815 => x"51",
          1816 => x"f5",
          1817 => x"2a",
          1818 => x"74",
          1819 => x"53",
          1820 => x"8f",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"80",
          1824 => x"73",
          1825 => x"3f",
          1826 => x"56",
          1827 => x"27",
          1828 => x"a0",
          1829 => x"3f",
          1830 => x"84",
          1831 => x"33",
          1832 => x"93",
          1833 => x"95",
          1834 => x"91",
          1835 => x"8d",
          1836 => x"89",
          1837 => x"fb",
          1838 => x"86",
          1839 => x"2a",
          1840 => x"51",
          1841 => x"2e",
          1842 => x"84",
          1843 => x"86",
          1844 => x"78",
          1845 => x"08",
          1846 => x"32",
          1847 => x"72",
          1848 => x"51",
          1849 => x"74",
          1850 => x"38",
          1851 => x"88",
          1852 => x"7a",
          1853 => x"55",
          1854 => x"3d",
          1855 => x"52",
          1856 => x"dc",
          1857 => x"c8",
          1858 => x"06",
          1859 => x"52",
          1860 => x"3f",
          1861 => x"08",
          1862 => x"27",
          1863 => x"14",
          1864 => x"f8",
          1865 => x"87",
          1866 => x"81",
          1867 => x"b0",
          1868 => x"7d",
          1869 => x"5f",
          1870 => x"75",
          1871 => x"07",
          1872 => x"54",
          1873 => x"26",
          1874 => x"ff",
          1875 => x"84",
          1876 => x"06",
          1877 => x"80",
          1878 => x"96",
          1879 => x"e0",
          1880 => x"73",
          1881 => x"57",
          1882 => x"06",
          1883 => x"54",
          1884 => x"a0",
          1885 => x"2a",
          1886 => x"54",
          1887 => x"38",
          1888 => x"76",
          1889 => x"38",
          1890 => x"fd",
          1891 => x"06",
          1892 => x"38",
          1893 => x"56",
          1894 => x"26",
          1895 => x"3d",
          1896 => x"05",
          1897 => x"ff",
          1898 => x"53",
          1899 => x"d9",
          1900 => x"38",
          1901 => x"56",
          1902 => x"27",
          1903 => x"a0",
          1904 => x"3f",
          1905 => x"3d",
          1906 => x"3d",
          1907 => x"70",
          1908 => x"52",
          1909 => x"73",
          1910 => x"3f",
          1911 => x"04",
          1912 => x"74",
          1913 => x"0c",
          1914 => x"05",
          1915 => x"fa",
          1916 => x"f8",
          1917 => x"80",
          1918 => x"0b",
          1919 => x"0c",
          1920 => x"04",
          1921 => x"81",
          1922 => x"76",
          1923 => x"0c",
          1924 => x"05",
          1925 => x"53",
          1926 => x"72",
          1927 => x"0c",
          1928 => x"04",
          1929 => x"77",
          1930 => x"e0",
          1931 => x"54",
          1932 => x"54",
          1933 => x"80",
          1934 => x"f8",
          1935 => x"71",
          1936 => x"c8",
          1937 => x"06",
          1938 => x"2e",
          1939 => x"72",
          1940 => x"38",
          1941 => x"70",
          1942 => x"25",
          1943 => x"73",
          1944 => x"38",
          1945 => x"86",
          1946 => x"54",
          1947 => x"73",
          1948 => x"ff",
          1949 => x"72",
          1950 => x"74",
          1951 => x"72",
          1952 => x"54",
          1953 => x"81",
          1954 => x"39",
          1955 => x"80",
          1956 => x"51",
          1957 => x"81",
          1958 => x"f8",
          1959 => x"3d",
          1960 => x"3d",
          1961 => x"e0",
          1962 => x"f8",
          1963 => x"53",
          1964 => x"fe",
          1965 => x"81",
          1966 => x"84",
          1967 => x"f8",
          1968 => x"7c",
          1969 => x"70",
          1970 => x"75",
          1971 => x"55",
          1972 => x"2e",
          1973 => x"87",
          1974 => x"76",
          1975 => x"73",
          1976 => x"81",
          1977 => x"81",
          1978 => x"77",
          1979 => x"70",
          1980 => x"58",
          1981 => x"09",
          1982 => x"c2",
          1983 => x"81",
          1984 => x"75",
          1985 => x"55",
          1986 => x"e2",
          1987 => x"90",
          1988 => x"f8",
          1989 => x"8f",
          1990 => x"81",
          1991 => x"75",
          1992 => x"55",
          1993 => x"81",
          1994 => x"27",
          1995 => x"d0",
          1996 => x"55",
          1997 => x"73",
          1998 => x"80",
          1999 => x"14",
          2000 => x"72",
          2001 => x"e0",
          2002 => x"80",
          2003 => x"39",
          2004 => x"55",
          2005 => x"80",
          2006 => x"e0",
          2007 => x"38",
          2008 => x"81",
          2009 => x"53",
          2010 => x"81",
          2011 => x"53",
          2012 => x"8e",
          2013 => x"70",
          2014 => x"55",
          2015 => x"27",
          2016 => x"77",
          2017 => x"74",
          2018 => x"76",
          2019 => x"77",
          2020 => x"70",
          2021 => x"55",
          2022 => x"77",
          2023 => x"38",
          2024 => x"74",
          2025 => x"55",
          2026 => x"c8",
          2027 => x"0d",
          2028 => x"0d",
          2029 => x"56",
          2030 => x"0c",
          2031 => x"70",
          2032 => x"73",
          2033 => x"81",
          2034 => x"81",
          2035 => x"ed",
          2036 => x"2e",
          2037 => x"8e",
          2038 => x"08",
          2039 => x"76",
          2040 => x"56",
          2041 => x"b0",
          2042 => x"06",
          2043 => x"75",
          2044 => x"76",
          2045 => x"70",
          2046 => x"73",
          2047 => x"8b",
          2048 => x"73",
          2049 => x"85",
          2050 => x"82",
          2051 => x"76",
          2052 => x"70",
          2053 => x"ac",
          2054 => x"a0",
          2055 => x"fa",
          2056 => x"53",
          2057 => x"57",
          2058 => x"98",
          2059 => x"39",
          2060 => x"80",
          2061 => x"26",
          2062 => x"86",
          2063 => x"80",
          2064 => x"57",
          2065 => x"74",
          2066 => x"38",
          2067 => x"27",
          2068 => x"14",
          2069 => x"06",
          2070 => x"14",
          2071 => x"06",
          2072 => x"74",
          2073 => x"f9",
          2074 => x"ff",
          2075 => x"89",
          2076 => x"38",
          2077 => x"c5",
          2078 => x"29",
          2079 => x"81",
          2080 => x"76",
          2081 => x"56",
          2082 => x"ba",
          2083 => x"2e",
          2084 => x"30",
          2085 => x"0c",
          2086 => x"81",
          2087 => x"8a",
          2088 => x"fd",
          2089 => x"98",
          2090 => x"2c",
          2091 => x"70",
          2092 => x"10",
          2093 => x"2b",
          2094 => x"54",
          2095 => x"0b",
          2096 => x"12",
          2097 => x"71",
          2098 => x"38",
          2099 => x"11",
          2100 => x"84",
          2101 => x"33",
          2102 => x"52",
          2103 => x"2e",
          2104 => x"83",
          2105 => x"72",
          2106 => x"0c",
          2107 => x"04",
          2108 => x"78",
          2109 => x"9f",
          2110 => x"33",
          2111 => x"71",
          2112 => x"38",
          2113 => x"81",
          2114 => x"f2",
          2115 => x"51",
          2116 => x"72",
          2117 => x"52",
          2118 => x"71",
          2119 => x"52",
          2120 => x"51",
          2121 => x"73",
          2122 => x"3d",
          2123 => x"3d",
          2124 => x"84",
          2125 => x"33",
          2126 => x"bb",
          2127 => x"f5",
          2128 => x"84",
          2129 => x"bc",
          2130 => x"51",
          2131 => x"58",
          2132 => x"2e",
          2133 => x"51",
          2134 => x"81",
          2135 => x"70",
          2136 => x"f4",
          2137 => x"19",
          2138 => x"56",
          2139 => x"3f",
          2140 => x"08",
          2141 => x"f5",
          2142 => x"84",
          2143 => x"bc",
          2144 => x"51",
          2145 => x"80",
          2146 => x"75",
          2147 => x"74",
          2148 => x"3f",
          2149 => x"33",
          2150 => x"74",
          2151 => x"34",
          2152 => x"06",
          2153 => x"27",
          2154 => x"0b",
          2155 => x"34",
          2156 => x"b6",
          2157 => x"90",
          2158 => x"80",
          2159 => x"81",
          2160 => x"55",
          2161 => x"8c",
          2162 => x"54",
          2163 => x"52",
          2164 => x"c8",
          2165 => x"f5",
          2166 => x"8a",
          2167 => x"9e",
          2168 => x"90",
          2169 => x"cb",
          2170 => x"3d",
          2171 => x"3d",
          2172 => x"80",
          2173 => x"90",
          2174 => x"d2",
          2175 => x"f8",
          2176 => x"d1",
          2177 => x"90",
          2178 => x"f8",
          2179 => x"70",
          2180 => x"fa",
          2181 => x"f8",
          2182 => x"2e",
          2183 => x"51",
          2184 => x"81",
          2185 => x"55",
          2186 => x"f8",
          2187 => x"9c",
          2188 => x"c8",
          2189 => x"70",
          2190 => x"80",
          2191 => x"53",
          2192 => x"17",
          2193 => x"52",
          2194 => x"3f",
          2195 => x"09",
          2196 => x"b1",
          2197 => x"0d",
          2198 => x"0d",
          2199 => x"ad",
          2200 => x"5a",
          2201 => x"58",
          2202 => x"f5",
          2203 => x"80",
          2204 => x"81",
          2205 => x"81",
          2206 => x"0b",
          2207 => x"08",
          2208 => x"f8",
          2209 => x"70",
          2210 => x"f9",
          2211 => x"f8",
          2212 => x"2e",
          2213 => x"51",
          2214 => x"81",
          2215 => x"81",
          2216 => x"80",
          2217 => x"c8",
          2218 => x"38",
          2219 => x"08",
          2220 => x"17",
          2221 => x"74",
          2222 => x"70",
          2223 => x"07",
          2224 => x"55",
          2225 => x"2e",
          2226 => x"ff",
          2227 => x"f5",
          2228 => x"11",
          2229 => x"80",
          2230 => x"81",
          2231 => x"80",
          2232 => x"81",
          2233 => x"ef",
          2234 => x"77",
          2235 => x"06",
          2236 => x"52",
          2237 => x"e8",
          2238 => x"d6",
          2239 => x"3d",
          2240 => x"f8",
          2241 => x"34",
          2242 => x"81",
          2243 => x"a9",
          2244 => x"f6",
          2245 => x"7e",
          2246 => x"72",
          2247 => x"5a",
          2248 => x"2e",
          2249 => x"a2",
          2250 => x"78",
          2251 => x"76",
          2252 => x"81",
          2253 => x"70",
          2254 => x"58",
          2255 => x"2e",
          2256 => x"86",
          2257 => x"26",
          2258 => x"54",
          2259 => x"81",
          2260 => x"70",
          2261 => x"d5",
          2262 => x"f8",
          2263 => x"79",
          2264 => x"51",
          2265 => x"81",
          2266 => x"80",
          2267 => x"15",
          2268 => x"81",
          2269 => x"74",
          2270 => x"38",
          2271 => x"ee",
          2272 => x"81",
          2273 => x"3d",
          2274 => x"f8",
          2275 => x"af",
          2276 => x"c8",
          2277 => x"99",
          2278 => x"78",
          2279 => x"fd",
          2280 => x"f8",
          2281 => x"ff",
          2282 => x"85",
          2283 => x"91",
          2284 => x"70",
          2285 => x"51",
          2286 => x"27",
          2287 => x"80",
          2288 => x"f8",
          2289 => x"3d",
          2290 => x"3d",
          2291 => x"08",
          2292 => x"81",
          2293 => x"5f",
          2294 => x"af",
          2295 => x"f5",
          2296 => x"81",
          2297 => x"81",
          2298 => x"f5",
          2299 => x"73",
          2300 => x"a8",
          2301 => x"3f",
          2302 => x"08",
          2303 => x"0c",
          2304 => x"08",
          2305 => x"fe",
          2306 => x"81",
          2307 => x"52",
          2308 => x"08",
          2309 => x"3f",
          2310 => x"08",
          2311 => x"38",
          2312 => x"51",
          2313 => x"80",
          2314 => x"f5",
          2315 => x"80",
          2316 => x"3d",
          2317 => x"80",
          2318 => x"81",
          2319 => x"56",
          2320 => x"08",
          2321 => x"81",
          2322 => x"38",
          2323 => x"08",
          2324 => x"3f",
          2325 => x"08",
          2326 => x"81",
          2327 => x"25",
          2328 => x"f8",
          2329 => x"05",
          2330 => x"55",
          2331 => x"80",
          2332 => x"ff",
          2333 => x"51",
          2334 => x"74",
          2335 => x"81",
          2336 => x"38",
          2337 => x"0b",
          2338 => x"34",
          2339 => x"dd",
          2340 => x"f8",
          2341 => x"2b",
          2342 => x"51",
          2343 => x"2e",
          2344 => x"81",
          2345 => x"f8",
          2346 => x"98",
          2347 => x"2c",
          2348 => x"33",
          2349 => x"70",
          2350 => x"98",
          2351 => x"84",
          2352 => x"c4",
          2353 => x"15",
          2354 => x"51",
          2355 => x"59",
          2356 => x"58",
          2357 => x"78",
          2358 => x"38",
          2359 => x"b4",
          2360 => x"80",
          2361 => x"ff",
          2362 => x"98",
          2363 => x"80",
          2364 => x"ce",
          2365 => x"74",
          2366 => x"f7",
          2367 => x"f8",
          2368 => x"ff",
          2369 => x"80",
          2370 => x"74",
          2371 => x"34",
          2372 => x"39",
          2373 => x"0a",
          2374 => x"0a",
          2375 => x"2c",
          2376 => x"06",
          2377 => x"73",
          2378 => x"38",
          2379 => x"52",
          2380 => x"ef",
          2381 => x"c8",
          2382 => x"06",
          2383 => x"38",
          2384 => x"56",
          2385 => x"80",
          2386 => x"1c",
          2387 => x"f8",
          2388 => x"98",
          2389 => x"2c",
          2390 => x"33",
          2391 => x"70",
          2392 => x"10",
          2393 => x"2b",
          2394 => x"11",
          2395 => x"51",
          2396 => x"51",
          2397 => x"2e",
          2398 => x"fe",
          2399 => x"e4",
          2400 => x"7d",
          2401 => x"81",
          2402 => x"80",
          2403 => x"e8",
          2404 => x"75",
          2405 => x"34",
          2406 => x"e8",
          2407 => x"3d",
          2408 => x"0c",
          2409 => x"8b",
          2410 => x"38",
          2411 => x"81",
          2412 => x"54",
          2413 => x"81",
          2414 => x"54",
          2415 => x"fd",
          2416 => x"f8",
          2417 => x"73",
          2418 => x"38",
          2419 => x"70",
          2420 => x"55",
          2421 => x"9e",
          2422 => x"54",
          2423 => x"15",
          2424 => x"80",
          2425 => x"ff",
          2426 => x"98",
          2427 => x"f4",
          2428 => x"55",
          2429 => x"f8",
          2430 => x"11",
          2431 => x"81",
          2432 => x"73",
          2433 => x"3d",
          2434 => x"81",
          2435 => x"54",
          2436 => x"89",
          2437 => x"54",
          2438 => x"f0",
          2439 => x"f4",
          2440 => x"80",
          2441 => x"ff",
          2442 => x"98",
          2443 => x"f0",
          2444 => x"56",
          2445 => x"25",
          2446 => x"1a",
          2447 => x"54",
          2448 => x"74",
          2449 => x"29",
          2450 => x"05",
          2451 => x"81",
          2452 => x"56",
          2453 => x"75",
          2454 => x"81",
          2455 => x"70",
          2456 => x"98",
          2457 => x"f0",
          2458 => x"56",
          2459 => x"25",
          2460 => x"88",
          2461 => x"3f",
          2462 => x"0a",
          2463 => x"0a",
          2464 => x"2c",
          2465 => x"33",
          2466 => x"73",
          2467 => x"38",
          2468 => x"81",
          2469 => x"70",
          2470 => x"55",
          2471 => x"2e",
          2472 => x"81",
          2473 => x"ff",
          2474 => x"81",
          2475 => x"ff",
          2476 => x"81",
          2477 => x"88",
          2478 => x"3f",
          2479 => x"33",
          2480 => x"70",
          2481 => x"f8",
          2482 => x"51",
          2483 => x"74",
          2484 => x"74",
          2485 => x"14",
          2486 => x"73",
          2487 => x"a9",
          2488 => x"80",
          2489 => x"80",
          2490 => x"98",
          2491 => x"f0",
          2492 => x"55",
          2493 => x"db",
          2494 => x"e7",
          2495 => x"f8",
          2496 => x"98",
          2497 => x"2c",
          2498 => x"33",
          2499 => x"57",
          2500 => x"fa",
          2501 => x"51",
          2502 => x"74",
          2503 => x"29",
          2504 => x"05",
          2505 => x"81",
          2506 => x"58",
          2507 => x"75",
          2508 => x"fa",
          2509 => x"f8",
          2510 => x"05",
          2511 => x"34",
          2512 => x"c5",
          2513 => x"f0",
          2514 => x"f7",
          2515 => x"f8",
          2516 => x"ff",
          2517 => x"98",
          2518 => x"f0",
          2519 => x"80",
          2520 => x"38",
          2521 => x"52",
          2522 => x"c2",
          2523 => x"39",
          2524 => x"84",
          2525 => x"f8",
          2526 => x"73",
          2527 => x"8c",
          2528 => x"e6",
          2529 => x"f8",
          2530 => x"05",
          2531 => x"f8",
          2532 => x"81",
          2533 => x"e3",
          2534 => x"f4",
          2535 => x"f0",
          2536 => x"73",
          2537 => x"e4",
          2538 => x"54",
          2539 => x"f0",
          2540 => x"2b",
          2541 => x"75",
          2542 => x"56",
          2543 => x"74",
          2544 => x"74",
          2545 => x"14",
          2546 => x"73",
          2547 => x"b9",
          2548 => x"80",
          2549 => x"80",
          2550 => x"98",
          2551 => x"f0",
          2552 => x"55",
          2553 => x"db",
          2554 => x"e5",
          2555 => x"f8",
          2556 => x"98",
          2557 => x"2c",
          2558 => x"33",
          2559 => x"57",
          2560 => x"f9",
          2561 => x"51",
          2562 => x"74",
          2563 => x"29",
          2564 => x"05",
          2565 => x"81",
          2566 => x"58",
          2567 => x"75",
          2568 => x"f8",
          2569 => x"f8",
          2570 => x"81",
          2571 => x"f8",
          2572 => x"56",
          2573 => x"27",
          2574 => x"81",
          2575 => x"81",
          2576 => x"74",
          2577 => x"52",
          2578 => x"3f",
          2579 => x"33",
          2580 => x"06",
          2581 => x"33",
          2582 => x"75",
          2583 => x"38",
          2584 => x"7a",
          2585 => x"f5",
          2586 => x"74",
          2587 => x"38",
          2588 => x"db",
          2589 => x"c8",
          2590 => x"f0",
          2591 => x"c8",
          2592 => x"06",
          2593 => x"74",
          2594 => x"c8",
          2595 => x"5b",
          2596 => x"7a",
          2597 => x"f4",
          2598 => x"11",
          2599 => x"74",
          2600 => x"38",
          2601 => x"a7",
          2602 => x"c8",
          2603 => x"f0",
          2604 => x"c8",
          2605 => x"06",
          2606 => x"74",
          2607 => x"c7",
          2608 => x"1b",
          2609 => x"39",
          2610 => x"74",
          2611 => x"bc",
          2612 => x"ca",
          2613 => x"e2",
          2614 => x"2e",
          2615 => x"93",
          2616 => x"bc",
          2617 => x"80",
          2618 => x"74",
          2619 => x"3f",
          2620 => x"7a",
          2621 => x"f4",
          2622 => x"11",
          2623 => x"74",
          2624 => x"38",
          2625 => x"c7",
          2626 => x"c8",
          2627 => x"f0",
          2628 => x"c8",
          2629 => x"06",
          2630 => x"74",
          2631 => x"c7",
          2632 => x"1b",
          2633 => x"ff",
          2634 => x"39",
          2635 => x"74",
          2636 => x"d8",
          2637 => x"ca",
          2638 => x"f8",
          2639 => x"f8",
          2640 => x"f8",
          2641 => x"ff",
          2642 => x"53",
          2643 => x"51",
          2644 => x"81",
          2645 => x"81",
          2646 => x"52",
          2647 => x"90",
          2648 => x"39",
          2649 => x"33",
          2650 => x"06",
          2651 => x"33",
          2652 => x"74",
          2653 => x"94",
          2654 => x"54",
          2655 => x"f4",
          2656 => x"70",
          2657 => x"e2",
          2658 => x"80",
          2659 => x"f4",
          2660 => x"80",
          2661 => x"38",
          2662 => x"ed",
          2663 => x"f4",
          2664 => x"54",
          2665 => x"f4",
          2666 => x"39",
          2667 => x"f8",
          2668 => x"0b",
          2669 => x"34",
          2670 => x"c8",
          2671 => x"0d",
          2672 => x"0d",
          2673 => x"33",
          2674 => x"70",
          2675 => x"38",
          2676 => x"11",
          2677 => x"81",
          2678 => x"83",
          2679 => x"fc",
          2680 => x"9b",
          2681 => x"84",
          2682 => x"33",
          2683 => x"51",
          2684 => x"80",
          2685 => x"84",
          2686 => x"92",
          2687 => x"51",
          2688 => x"80",
          2689 => x"81",
          2690 => x"72",
          2691 => x"92",
          2692 => x"81",
          2693 => x"0b",
          2694 => x"8c",
          2695 => x"71",
          2696 => x"06",
          2697 => x"80",
          2698 => x"87",
          2699 => x"08",
          2700 => x"38",
          2701 => x"80",
          2702 => x"71",
          2703 => x"c0",
          2704 => x"51",
          2705 => x"87",
          2706 => x"f5",
          2707 => x"81",
          2708 => x"33",
          2709 => x"f8",
          2710 => x"3d",
          2711 => x"3d",
          2712 => x"64",
          2713 => x"bf",
          2714 => x"40",
          2715 => x"74",
          2716 => x"cd",
          2717 => x"c8",
          2718 => x"7a",
          2719 => x"81",
          2720 => x"72",
          2721 => x"87",
          2722 => x"11",
          2723 => x"8c",
          2724 => x"92",
          2725 => x"5a",
          2726 => x"58",
          2727 => x"c0",
          2728 => x"76",
          2729 => x"76",
          2730 => x"70",
          2731 => x"81",
          2732 => x"54",
          2733 => x"8e",
          2734 => x"52",
          2735 => x"81",
          2736 => x"81",
          2737 => x"74",
          2738 => x"53",
          2739 => x"83",
          2740 => x"78",
          2741 => x"8f",
          2742 => x"2e",
          2743 => x"c0",
          2744 => x"52",
          2745 => x"87",
          2746 => x"08",
          2747 => x"2e",
          2748 => x"84",
          2749 => x"38",
          2750 => x"87",
          2751 => x"15",
          2752 => x"70",
          2753 => x"52",
          2754 => x"ff",
          2755 => x"39",
          2756 => x"81",
          2757 => x"ff",
          2758 => x"57",
          2759 => x"90",
          2760 => x"80",
          2761 => x"71",
          2762 => x"78",
          2763 => x"38",
          2764 => x"80",
          2765 => x"80",
          2766 => x"81",
          2767 => x"72",
          2768 => x"0c",
          2769 => x"04",
          2770 => x"60",
          2771 => x"8c",
          2772 => x"33",
          2773 => x"5b",
          2774 => x"74",
          2775 => x"e1",
          2776 => x"c8",
          2777 => x"79",
          2778 => x"78",
          2779 => x"06",
          2780 => x"77",
          2781 => x"87",
          2782 => x"11",
          2783 => x"8c",
          2784 => x"92",
          2785 => x"59",
          2786 => x"85",
          2787 => x"98",
          2788 => x"7d",
          2789 => x"0c",
          2790 => x"08",
          2791 => x"70",
          2792 => x"53",
          2793 => x"2e",
          2794 => x"70",
          2795 => x"33",
          2796 => x"18",
          2797 => x"2a",
          2798 => x"51",
          2799 => x"2e",
          2800 => x"c0",
          2801 => x"52",
          2802 => x"87",
          2803 => x"08",
          2804 => x"2e",
          2805 => x"84",
          2806 => x"38",
          2807 => x"87",
          2808 => x"15",
          2809 => x"70",
          2810 => x"52",
          2811 => x"ff",
          2812 => x"39",
          2813 => x"81",
          2814 => x"80",
          2815 => x"52",
          2816 => x"90",
          2817 => x"80",
          2818 => x"71",
          2819 => x"7a",
          2820 => x"38",
          2821 => x"80",
          2822 => x"80",
          2823 => x"81",
          2824 => x"72",
          2825 => x"0c",
          2826 => x"04",
          2827 => x"7a",
          2828 => x"a3",
          2829 => x"88",
          2830 => x"33",
          2831 => x"56",
          2832 => x"3f",
          2833 => x"08",
          2834 => x"83",
          2835 => x"fe",
          2836 => x"87",
          2837 => x"0c",
          2838 => x"76",
          2839 => x"38",
          2840 => x"93",
          2841 => x"2b",
          2842 => x"8c",
          2843 => x"71",
          2844 => x"38",
          2845 => x"71",
          2846 => x"c6",
          2847 => x"39",
          2848 => x"81",
          2849 => x"06",
          2850 => x"71",
          2851 => x"38",
          2852 => x"8c",
          2853 => x"e8",
          2854 => x"98",
          2855 => x"71",
          2856 => x"73",
          2857 => x"92",
          2858 => x"72",
          2859 => x"06",
          2860 => x"f7",
          2861 => x"80",
          2862 => x"88",
          2863 => x"0c",
          2864 => x"80",
          2865 => x"56",
          2866 => x"56",
          2867 => x"81",
          2868 => x"88",
          2869 => x"fe",
          2870 => x"81",
          2871 => x"33",
          2872 => x"07",
          2873 => x"0c",
          2874 => x"3d",
          2875 => x"3d",
          2876 => x"11",
          2877 => x"33",
          2878 => x"71",
          2879 => x"81",
          2880 => x"72",
          2881 => x"75",
          2882 => x"81",
          2883 => x"52",
          2884 => x"54",
          2885 => x"0d",
          2886 => x"0d",
          2887 => x"05",
          2888 => x"52",
          2889 => x"70",
          2890 => x"34",
          2891 => x"51",
          2892 => x"83",
          2893 => x"ff",
          2894 => x"75",
          2895 => x"72",
          2896 => x"54",
          2897 => x"2a",
          2898 => x"70",
          2899 => x"34",
          2900 => x"51",
          2901 => x"81",
          2902 => x"70",
          2903 => x"70",
          2904 => x"3d",
          2905 => x"3d",
          2906 => x"77",
          2907 => x"70",
          2908 => x"38",
          2909 => x"05",
          2910 => x"70",
          2911 => x"34",
          2912 => x"eb",
          2913 => x"0d",
          2914 => x"0d",
          2915 => x"54",
          2916 => x"72",
          2917 => x"54",
          2918 => x"51",
          2919 => x"84",
          2920 => x"fc",
          2921 => x"77",
          2922 => x"53",
          2923 => x"05",
          2924 => x"70",
          2925 => x"33",
          2926 => x"ff",
          2927 => x"52",
          2928 => x"2e",
          2929 => x"80",
          2930 => x"71",
          2931 => x"0c",
          2932 => x"04",
          2933 => x"74",
          2934 => x"89",
          2935 => x"2e",
          2936 => x"11",
          2937 => x"52",
          2938 => x"70",
          2939 => x"c8",
          2940 => x"0d",
          2941 => x"81",
          2942 => x"04",
          2943 => x"f8",
          2944 => x"f7",
          2945 => x"56",
          2946 => x"17",
          2947 => x"74",
          2948 => x"d6",
          2949 => x"b0",
          2950 => x"b4",
          2951 => x"81",
          2952 => x"59",
          2953 => x"81",
          2954 => x"7a",
          2955 => x"06",
          2956 => x"f8",
          2957 => x"17",
          2958 => x"08",
          2959 => x"08",
          2960 => x"08",
          2961 => x"74",
          2962 => x"38",
          2963 => x"55",
          2964 => x"09",
          2965 => x"38",
          2966 => x"18",
          2967 => x"81",
          2968 => x"f9",
          2969 => x"39",
          2970 => x"81",
          2971 => x"8b",
          2972 => x"fa",
          2973 => x"7a",
          2974 => x"57",
          2975 => x"08",
          2976 => x"75",
          2977 => x"3f",
          2978 => x"08",
          2979 => x"c8",
          2980 => x"81",
          2981 => x"b4",
          2982 => x"16",
          2983 => x"be",
          2984 => x"c8",
          2985 => x"85",
          2986 => x"81",
          2987 => x"17",
          2988 => x"f8",
          2989 => x"3d",
          2990 => x"3d",
          2991 => x"52",
          2992 => x"3f",
          2993 => x"08",
          2994 => x"c8",
          2995 => x"38",
          2996 => x"74",
          2997 => x"81",
          2998 => x"38",
          2999 => x"59",
          3000 => x"09",
          3001 => x"e3",
          3002 => x"53",
          3003 => x"08",
          3004 => x"70",
          3005 => x"91",
          3006 => x"d5",
          3007 => x"17",
          3008 => x"3f",
          3009 => x"a4",
          3010 => x"51",
          3011 => x"86",
          3012 => x"f2",
          3013 => x"17",
          3014 => x"3f",
          3015 => x"52",
          3016 => x"51",
          3017 => x"8c",
          3018 => x"84",
          3019 => x"fc",
          3020 => x"17",
          3021 => x"70",
          3022 => x"79",
          3023 => x"52",
          3024 => x"51",
          3025 => x"77",
          3026 => x"80",
          3027 => x"81",
          3028 => x"f9",
          3029 => x"f8",
          3030 => x"2e",
          3031 => x"58",
          3032 => x"c8",
          3033 => x"0d",
          3034 => x"0d",
          3035 => x"98",
          3036 => x"05",
          3037 => x"80",
          3038 => x"27",
          3039 => x"14",
          3040 => x"29",
          3041 => x"05",
          3042 => x"81",
          3043 => x"87",
          3044 => x"f9",
          3045 => x"7a",
          3046 => x"54",
          3047 => x"27",
          3048 => x"76",
          3049 => x"27",
          3050 => x"ff",
          3051 => x"58",
          3052 => x"80",
          3053 => x"82",
          3054 => x"72",
          3055 => x"38",
          3056 => x"72",
          3057 => x"8e",
          3058 => x"39",
          3059 => x"17",
          3060 => x"a4",
          3061 => x"53",
          3062 => x"fd",
          3063 => x"f8",
          3064 => x"9f",
          3065 => x"ff",
          3066 => x"11",
          3067 => x"70",
          3068 => x"18",
          3069 => x"76",
          3070 => x"53",
          3071 => x"81",
          3072 => x"80",
          3073 => x"83",
          3074 => x"b4",
          3075 => x"88",
          3076 => x"79",
          3077 => x"84",
          3078 => x"58",
          3079 => x"80",
          3080 => x"9f",
          3081 => x"80",
          3082 => x"88",
          3083 => x"08",
          3084 => x"51",
          3085 => x"81",
          3086 => x"80",
          3087 => x"10",
          3088 => x"74",
          3089 => x"51",
          3090 => x"81",
          3091 => x"83",
          3092 => x"58",
          3093 => x"87",
          3094 => x"08",
          3095 => x"51",
          3096 => x"81",
          3097 => x"9b",
          3098 => x"2b",
          3099 => x"74",
          3100 => x"51",
          3101 => x"81",
          3102 => x"f0",
          3103 => x"83",
          3104 => x"77",
          3105 => x"0c",
          3106 => x"04",
          3107 => x"7a",
          3108 => x"58",
          3109 => x"81",
          3110 => x"9e",
          3111 => x"17",
          3112 => x"96",
          3113 => x"53",
          3114 => x"81",
          3115 => x"79",
          3116 => x"72",
          3117 => x"38",
          3118 => x"72",
          3119 => x"b8",
          3120 => x"39",
          3121 => x"17",
          3122 => x"a4",
          3123 => x"53",
          3124 => x"fb",
          3125 => x"f8",
          3126 => x"81",
          3127 => x"81",
          3128 => x"83",
          3129 => x"b4",
          3130 => x"78",
          3131 => x"56",
          3132 => x"76",
          3133 => x"38",
          3134 => x"9f",
          3135 => x"33",
          3136 => x"07",
          3137 => x"74",
          3138 => x"83",
          3139 => x"89",
          3140 => x"08",
          3141 => x"51",
          3142 => x"81",
          3143 => x"59",
          3144 => x"08",
          3145 => x"74",
          3146 => x"16",
          3147 => x"84",
          3148 => x"76",
          3149 => x"88",
          3150 => x"81",
          3151 => x"8f",
          3152 => x"53",
          3153 => x"80",
          3154 => x"88",
          3155 => x"08",
          3156 => x"51",
          3157 => x"81",
          3158 => x"59",
          3159 => x"08",
          3160 => x"77",
          3161 => x"06",
          3162 => x"83",
          3163 => x"05",
          3164 => x"f7",
          3165 => x"39",
          3166 => x"a4",
          3167 => x"52",
          3168 => x"ef",
          3169 => x"c8",
          3170 => x"f8",
          3171 => x"38",
          3172 => x"06",
          3173 => x"83",
          3174 => x"18",
          3175 => x"54",
          3176 => x"f6",
          3177 => x"f8",
          3178 => x"0a",
          3179 => x"52",
          3180 => x"83",
          3181 => x"83",
          3182 => x"81",
          3183 => x"8a",
          3184 => x"f8",
          3185 => x"7c",
          3186 => x"59",
          3187 => x"81",
          3188 => x"38",
          3189 => x"08",
          3190 => x"73",
          3191 => x"38",
          3192 => x"52",
          3193 => x"a4",
          3194 => x"c8",
          3195 => x"f8",
          3196 => x"f2",
          3197 => x"82",
          3198 => x"39",
          3199 => x"e6",
          3200 => x"c8",
          3201 => x"de",
          3202 => x"78",
          3203 => x"3f",
          3204 => x"08",
          3205 => x"c8",
          3206 => x"80",
          3207 => x"f8",
          3208 => x"2e",
          3209 => x"f8",
          3210 => x"2e",
          3211 => x"53",
          3212 => x"51",
          3213 => x"81",
          3214 => x"c5",
          3215 => x"08",
          3216 => x"18",
          3217 => x"57",
          3218 => x"90",
          3219 => x"90",
          3220 => x"16",
          3221 => x"54",
          3222 => x"34",
          3223 => x"78",
          3224 => x"38",
          3225 => x"81",
          3226 => x"8a",
          3227 => x"f6",
          3228 => x"7e",
          3229 => x"5b",
          3230 => x"38",
          3231 => x"58",
          3232 => x"88",
          3233 => x"08",
          3234 => x"38",
          3235 => x"39",
          3236 => x"51",
          3237 => x"81",
          3238 => x"f8",
          3239 => x"82",
          3240 => x"f8",
          3241 => x"81",
          3242 => x"ff",
          3243 => x"38",
          3244 => x"81",
          3245 => x"26",
          3246 => x"79",
          3247 => x"08",
          3248 => x"73",
          3249 => x"b9",
          3250 => x"2e",
          3251 => x"80",
          3252 => x"1a",
          3253 => x"08",
          3254 => x"38",
          3255 => x"52",
          3256 => x"af",
          3257 => x"81",
          3258 => x"81",
          3259 => x"06",
          3260 => x"f8",
          3261 => x"81",
          3262 => x"09",
          3263 => x"72",
          3264 => x"70",
          3265 => x"f8",
          3266 => x"51",
          3267 => x"73",
          3268 => x"81",
          3269 => x"80",
          3270 => x"8c",
          3271 => x"81",
          3272 => x"38",
          3273 => x"08",
          3274 => x"73",
          3275 => x"75",
          3276 => x"77",
          3277 => x"56",
          3278 => x"76",
          3279 => x"82",
          3280 => x"26",
          3281 => x"75",
          3282 => x"f8",
          3283 => x"f8",
          3284 => x"2e",
          3285 => x"59",
          3286 => x"08",
          3287 => x"81",
          3288 => x"81",
          3289 => x"59",
          3290 => x"08",
          3291 => x"70",
          3292 => x"25",
          3293 => x"51",
          3294 => x"73",
          3295 => x"75",
          3296 => x"81",
          3297 => x"38",
          3298 => x"f5",
          3299 => x"75",
          3300 => x"f9",
          3301 => x"f8",
          3302 => x"f8",
          3303 => x"70",
          3304 => x"08",
          3305 => x"51",
          3306 => x"80",
          3307 => x"73",
          3308 => x"38",
          3309 => x"52",
          3310 => x"d0",
          3311 => x"c8",
          3312 => x"a5",
          3313 => x"18",
          3314 => x"08",
          3315 => x"18",
          3316 => x"74",
          3317 => x"38",
          3318 => x"18",
          3319 => x"33",
          3320 => x"73",
          3321 => x"97",
          3322 => x"74",
          3323 => x"38",
          3324 => x"55",
          3325 => x"f8",
          3326 => x"85",
          3327 => x"75",
          3328 => x"f8",
          3329 => x"3d",
          3330 => x"3d",
          3331 => x"52",
          3332 => x"3f",
          3333 => x"08",
          3334 => x"81",
          3335 => x"80",
          3336 => x"52",
          3337 => x"c1",
          3338 => x"c8",
          3339 => x"c8",
          3340 => x"0c",
          3341 => x"53",
          3342 => x"15",
          3343 => x"f2",
          3344 => x"56",
          3345 => x"16",
          3346 => x"22",
          3347 => x"27",
          3348 => x"54",
          3349 => x"76",
          3350 => x"33",
          3351 => x"3f",
          3352 => x"08",
          3353 => x"38",
          3354 => x"76",
          3355 => x"70",
          3356 => x"9f",
          3357 => x"56",
          3358 => x"f8",
          3359 => x"3d",
          3360 => x"3d",
          3361 => x"71",
          3362 => x"57",
          3363 => x"0a",
          3364 => x"38",
          3365 => x"53",
          3366 => x"38",
          3367 => x"0c",
          3368 => x"54",
          3369 => x"75",
          3370 => x"73",
          3371 => x"a8",
          3372 => x"73",
          3373 => x"85",
          3374 => x"0b",
          3375 => x"5a",
          3376 => x"27",
          3377 => x"a8",
          3378 => x"18",
          3379 => x"39",
          3380 => x"70",
          3381 => x"58",
          3382 => x"b2",
          3383 => x"76",
          3384 => x"3f",
          3385 => x"08",
          3386 => x"c8",
          3387 => x"bd",
          3388 => x"81",
          3389 => x"27",
          3390 => x"16",
          3391 => x"c8",
          3392 => x"38",
          3393 => x"39",
          3394 => x"55",
          3395 => x"52",
          3396 => x"d5",
          3397 => x"c8",
          3398 => x"0c",
          3399 => x"0c",
          3400 => x"53",
          3401 => x"80",
          3402 => x"85",
          3403 => x"94",
          3404 => x"2a",
          3405 => x"0c",
          3406 => x"06",
          3407 => x"9c",
          3408 => x"58",
          3409 => x"c8",
          3410 => x"0d",
          3411 => x"0d",
          3412 => x"90",
          3413 => x"05",
          3414 => x"f0",
          3415 => x"27",
          3416 => x"0b",
          3417 => x"98",
          3418 => x"84",
          3419 => x"2e",
          3420 => x"76",
          3421 => x"58",
          3422 => x"38",
          3423 => x"15",
          3424 => x"08",
          3425 => x"38",
          3426 => x"88",
          3427 => x"53",
          3428 => x"81",
          3429 => x"c0",
          3430 => x"22",
          3431 => x"89",
          3432 => x"72",
          3433 => x"74",
          3434 => x"f3",
          3435 => x"f8",
          3436 => x"82",
          3437 => x"81",
          3438 => x"27",
          3439 => x"81",
          3440 => x"c8",
          3441 => x"80",
          3442 => x"16",
          3443 => x"c8",
          3444 => x"ca",
          3445 => x"38",
          3446 => x"0c",
          3447 => x"dd",
          3448 => x"08",
          3449 => x"f9",
          3450 => x"f8",
          3451 => x"87",
          3452 => x"c8",
          3453 => x"80",
          3454 => x"55",
          3455 => x"08",
          3456 => x"38",
          3457 => x"f8",
          3458 => x"2e",
          3459 => x"f8",
          3460 => x"75",
          3461 => x"3f",
          3462 => x"08",
          3463 => x"94",
          3464 => x"52",
          3465 => x"c1",
          3466 => x"c8",
          3467 => x"0c",
          3468 => x"0c",
          3469 => x"05",
          3470 => x"80",
          3471 => x"f8",
          3472 => x"3d",
          3473 => x"3d",
          3474 => x"71",
          3475 => x"57",
          3476 => x"51",
          3477 => x"81",
          3478 => x"54",
          3479 => x"08",
          3480 => x"81",
          3481 => x"56",
          3482 => x"52",
          3483 => x"83",
          3484 => x"c8",
          3485 => x"f8",
          3486 => x"d2",
          3487 => x"c8",
          3488 => x"08",
          3489 => x"54",
          3490 => x"e5",
          3491 => x"06",
          3492 => x"58",
          3493 => x"08",
          3494 => x"38",
          3495 => x"75",
          3496 => x"80",
          3497 => x"81",
          3498 => x"7a",
          3499 => x"06",
          3500 => x"39",
          3501 => x"08",
          3502 => x"76",
          3503 => x"3f",
          3504 => x"08",
          3505 => x"c8",
          3506 => x"ff",
          3507 => x"84",
          3508 => x"06",
          3509 => x"54",
          3510 => x"c8",
          3511 => x"0d",
          3512 => x"0d",
          3513 => x"52",
          3514 => x"3f",
          3515 => x"08",
          3516 => x"06",
          3517 => x"51",
          3518 => x"83",
          3519 => x"06",
          3520 => x"14",
          3521 => x"3f",
          3522 => x"08",
          3523 => x"07",
          3524 => x"f8",
          3525 => x"3d",
          3526 => x"3d",
          3527 => x"70",
          3528 => x"06",
          3529 => x"53",
          3530 => x"ed",
          3531 => x"33",
          3532 => x"83",
          3533 => x"06",
          3534 => x"90",
          3535 => x"15",
          3536 => x"3f",
          3537 => x"04",
          3538 => x"7b",
          3539 => x"84",
          3540 => x"58",
          3541 => x"80",
          3542 => x"38",
          3543 => x"52",
          3544 => x"8f",
          3545 => x"c8",
          3546 => x"f8",
          3547 => x"f5",
          3548 => x"08",
          3549 => x"53",
          3550 => x"84",
          3551 => x"39",
          3552 => x"70",
          3553 => x"81",
          3554 => x"51",
          3555 => x"16",
          3556 => x"c8",
          3557 => x"81",
          3558 => x"38",
          3559 => x"ae",
          3560 => x"81",
          3561 => x"54",
          3562 => x"2e",
          3563 => x"8f",
          3564 => x"81",
          3565 => x"76",
          3566 => x"54",
          3567 => x"09",
          3568 => x"38",
          3569 => x"7a",
          3570 => x"80",
          3571 => x"fa",
          3572 => x"f8",
          3573 => x"81",
          3574 => x"89",
          3575 => x"08",
          3576 => x"86",
          3577 => x"98",
          3578 => x"81",
          3579 => x"8b",
          3580 => x"fb",
          3581 => x"70",
          3582 => x"81",
          3583 => x"fc",
          3584 => x"f8",
          3585 => x"81",
          3586 => x"b4",
          3587 => x"08",
          3588 => x"ec",
          3589 => x"f8",
          3590 => x"81",
          3591 => x"a0",
          3592 => x"81",
          3593 => x"52",
          3594 => x"51",
          3595 => x"8b",
          3596 => x"52",
          3597 => x"51",
          3598 => x"81",
          3599 => x"34",
          3600 => x"c8",
          3601 => x"0d",
          3602 => x"0d",
          3603 => x"98",
          3604 => x"70",
          3605 => x"ec",
          3606 => x"f8",
          3607 => x"38",
          3608 => x"53",
          3609 => x"81",
          3610 => x"34",
          3611 => x"04",
          3612 => x"78",
          3613 => x"80",
          3614 => x"34",
          3615 => x"80",
          3616 => x"38",
          3617 => x"18",
          3618 => x"9c",
          3619 => x"70",
          3620 => x"56",
          3621 => x"a0",
          3622 => x"71",
          3623 => x"81",
          3624 => x"81",
          3625 => x"89",
          3626 => x"06",
          3627 => x"73",
          3628 => x"55",
          3629 => x"55",
          3630 => x"81",
          3631 => x"81",
          3632 => x"74",
          3633 => x"75",
          3634 => x"52",
          3635 => x"13",
          3636 => x"08",
          3637 => x"33",
          3638 => x"9c",
          3639 => x"11",
          3640 => x"8a",
          3641 => x"c8",
          3642 => x"96",
          3643 => x"e7",
          3644 => x"c8",
          3645 => x"23",
          3646 => x"e7",
          3647 => x"f8",
          3648 => x"17",
          3649 => x"0d",
          3650 => x"0d",
          3651 => x"5e",
          3652 => x"70",
          3653 => x"55",
          3654 => x"83",
          3655 => x"73",
          3656 => x"91",
          3657 => x"2e",
          3658 => x"1d",
          3659 => x"0c",
          3660 => x"15",
          3661 => x"70",
          3662 => x"56",
          3663 => x"09",
          3664 => x"38",
          3665 => x"80",
          3666 => x"30",
          3667 => x"78",
          3668 => x"54",
          3669 => x"73",
          3670 => x"60",
          3671 => x"54",
          3672 => x"96",
          3673 => x"0b",
          3674 => x"80",
          3675 => x"f6",
          3676 => x"f8",
          3677 => x"85",
          3678 => x"3d",
          3679 => x"5c",
          3680 => x"53",
          3681 => x"51",
          3682 => x"80",
          3683 => x"88",
          3684 => x"5c",
          3685 => x"09",
          3686 => x"d4",
          3687 => x"70",
          3688 => x"71",
          3689 => x"30",
          3690 => x"73",
          3691 => x"51",
          3692 => x"57",
          3693 => x"38",
          3694 => x"75",
          3695 => x"17",
          3696 => x"75",
          3697 => x"30",
          3698 => x"51",
          3699 => x"80",
          3700 => x"38",
          3701 => x"87",
          3702 => x"26",
          3703 => x"77",
          3704 => x"a4",
          3705 => x"27",
          3706 => x"a0",
          3707 => x"39",
          3708 => x"33",
          3709 => x"57",
          3710 => x"27",
          3711 => x"75",
          3712 => x"30",
          3713 => x"32",
          3714 => x"80",
          3715 => x"25",
          3716 => x"56",
          3717 => x"80",
          3718 => x"84",
          3719 => x"58",
          3720 => x"70",
          3721 => x"55",
          3722 => x"09",
          3723 => x"38",
          3724 => x"80",
          3725 => x"30",
          3726 => x"77",
          3727 => x"54",
          3728 => x"81",
          3729 => x"ae",
          3730 => x"06",
          3731 => x"54",
          3732 => x"74",
          3733 => x"80",
          3734 => x"7b",
          3735 => x"30",
          3736 => x"70",
          3737 => x"25",
          3738 => x"07",
          3739 => x"51",
          3740 => x"a7",
          3741 => x"8b",
          3742 => x"39",
          3743 => x"54",
          3744 => x"8c",
          3745 => x"ff",
          3746 => x"d8",
          3747 => x"54",
          3748 => x"e1",
          3749 => x"c8",
          3750 => x"b2",
          3751 => x"70",
          3752 => x"71",
          3753 => x"54",
          3754 => x"81",
          3755 => x"80",
          3756 => x"38",
          3757 => x"76",
          3758 => x"df",
          3759 => x"54",
          3760 => x"81",
          3761 => x"55",
          3762 => x"34",
          3763 => x"52",
          3764 => x"51",
          3765 => x"81",
          3766 => x"bf",
          3767 => x"16",
          3768 => x"26",
          3769 => x"16",
          3770 => x"06",
          3771 => x"17",
          3772 => x"34",
          3773 => x"fd",
          3774 => x"19",
          3775 => x"80",
          3776 => x"79",
          3777 => x"81",
          3778 => x"81",
          3779 => x"85",
          3780 => x"54",
          3781 => x"8f",
          3782 => x"86",
          3783 => x"39",
          3784 => x"f3",
          3785 => x"73",
          3786 => x"80",
          3787 => x"52",
          3788 => x"ce",
          3789 => x"c8",
          3790 => x"f8",
          3791 => x"d7",
          3792 => x"08",
          3793 => x"e6",
          3794 => x"f8",
          3795 => x"81",
          3796 => x"80",
          3797 => x"1b",
          3798 => x"55",
          3799 => x"2e",
          3800 => x"8b",
          3801 => x"06",
          3802 => x"1c",
          3803 => x"33",
          3804 => x"70",
          3805 => x"55",
          3806 => x"38",
          3807 => x"52",
          3808 => x"9f",
          3809 => x"c8",
          3810 => x"8b",
          3811 => x"7a",
          3812 => x"3f",
          3813 => x"75",
          3814 => x"57",
          3815 => x"2e",
          3816 => x"84",
          3817 => x"06",
          3818 => x"75",
          3819 => x"81",
          3820 => x"2a",
          3821 => x"73",
          3822 => x"38",
          3823 => x"54",
          3824 => x"fb",
          3825 => x"80",
          3826 => x"34",
          3827 => x"c1",
          3828 => x"06",
          3829 => x"38",
          3830 => x"39",
          3831 => x"70",
          3832 => x"54",
          3833 => x"86",
          3834 => x"84",
          3835 => x"06",
          3836 => x"73",
          3837 => x"38",
          3838 => x"83",
          3839 => x"b4",
          3840 => x"51",
          3841 => x"81",
          3842 => x"88",
          3843 => x"ea",
          3844 => x"f8",
          3845 => x"3d",
          3846 => x"3d",
          3847 => x"ff",
          3848 => x"71",
          3849 => x"5c",
          3850 => x"80",
          3851 => x"38",
          3852 => x"05",
          3853 => x"a0",
          3854 => x"71",
          3855 => x"38",
          3856 => x"71",
          3857 => x"81",
          3858 => x"38",
          3859 => x"11",
          3860 => x"06",
          3861 => x"70",
          3862 => x"38",
          3863 => x"81",
          3864 => x"05",
          3865 => x"76",
          3866 => x"38",
          3867 => x"e6",
          3868 => x"77",
          3869 => x"57",
          3870 => x"05",
          3871 => x"70",
          3872 => x"33",
          3873 => x"53",
          3874 => x"99",
          3875 => x"e0",
          3876 => x"ff",
          3877 => x"ff",
          3878 => x"70",
          3879 => x"38",
          3880 => x"81",
          3881 => x"51",
          3882 => x"9f",
          3883 => x"72",
          3884 => x"81",
          3885 => x"70",
          3886 => x"72",
          3887 => x"32",
          3888 => x"72",
          3889 => x"73",
          3890 => x"53",
          3891 => x"70",
          3892 => x"38",
          3893 => x"19",
          3894 => x"75",
          3895 => x"38",
          3896 => x"83",
          3897 => x"74",
          3898 => x"59",
          3899 => x"39",
          3900 => x"33",
          3901 => x"f8",
          3902 => x"3d",
          3903 => x"3d",
          3904 => x"80",
          3905 => x"34",
          3906 => x"17",
          3907 => x"75",
          3908 => x"3f",
          3909 => x"f8",
          3910 => x"80",
          3911 => x"16",
          3912 => x"3f",
          3913 => x"08",
          3914 => x"06",
          3915 => x"73",
          3916 => x"2e",
          3917 => x"80",
          3918 => x"0b",
          3919 => x"56",
          3920 => x"e9",
          3921 => x"06",
          3922 => x"57",
          3923 => x"32",
          3924 => x"80",
          3925 => x"51",
          3926 => x"8a",
          3927 => x"e8",
          3928 => x"06",
          3929 => x"53",
          3930 => x"52",
          3931 => x"51",
          3932 => x"81",
          3933 => x"55",
          3934 => x"08",
          3935 => x"38",
          3936 => x"e6",
          3937 => x"86",
          3938 => x"97",
          3939 => x"c8",
          3940 => x"f8",
          3941 => x"2e",
          3942 => x"55",
          3943 => x"c8",
          3944 => x"0d",
          3945 => x"0d",
          3946 => x"05",
          3947 => x"33",
          3948 => x"75",
          3949 => x"fc",
          3950 => x"f8",
          3951 => x"8b",
          3952 => x"81",
          3953 => x"24",
          3954 => x"81",
          3955 => x"84",
          3956 => x"f8",
          3957 => x"55",
          3958 => x"73",
          3959 => x"e6",
          3960 => x"0c",
          3961 => x"06",
          3962 => x"57",
          3963 => x"ae",
          3964 => x"33",
          3965 => x"3f",
          3966 => x"08",
          3967 => x"70",
          3968 => x"55",
          3969 => x"76",
          3970 => x"b8",
          3971 => x"2a",
          3972 => x"51",
          3973 => x"72",
          3974 => x"86",
          3975 => x"74",
          3976 => x"15",
          3977 => x"81",
          3978 => x"d7",
          3979 => x"f8",
          3980 => x"ff",
          3981 => x"06",
          3982 => x"56",
          3983 => x"38",
          3984 => x"8f",
          3985 => x"2a",
          3986 => x"51",
          3987 => x"72",
          3988 => x"80",
          3989 => x"52",
          3990 => x"3f",
          3991 => x"08",
          3992 => x"57",
          3993 => x"09",
          3994 => x"e2",
          3995 => x"74",
          3996 => x"56",
          3997 => x"33",
          3998 => x"72",
          3999 => x"38",
          4000 => x"51",
          4001 => x"81",
          4002 => x"57",
          4003 => x"84",
          4004 => x"ff",
          4005 => x"56",
          4006 => x"25",
          4007 => x"0b",
          4008 => x"56",
          4009 => x"05",
          4010 => x"83",
          4011 => x"2e",
          4012 => x"52",
          4013 => x"c6",
          4014 => x"c8",
          4015 => x"06",
          4016 => x"27",
          4017 => x"16",
          4018 => x"27",
          4019 => x"56",
          4020 => x"84",
          4021 => x"56",
          4022 => x"84",
          4023 => x"14",
          4024 => x"3f",
          4025 => x"08",
          4026 => x"06",
          4027 => x"80",
          4028 => x"06",
          4029 => x"80",
          4030 => x"db",
          4031 => x"f8",
          4032 => x"ff",
          4033 => x"77",
          4034 => x"d8",
          4035 => x"de",
          4036 => x"c8",
          4037 => x"9c",
          4038 => x"c4",
          4039 => x"15",
          4040 => x"14",
          4041 => x"70",
          4042 => x"51",
          4043 => x"56",
          4044 => x"84",
          4045 => x"81",
          4046 => x"71",
          4047 => x"16",
          4048 => x"53",
          4049 => x"23",
          4050 => x"8b",
          4051 => x"73",
          4052 => x"80",
          4053 => x"8d",
          4054 => x"39",
          4055 => x"51",
          4056 => x"81",
          4057 => x"53",
          4058 => x"08",
          4059 => x"72",
          4060 => x"8d",
          4061 => x"ce",
          4062 => x"14",
          4063 => x"3f",
          4064 => x"08",
          4065 => x"06",
          4066 => x"38",
          4067 => x"51",
          4068 => x"81",
          4069 => x"55",
          4070 => x"51",
          4071 => x"81",
          4072 => x"83",
          4073 => x"53",
          4074 => x"80",
          4075 => x"38",
          4076 => x"78",
          4077 => x"2a",
          4078 => x"78",
          4079 => x"86",
          4080 => x"22",
          4081 => x"31",
          4082 => x"e1",
          4083 => x"c8",
          4084 => x"f8",
          4085 => x"2e",
          4086 => x"81",
          4087 => x"80",
          4088 => x"f5",
          4089 => x"83",
          4090 => x"ff",
          4091 => x"38",
          4092 => x"9f",
          4093 => x"38",
          4094 => x"39",
          4095 => x"80",
          4096 => x"38",
          4097 => x"98",
          4098 => x"a0",
          4099 => x"1c",
          4100 => x"0c",
          4101 => x"17",
          4102 => x"76",
          4103 => x"81",
          4104 => x"80",
          4105 => x"d9",
          4106 => x"f8",
          4107 => x"ff",
          4108 => x"8d",
          4109 => x"8e",
          4110 => x"8a",
          4111 => x"14",
          4112 => x"3f",
          4113 => x"08",
          4114 => x"74",
          4115 => x"a2",
          4116 => x"79",
          4117 => x"ee",
          4118 => x"a8",
          4119 => x"15",
          4120 => x"2e",
          4121 => x"10",
          4122 => x"2a",
          4123 => x"05",
          4124 => x"ff",
          4125 => x"53",
          4126 => x"9c",
          4127 => x"81",
          4128 => x"0b",
          4129 => x"ff",
          4130 => x"0c",
          4131 => x"84",
          4132 => x"83",
          4133 => x"06",
          4134 => x"80",
          4135 => x"d8",
          4136 => x"f8",
          4137 => x"ff",
          4138 => x"72",
          4139 => x"81",
          4140 => x"38",
          4141 => x"73",
          4142 => x"3f",
          4143 => x"08",
          4144 => x"81",
          4145 => x"84",
          4146 => x"b2",
          4147 => x"87",
          4148 => x"c8",
          4149 => x"ff",
          4150 => x"82",
          4151 => x"09",
          4152 => x"c8",
          4153 => x"51",
          4154 => x"81",
          4155 => x"84",
          4156 => x"d2",
          4157 => x"06",
          4158 => x"98",
          4159 => x"ee",
          4160 => x"c8",
          4161 => x"85",
          4162 => x"09",
          4163 => x"38",
          4164 => x"51",
          4165 => x"81",
          4166 => x"90",
          4167 => x"a0",
          4168 => x"ca",
          4169 => x"c8",
          4170 => x"0c",
          4171 => x"81",
          4172 => x"81",
          4173 => x"81",
          4174 => x"72",
          4175 => x"80",
          4176 => x"0c",
          4177 => x"81",
          4178 => x"90",
          4179 => x"fb",
          4180 => x"54",
          4181 => x"80",
          4182 => x"73",
          4183 => x"80",
          4184 => x"72",
          4185 => x"80",
          4186 => x"86",
          4187 => x"15",
          4188 => x"71",
          4189 => x"81",
          4190 => x"81",
          4191 => x"d0",
          4192 => x"f8",
          4193 => x"06",
          4194 => x"38",
          4195 => x"54",
          4196 => x"80",
          4197 => x"71",
          4198 => x"81",
          4199 => x"87",
          4200 => x"fa",
          4201 => x"ab",
          4202 => x"58",
          4203 => x"05",
          4204 => x"e6",
          4205 => x"80",
          4206 => x"c8",
          4207 => x"38",
          4208 => x"08",
          4209 => x"f8",
          4210 => x"08",
          4211 => x"80",
          4212 => x"80",
          4213 => x"54",
          4214 => x"84",
          4215 => x"34",
          4216 => x"75",
          4217 => x"2e",
          4218 => x"53",
          4219 => x"53",
          4220 => x"f7",
          4221 => x"f8",
          4222 => x"73",
          4223 => x"0c",
          4224 => x"04",
          4225 => x"67",
          4226 => x"80",
          4227 => x"59",
          4228 => x"78",
          4229 => x"c8",
          4230 => x"06",
          4231 => x"3d",
          4232 => x"99",
          4233 => x"52",
          4234 => x"3f",
          4235 => x"08",
          4236 => x"c8",
          4237 => x"38",
          4238 => x"52",
          4239 => x"52",
          4240 => x"3f",
          4241 => x"08",
          4242 => x"c8",
          4243 => x"02",
          4244 => x"33",
          4245 => x"55",
          4246 => x"25",
          4247 => x"55",
          4248 => x"54",
          4249 => x"81",
          4250 => x"80",
          4251 => x"74",
          4252 => x"81",
          4253 => x"75",
          4254 => x"3f",
          4255 => x"08",
          4256 => x"02",
          4257 => x"91",
          4258 => x"81",
          4259 => x"82",
          4260 => x"06",
          4261 => x"80",
          4262 => x"88",
          4263 => x"39",
          4264 => x"58",
          4265 => x"38",
          4266 => x"70",
          4267 => x"54",
          4268 => x"81",
          4269 => x"52",
          4270 => x"a5",
          4271 => x"c8",
          4272 => x"88",
          4273 => x"62",
          4274 => x"d4",
          4275 => x"54",
          4276 => x"15",
          4277 => x"62",
          4278 => x"e8",
          4279 => x"52",
          4280 => x"51",
          4281 => x"7a",
          4282 => x"83",
          4283 => x"80",
          4284 => x"38",
          4285 => x"08",
          4286 => x"53",
          4287 => x"3d",
          4288 => x"dd",
          4289 => x"f8",
          4290 => x"81",
          4291 => x"82",
          4292 => x"39",
          4293 => x"38",
          4294 => x"33",
          4295 => x"70",
          4296 => x"55",
          4297 => x"2e",
          4298 => x"55",
          4299 => x"77",
          4300 => x"81",
          4301 => x"73",
          4302 => x"38",
          4303 => x"54",
          4304 => x"a0",
          4305 => x"82",
          4306 => x"52",
          4307 => x"a3",
          4308 => x"c8",
          4309 => x"18",
          4310 => x"55",
          4311 => x"c8",
          4312 => x"38",
          4313 => x"70",
          4314 => x"54",
          4315 => x"86",
          4316 => x"c0",
          4317 => x"b0",
          4318 => x"1b",
          4319 => x"1b",
          4320 => x"70",
          4321 => x"d9",
          4322 => x"c8",
          4323 => x"c8",
          4324 => x"0c",
          4325 => x"52",
          4326 => x"3f",
          4327 => x"08",
          4328 => x"08",
          4329 => x"77",
          4330 => x"86",
          4331 => x"1a",
          4332 => x"1a",
          4333 => x"91",
          4334 => x"0b",
          4335 => x"80",
          4336 => x"0c",
          4337 => x"70",
          4338 => x"54",
          4339 => x"81",
          4340 => x"f8",
          4341 => x"2e",
          4342 => x"81",
          4343 => x"94",
          4344 => x"17",
          4345 => x"2b",
          4346 => x"57",
          4347 => x"52",
          4348 => x"9f",
          4349 => x"c8",
          4350 => x"f8",
          4351 => x"26",
          4352 => x"55",
          4353 => x"08",
          4354 => x"81",
          4355 => x"79",
          4356 => x"31",
          4357 => x"70",
          4358 => x"25",
          4359 => x"76",
          4360 => x"81",
          4361 => x"55",
          4362 => x"38",
          4363 => x"0c",
          4364 => x"75",
          4365 => x"54",
          4366 => x"a2",
          4367 => x"7a",
          4368 => x"3f",
          4369 => x"08",
          4370 => x"55",
          4371 => x"89",
          4372 => x"c8",
          4373 => x"1a",
          4374 => x"80",
          4375 => x"54",
          4376 => x"c8",
          4377 => x"0d",
          4378 => x"0d",
          4379 => x"64",
          4380 => x"59",
          4381 => x"90",
          4382 => x"52",
          4383 => x"cf",
          4384 => x"c8",
          4385 => x"f8",
          4386 => x"38",
          4387 => x"55",
          4388 => x"86",
          4389 => x"82",
          4390 => x"19",
          4391 => x"55",
          4392 => x"80",
          4393 => x"38",
          4394 => x"0b",
          4395 => x"82",
          4396 => x"39",
          4397 => x"1a",
          4398 => x"82",
          4399 => x"19",
          4400 => x"08",
          4401 => x"7c",
          4402 => x"74",
          4403 => x"2e",
          4404 => x"94",
          4405 => x"83",
          4406 => x"56",
          4407 => x"38",
          4408 => x"22",
          4409 => x"89",
          4410 => x"55",
          4411 => x"75",
          4412 => x"19",
          4413 => x"39",
          4414 => x"52",
          4415 => x"93",
          4416 => x"c8",
          4417 => x"75",
          4418 => x"38",
          4419 => x"ff",
          4420 => x"98",
          4421 => x"19",
          4422 => x"51",
          4423 => x"81",
          4424 => x"80",
          4425 => x"38",
          4426 => x"08",
          4427 => x"2a",
          4428 => x"80",
          4429 => x"38",
          4430 => x"8a",
          4431 => x"5c",
          4432 => x"27",
          4433 => x"7a",
          4434 => x"54",
          4435 => x"52",
          4436 => x"51",
          4437 => x"81",
          4438 => x"fe",
          4439 => x"83",
          4440 => x"56",
          4441 => x"9f",
          4442 => x"08",
          4443 => x"74",
          4444 => x"38",
          4445 => x"b4",
          4446 => x"16",
          4447 => x"89",
          4448 => x"51",
          4449 => x"77",
          4450 => x"b9",
          4451 => x"1a",
          4452 => x"08",
          4453 => x"84",
          4454 => x"57",
          4455 => x"27",
          4456 => x"56",
          4457 => x"52",
          4458 => x"c7",
          4459 => x"c8",
          4460 => x"38",
          4461 => x"19",
          4462 => x"06",
          4463 => x"52",
          4464 => x"a2",
          4465 => x"31",
          4466 => x"7f",
          4467 => x"94",
          4468 => x"94",
          4469 => x"5c",
          4470 => x"80",
          4471 => x"f8",
          4472 => x"3d",
          4473 => x"3d",
          4474 => x"65",
          4475 => x"5d",
          4476 => x"0c",
          4477 => x"05",
          4478 => x"f6",
          4479 => x"f8",
          4480 => x"81",
          4481 => x"8a",
          4482 => x"33",
          4483 => x"2e",
          4484 => x"56",
          4485 => x"90",
          4486 => x"81",
          4487 => x"06",
          4488 => x"87",
          4489 => x"2e",
          4490 => x"95",
          4491 => x"91",
          4492 => x"56",
          4493 => x"81",
          4494 => x"34",
          4495 => x"8e",
          4496 => x"08",
          4497 => x"56",
          4498 => x"84",
          4499 => x"5c",
          4500 => x"82",
          4501 => x"18",
          4502 => x"ff",
          4503 => x"74",
          4504 => x"7e",
          4505 => x"ff",
          4506 => x"2a",
          4507 => x"7a",
          4508 => x"8c",
          4509 => x"08",
          4510 => x"38",
          4511 => x"39",
          4512 => x"52",
          4513 => x"e7",
          4514 => x"c8",
          4515 => x"f8",
          4516 => x"2e",
          4517 => x"74",
          4518 => x"91",
          4519 => x"2e",
          4520 => x"74",
          4521 => x"88",
          4522 => x"38",
          4523 => x"0c",
          4524 => x"15",
          4525 => x"08",
          4526 => x"06",
          4527 => x"51",
          4528 => x"81",
          4529 => x"fe",
          4530 => x"18",
          4531 => x"51",
          4532 => x"81",
          4533 => x"80",
          4534 => x"38",
          4535 => x"08",
          4536 => x"2a",
          4537 => x"80",
          4538 => x"38",
          4539 => x"8a",
          4540 => x"5b",
          4541 => x"27",
          4542 => x"7b",
          4543 => x"54",
          4544 => x"52",
          4545 => x"51",
          4546 => x"81",
          4547 => x"fe",
          4548 => x"b0",
          4549 => x"31",
          4550 => x"79",
          4551 => x"84",
          4552 => x"16",
          4553 => x"89",
          4554 => x"52",
          4555 => x"cc",
          4556 => x"55",
          4557 => x"16",
          4558 => x"2b",
          4559 => x"39",
          4560 => x"94",
          4561 => x"93",
          4562 => x"cd",
          4563 => x"f8",
          4564 => x"e3",
          4565 => x"b0",
          4566 => x"76",
          4567 => x"94",
          4568 => x"ff",
          4569 => x"71",
          4570 => x"7b",
          4571 => x"38",
          4572 => x"18",
          4573 => x"51",
          4574 => x"81",
          4575 => x"fd",
          4576 => x"53",
          4577 => x"18",
          4578 => x"06",
          4579 => x"51",
          4580 => x"7e",
          4581 => x"83",
          4582 => x"76",
          4583 => x"17",
          4584 => x"1e",
          4585 => x"18",
          4586 => x"0c",
          4587 => x"58",
          4588 => x"74",
          4589 => x"38",
          4590 => x"8c",
          4591 => x"90",
          4592 => x"33",
          4593 => x"55",
          4594 => x"34",
          4595 => x"81",
          4596 => x"90",
          4597 => x"f8",
          4598 => x"8b",
          4599 => x"53",
          4600 => x"f2",
          4601 => x"f8",
          4602 => x"81",
          4603 => x"80",
          4604 => x"16",
          4605 => x"2a",
          4606 => x"51",
          4607 => x"80",
          4608 => x"38",
          4609 => x"52",
          4610 => x"e7",
          4611 => x"c8",
          4612 => x"f8",
          4613 => x"d4",
          4614 => x"08",
          4615 => x"a0",
          4616 => x"73",
          4617 => x"88",
          4618 => x"74",
          4619 => x"51",
          4620 => x"8c",
          4621 => x"9c",
          4622 => x"fb",
          4623 => x"b2",
          4624 => x"15",
          4625 => x"3f",
          4626 => x"15",
          4627 => x"3f",
          4628 => x"0b",
          4629 => x"78",
          4630 => x"3f",
          4631 => x"08",
          4632 => x"81",
          4633 => x"57",
          4634 => x"34",
          4635 => x"c8",
          4636 => x"0d",
          4637 => x"0d",
          4638 => x"54",
          4639 => x"81",
          4640 => x"53",
          4641 => x"08",
          4642 => x"3d",
          4643 => x"73",
          4644 => x"3f",
          4645 => x"08",
          4646 => x"c8",
          4647 => x"81",
          4648 => x"74",
          4649 => x"f8",
          4650 => x"3d",
          4651 => x"3d",
          4652 => x"51",
          4653 => x"8b",
          4654 => x"81",
          4655 => x"24",
          4656 => x"f8",
          4657 => x"f9",
          4658 => x"52",
          4659 => x"c8",
          4660 => x"0d",
          4661 => x"0d",
          4662 => x"3d",
          4663 => x"94",
          4664 => x"c1",
          4665 => x"c8",
          4666 => x"f8",
          4667 => x"e0",
          4668 => x"63",
          4669 => x"d4",
          4670 => x"8d",
          4671 => x"c8",
          4672 => x"f8",
          4673 => x"38",
          4674 => x"05",
          4675 => x"2b",
          4676 => x"80",
          4677 => x"76",
          4678 => x"0c",
          4679 => x"02",
          4680 => x"70",
          4681 => x"81",
          4682 => x"56",
          4683 => x"9e",
          4684 => x"53",
          4685 => x"db",
          4686 => x"f8",
          4687 => x"15",
          4688 => x"81",
          4689 => x"84",
          4690 => x"06",
          4691 => x"55",
          4692 => x"c8",
          4693 => x"0d",
          4694 => x"0d",
          4695 => x"5b",
          4696 => x"80",
          4697 => x"ff",
          4698 => x"9f",
          4699 => x"b5",
          4700 => x"c8",
          4701 => x"f8",
          4702 => x"fc",
          4703 => x"7a",
          4704 => x"08",
          4705 => x"64",
          4706 => x"2e",
          4707 => x"a0",
          4708 => x"70",
          4709 => x"ea",
          4710 => x"c8",
          4711 => x"f8",
          4712 => x"d4",
          4713 => x"7b",
          4714 => x"3f",
          4715 => x"08",
          4716 => x"c8",
          4717 => x"38",
          4718 => x"51",
          4719 => x"81",
          4720 => x"45",
          4721 => x"51",
          4722 => x"81",
          4723 => x"57",
          4724 => x"08",
          4725 => x"80",
          4726 => x"da",
          4727 => x"f8",
          4728 => x"81",
          4729 => x"a4",
          4730 => x"7b",
          4731 => x"3f",
          4732 => x"c8",
          4733 => x"38",
          4734 => x"51",
          4735 => x"81",
          4736 => x"57",
          4737 => x"08",
          4738 => x"38",
          4739 => x"09",
          4740 => x"38",
          4741 => x"e0",
          4742 => x"dc",
          4743 => x"ff",
          4744 => x"74",
          4745 => x"3f",
          4746 => x"78",
          4747 => x"33",
          4748 => x"56",
          4749 => x"91",
          4750 => x"05",
          4751 => x"81",
          4752 => x"56",
          4753 => x"f5",
          4754 => x"54",
          4755 => x"81",
          4756 => x"80",
          4757 => x"78",
          4758 => x"55",
          4759 => x"11",
          4760 => x"18",
          4761 => x"58",
          4762 => x"34",
          4763 => x"ff",
          4764 => x"55",
          4765 => x"34",
          4766 => x"77",
          4767 => x"81",
          4768 => x"ff",
          4769 => x"55",
          4770 => x"34",
          4771 => x"f9",
          4772 => x"84",
          4773 => x"c8",
          4774 => x"70",
          4775 => x"56",
          4776 => x"76",
          4777 => x"81",
          4778 => x"70",
          4779 => x"56",
          4780 => x"82",
          4781 => x"78",
          4782 => x"80",
          4783 => x"27",
          4784 => x"19",
          4785 => x"7a",
          4786 => x"5c",
          4787 => x"55",
          4788 => x"7a",
          4789 => x"5c",
          4790 => x"2e",
          4791 => x"85",
          4792 => x"94",
          4793 => x"81",
          4794 => x"73",
          4795 => x"81",
          4796 => x"7a",
          4797 => x"38",
          4798 => x"76",
          4799 => x"0c",
          4800 => x"04",
          4801 => x"7b",
          4802 => x"fc",
          4803 => x"53",
          4804 => x"bb",
          4805 => x"c8",
          4806 => x"f8",
          4807 => x"fa",
          4808 => x"33",
          4809 => x"f2",
          4810 => x"08",
          4811 => x"27",
          4812 => x"15",
          4813 => x"2a",
          4814 => x"51",
          4815 => x"83",
          4816 => x"94",
          4817 => x"80",
          4818 => x"0c",
          4819 => x"2e",
          4820 => x"79",
          4821 => x"70",
          4822 => x"51",
          4823 => x"2e",
          4824 => x"52",
          4825 => x"fe",
          4826 => x"81",
          4827 => x"ff",
          4828 => x"70",
          4829 => x"fe",
          4830 => x"81",
          4831 => x"73",
          4832 => x"76",
          4833 => x"06",
          4834 => x"0c",
          4835 => x"98",
          4836 => x"58",
          4837 => x"39",
          4838 => x"54",
          4839 => x"73",
          4840 => x"cd",
          4841 => x"f8",
          4842 => x"81",
          4843 => x"81",
          4844 => x"38",
          4845 => x"08",
          4846 => x"9b",
          4847 => x"c8",
          4848 => x"0c",
          4849 => x"0c",
          4850 => x"81",
          4851 => x"76",
          4852 => x"38",
          4853 => x"94",
          4854 => x"94",
          4855 => x"16",
          4856 => x"2a",
          4857 => x"51",
          4858 => x"72",
          4859 => x"38",
          4860 => x"51",
          4861 => x"81",
          4862 => x"54",
          4863 => x"08",
          4864 => x"f8",
          4865 => x"a7",
          4866 => x"74",
          4867 => x"3f",
          4868 => x"08",
          4869 => x"2e",
          4870 => x"74",
          4871 => x"79",
          4872 => x"14",
          4873 => x"38",
          4874 => x"0c",
          4875 => x"94",
          4876 => x"94",
          4877 => x"83",
          4878 => x"72",
          4879 => x"38",
          4880 => x"51",
          4881 => x"81",
          4882 => x"94",
          4883 => x"91",
          4884 => x"53",
          4885 => x"81",
          4886 => x"34",
          4887 => x"39",
          4888 => x"81",
          4889 => x"05",
          4890 => x"08",
          4891 => x"08",
          4892 => x"38",
          4893 => x"0c",
          4894 => x"80",
          4895 => x"72",
          4896 => x"73",
          4897 => x"53",
          4898 => x"8c",
          4899 => x"16",
          4900 => x"38",
          4901 => x"0c",
          4902 => x"81",
          4903 => x"8b",
          4904 => x"f9",
          4905 => x"56",
          4906 => x"80",
          4907 => x"38",
          4908 => x"3d",
          4909 => x"8a",
          4910 => x"51",
          4911 => x"81",
          4912 => x"55",
          4913 => x"08",
          4914 => x"77",
          4915 => x"52",
          4916 => x"b5",
          4917 => x"c8",
          4918 => x"f8",
          4919 => x"c3",
          4920 => x"33",
          4921 => x"55",
          4922 => x"24",
          4923 => x"16",
          4924 => x"2a",
          4925 => x"51",
          4926 => x"80",
          4927 => x"9c",
          4928 => x"77",
          4929 => x"3f",
          4930 => x"08",
          4931 => x"77",
          4932 => x"22",
          4933 => x"74",
          4934 => x"ce",
          4935 => x"f8",
          4936 => x"74",
          4937 => x"81",
          4938 => x"85",
          4939 => x"74",
          4940 => x"38",
          4941 => x"74",
          4942 => x"f8",
          4943 => x"3d",
          4944 => x"3d",
          4945 => x"3d",
          4946 => x"70",
          4947 => x"ff",
          4948 => x"c8",
          4949 => x"81",
          4950 => x"73",
          4951 => x"0d",
          4952 => x"0d",
          4953 => x"3d",
          4954 => x"71",
          4955 => x"e7",
          4956 => x"f8",
          4957 => x"81",
          4958 => x"80",
          4959 => x"93",
          4960 => x"c8",
          4961 => x"51",
          4962 => x"81",
          4963 => x"53",
          4964 => x"81",
          4965 => x"52",
          4966 => x"ac",
          4967 => x"c8",
          4968 => x"f8",
          4969 => x"2e",
          4970 => x"85",
          4971 => x"87",
          4972 => x"c8",
          4973 => x"74",
          4974 => x"d5",
          4975 => x"52",
          4976 => x"89",
          4977 => x"c8",
          4978 => x"70",
          4979 => x"07",
          4980 => x"81",
          4981 => x"06",
          4982 => x"54",
          4983 => x"c8",
          4984 => x"0d",
          4985 => x"0d",
          4986 => x"53",
          4987 => x"53",
          4988 => x"56",
          4989 => x"81",
          4990 => x"55",
          4991 => x"08",
          4992 => x"52",
          4993 => x"81",
          4994 => x"c8",
          4995 => x"f8",
          4996 => x"38",
          4997 => x"05",
          4998 => x"2b",
          4999 => x"80",
          5000 => x"86",
          5001 => x"76",
          5002 => x"38",
          5003 => x"51",
          5004 => x"74",
          5005 => x"0c",
          5006 => x"04",
          5007 => x"63",
          5008 => x"80",
          5009 => x"ec",
          5010 => x"3d",
          5011 => x"3f",
          5012 => x"08",
          5013 => x"c8",
          5014 => x"38",
          5015 => x"73",
          5016 => x"08",
          5017 => x"13",
          5018 => x"58",
          5019 => x"26",
          5020 => x"7c",
          5021 => x"39",
          5022 => x"cc",
          5023 => x"81",
          5024 => x"f8",
          5025 => x"33",
          5026 => x"81",
          5027 => x"06",
          5028 => x"75",
          5029 => x"52",
          5030 => x"05",
          5031 => x"3f",
          5032 => x"08",
          5033 => x"38",
          5034 => x"08",
          5035 => x"38",
          5036 => x"08",
          5037 => x"f8",
          5038 => x"80",
          5039 => x"81",
          5040 => x"59",
          5041 => x"14",
          5042 => x"ca",
          5043 => x"39",
          5044 => x"81",
          5045 => x"57",
          5046 => x"38",
          5047 => x"18",
          5048 => x"ff",
          5049 => x"81",
          5050 => x"5b",
          5051 => x"08",
          5052 => x"7c",
          5053 => x"12",
          5054 => x"52",
          5055 => x"82",
          5056 => x"06",
          5057 => x"14",
          5058 => x"cb",
          5059 => x"c8",
          5060 => x"ff",
          5061 => x"70",
          5062 => x"82",
          5063 => x"51",
          5064 => x"b4",
          5065 => x"bb",
          5066 => x"f8",
          5067 => x"0a",
          5068 => x"70",
          5069 => x"84",
          5070 => x"51",
          5071 => x"ff",
          5072 => x"56",
          5073 => x"38",
          5074 => x"7c",
          5075 => x"0c",
          5076 => x"81",
          5077 => x"74",
          5078 => x"7a",
          5079 => x"0c",
          5080 => x"04",
          5081 => x"79",
          5082 => x"05",
          5083 => x"57",
          5084 => x"81",
          5085 => x"56",
          5086 => x"08",
          5087 => x"91",
          5088 => x"75",
          5089 => x"90",
          5090 => x"81",
          5091 => x"06",
          5092 => x"87",
          5093 => x"2e",
          5094 => x"94",
          5095 => x"73",
          5096 => x"27",
          5097 => x"73",
          5098 => x"f8",
          5099 => x"88",
          5100 => x"76",
          5101 => x"3f",
          5102 => x"08",
          5103 => x"0c",
          5104 => x"39",
          5105 => x"52",
          5106 => x"bf",
          5107 => x"f8",
          5108 => x"2e",
          5109 => x"83",
          5110 => x"81",
          5111 => x"81",
          5112 => x"06",
          5113 => x"56",
          5114 => x"a0",
          5115 => x"81",
          5116 => x"98",
          5117 => x"94",
          5118 => x"08",
          5119 => x"c8",
          5120 => x"51",
          5121 => x"81",
          5122 => x"56",
          5123 => x"8c",
          5124 => x"17",
          5125 => x"07",
          5126 => x"18",
          5127 => x"2e",
          5128 => x"91",
          5129 => x"55",
          5130 => x"c8",
          5131 => x"0d",
          5132 => x"0d",
          5133 => x"3d",
          5134 => x"52",
          5135 => x"da",
          5136 => x"f8",
          5137 => x"81",
          5138 => x"81",
          5139 => x"45",
          5140 => x"52",
          5141 => x"52",
          5142 => x"3f",
          5143 => x"08",
          5144 => x"c8",
          5145 => x"38",
          5146 => x"05",
          5147 => x"2a",
          5148 => x"51",
          5149 => x"55",
          5150 => x"38",
          5151 => x"54",
          5152 => x"81",
          5153 => x"80",
          5154 => x"70",
          5155 => x"54",
          5156 => x"81",
          5157 => x"52",
          5158 => x"c5",
          5159 => x"c8",
          5160 => x"2a",
          5161 => x"51",
          5162 => x"80",
          5163 => x"38",
          5164 => x"f8",
          5165 => x"15",
          5166 => x"86",
          5167 => x"81",
          5168 => x"5c",
          5169 => x"3d",
          5170 => x"c7",
          5171 => x"f8",
          5172 => x"81",
          5173 => x"80",
          5174 => x"f8",
          5175 => x"73",
          5176 => x"3f",
          5177 => x"08",
          5178 => x"c8",
          5179 => x"87",
          5180 => x"39",
          5181 => x"08",
          5182 => x"38",
          5183 => x"08",
          5184 => x"77",
          5185 => x"3f",
          5186 => x"08",
          5187 => x"08",
          5188 => x"f8",
          5189 => x"80",
          5190 => x"55",
          5191 => x"94",
          5192 => x"2e",
          5193 => x"53",
          5194 => x"51",
          5195 => x"81",
          5196 => x"55",
          5197 => x"78",
          5198 => x"fe",
          5199 => x"c8",
          5200 => x"81",
          5201 => x"a0",
          5202 => x"e9",
          5203 => x"53",
          5204 => x"05",
          5205 => x"51",
          5206 => x"81",
          5207 => x"54",
          5208 => x"08",
          5209 => x"78",
          5210 => x"8e",
          5211 => x"58",
          5212 => x"81",
          5213 => x"54",
          5214 => x"08",
          5215 => x"54",
          5216 => x"81",
          5217 => x"84",
          5218 => x"06",
          5219 => x"02",
          5220 => x"33",
          5221 => x"81",
          5222 => x"86",
          5223 => x"f6",
          5224 => x"74",
          5225 => x"70",
          5226 => x"c3",
          5227 => x"c8",
          5228 => x"56",
          5229 => x"08",
          5230 => x"54",
          5231 => x"08",
          5232 => x"81",
          5233 => x"82",
          5234 => x"c8",
          5235 => x"09",
          5236 => x"38",
          5237 => x"b4",
          5238 => x"b0",
          5239 => x"c8",
          5240 => x"51",
          5241 => x"81",
          5242 => x"54",
          5243 => x"08",
          5244 => x"8b",
          5245 => x"b4",
          5246 => x"b7",
          5247 => x"54",
          5248 => x"15",
          5249 => x"90",
          5250 => x"34",
          5251 => x"0a",
          5252 => x"19",
          5253 => x"9f",
          5254 => x"78",
          5255 => x"51",
          5256 => x"a0",
          5257 => x"11",
          5258 => x"05",
          5259 => x"b6",
          5260 => x"ae",
          5261 => x"15",
          5262 => x"78",
          5263 => x"53",
          5264 => x"3f",
          5265 => x"0b",
          5266 => x"77",
          5267 => x"3f",
          5268 => x"08",
          5269 => x"c8",
          5270 => x"82",
          5271 => x"52",
          5272 => x"51",
          5273 => x"3f",
          5274 => x"52",
          5275 => x"aa",
          5276 => x"90",
          5277 => x"34",
          5278 => x"0b",
          5279 => x"78",
          5280 => x"b6",
          5281 => x"c8",
          5282 => x"39",
          5283 => x"52",
          5284 => x"be",
          5285 => x"81",
          5286 => x"99",
          5287 => x"da",
          5288 => x"3d",
          5289 => x"d2",
          5290 => x"53",
          5291 => x"84",
          5292 => x"3d",
          5293 => x"3f",
          5294 => x"08",
          5295 => x"c8",
          5296 => x"38",
          5297 => x"3d",
          5298 => x"3d",
          5299 => x"cc",
          5300 => x"f8",
          5301 => x"81",
          5302 => x"82",
          5303 => x"81",
          5304 => x"81",
          5305 => x"86",
          5306 => x"aa",
          5307 => x"a4",
          5308 => x"a8",
          5309 => x"05",
          5310 => x"ea",
          5311 => x"77",
          5312 => x"70",
          5313 => x"b4",
          5314 => x"3d",
          5315 => x"51",
          5316 => x"81",
          5317 => x"55",
          5318 => x"08",
          5319 => x"6f",
          5320 => x"06",
          5321 => x"a2",
          5322 => x"92",
          5323 => x"81",
          5324 => x"f8",
          5325 => x"2e",
          5326 => x"81",
          5327 => x"51",
          5328 => x"81",
          5329 => x"55",
          5330 => x"08",
          5331 => x"68",
          5332 => x"a8",
          5333 => x"05",
          5334 => x"51",
          5335 => x"3f",
          5336 => x"33",
          5337 => x"8b",
          5338 => x"84",
          5339 => x"06",
          5340 => x"73",
          5341 => x"a0",
          5342 => x"8b",
          5343 => x"54",
          5344 => x"15",
          5345 => x"33",
          5346 => x"70",
          5347 => x"55",
          5348 => x"2e",
          5349 => x"6e",
          5350 => x"df",
          5351 => x"78",
          5352 => x"3f",
          5353 => x"08",
          5354 => x"ff",
          5355 => x"82",
          5356 => x"c8",
          5357 => x"80",
          5358 => x"f8",
          5359 => x"78",
          5360 => x"af",
          5361 => x"c8",
          5362 => x"d4",
          5363 => x"55",
          5364 => x"08",
          5365 => x"81",
          5366 => x"73",
          5367 => x"81",
          5368 => x"63",
          5369 => x"76",
          5370 => x"3f",
          5371 => x"0b",
          5372 => x"87",
          5373 => x"c8",
          5374 => x"77",
          5375 => x"3f",
          5376 => x"08",
          5377 => x"c8",
          5378 => x"78",
          5379 => x"aa",
          5380 => x"c8",
          5381 => x"81",
          5382 => x"a8",
          5383 => x"ed",
          5384 => x"80",
          5385 => x"02",
          5386 => x"df",
          5387 => x"57",
          5388 => x"3d",
          5389 => x"96",
          5390 => x"e9",
          5391 => x"c8",
          5392 => x"f8",
          5393 => x"cf",
          5394 => x"65",
          5395 => x"d4",
          5396 => x"b5",
          5397 => x"c8",
          5398 => x"f8",
          5399 => x"38",
          5400 => x"05",
          5401 => x"06",
          5402 => x"73",
          5403 => x"a7",
          5404 => x"09",
          5405 => x"71",
          5406 => x"06",
          5407 => x"55",
          5408 => x"15",
          5409 => x"81",
          5410 => x"34",
          5411 => x"b4",
          5412 => x"f8",
          5413 => x"74",
          5414 => x"0c",
          5415 => x"04",
          5416 => x"64",
          5417 => x"93",
          5418 => x"52",
          5419 => x"d1",
          5420 => x"f8",
          5421 => x"81",
          5422 => x"80",
          5423 => x"58",
          5424 => x"3d",
          5425 => x"c8",
          5426 => x"f8",
          5427 => x"81",
          5428 => x"b4",
          5429 => x"c7",
          5430 => x"a0",
          5431 => x"55",
          5432 => x"84",
          5433 => x"17",
          5434 => x"2b",
          5435 => x"96",
          5436 => x"b0",
          5437 => x"54",
          5438 => x"15",
          5439 => x"ff",
          5440 => x"81",
          5441 => x"55",
          5442 => x"c8",
          5443 => x"0d",
          5444 => x"0d",
          5445 => x"5a",
          5446 => x"3d",
          5447 => x"99",
          5448 => x"81",
          5449 => x"c8",
          5450 => x"c8",
          5451 => x"81",
          5452 => x"07",
          5453 => x"55",
          5454 => x"2e",
          5455 => x"81",
          5456 => x"55",
          5457 => x"2e",
          5458 => x"7b",
          5459 => x"80",
          5460 => x"70",
          5461 => x"be",
          5462 => x"f8",
          5463 => x"81",
          5464 => x"80",
          5465 => x"52",
          5466 => x"dc",
          5467 => x"c8",
          5468 => x"f8",
          5469 => x"38",
          5470 => x"08",
          5471 => x"08",
          5472 => x"56",
          5473 => x"19",
          5474 => x"59",
          5475 => x"74",
          5476 => x"56",
          5477 => x"ec",
          5478 => x"75",
          5479 => x"74",
          5480 => x"2e",
          5481 => x"16",
          5482 => x"33",
          5483 => x"73",
          5484 => x"38",
          5485 => x"84",
          5486 => x"06",
          5487 => x"7a",
          5488 => x"76",
          5489 => x"07",
          5490 => x"54",
          5491 => x"80",
          5492 => x"80",
          5493 => x"7b",
          5494 => x"53",
          5495 => x"93",
          5496 => x"c8",
          5497 => x"f8",
          5498 => x"38",
          5499 => x"55",
          5500 => x"56",
          5501 => x"8b",
          5502 => x"56",
          5503 => x"83",
          5504 => x"75",
          5505 => x"51",
          5506 => x"3f",
          5507 => x"08",
          5508 => x"81",
          5509 => x"98",
          5510 => x"e6",
          5511 => x"53",
          5512 => x"b8",
          5513 => x"3d",
          5514 => x"3f",
          5515 => x"08",
          5516 => x"08",
          5517 => x"f8",
          5518 => x"98",
          5519 => x"a0",
          5520 => x"70",
          5521 => x"ae",
          5522 => x"6d",
          5523 => x"81",
          5524 => x"57",
          5525 => x"74",
          5526 => x"38",
          5527 => x"81",
          5528 => x"81",
          5529 => x"52",
          5530 => x"89",
          5531 => x"c8",
          5532 => x"a5",
          5533 => x"33",
          5534 => x"54",
          5535 => x"3f",
          5536 => x"08",
          5537 => x"38",
          5538 => x"76",
          5539 => x"05",
          5540 => x"39",
          5541 => x"08",
          5542 => x"15",
          5543 => x"ff",
          5544 => x"73",
          5545 => x"38",
          5546 => x"83",
          5547 => x"56",
          5548 => x"75",
          5549 => x"81",
          5550 => x"33",
          5551 => x"2e",
          5552 => x"52",
          5553 => x"51",
          5554 => x"3f",
          5555 => x"08",
          5556 => x"ff",
          5557 => x"38",
          5558 => x"88",
          5559 => x"8a",
          5560 => x"38",
          5561 => x"ec",
          5562 => x"75",
          5563 => x"74",
          5564 => x"73",
          5565 => x"05",
          5566 => x"17",
          5567 => x"70",
          5568 => x"34",
          5569 => x"70",
          5570 => x"ff",
          5571 => x"55",
          5572 => x"26",
          5573 => x"8b",
          5574 => x"86",
          5575 => x"e5",
          5576 => x"38",
          5577 => x"99",
          5578 => x"05",
          5579 => x"70",
          5580 => x"73",
          5581 => x"81",
          5582 => x"ff",
          5583 => x"ed",
          5584 => x"80",
          5585 => x"91",
          5586 => x"55",
          5587 => x"3f",
          5588 => x"08",
          5589 => x"c8",
          5590 => x"38",
          5591 => x"51",
          5592 => x"3f",
          5593 => x"08",
          5594 => x"c8",
          5595 => x"76",
          5596 => x"67",
          5597 => x"34",
          5598 => x"81",
          5599 => x"84",
          5600 => x"06",
          5601 => x"80",
          5602 => x"2e",
          5603 => x"81",
          5604 => x"ff",
          5605 => x"81",
          5606 => x"54",
          5607 => x"08",
          5608 => x"53",
          5609 => x"08",
          5610 => x"ff",
          5611 => x"67",
          5612 => x"8b",
          5613 => x"53",
          5614 => x"51",
          5615 => x"3f",
          5616 => x"0b",
          5617 => x"79",
          5618 => x"ee",
          5619 => x"c8",
          5620 => x"55",
          5621 => x"c8",
          5622 => x"0d",
          5623 => x"0d",
          5624 => x"88",
          5625 => x"05",
          5626 => x"fc",
          5627 => x"54",
          5628 => x"d2",
          5629 => x"f8",
          5630 => x"81",
          5631 => x"82",
          5632 => x"1a",
          5633 => x"82",
          5634 => x"80",
          5635 => x"8c",
          5636 => x"78",
          5637 => x"1a",
          5638 => x"2a",
          5639 => x"51",
          5640 => x"90",
          5641 => x"82",
          5642 => x"58",
          5643 => x"81",
          5644 => x"39",
          5645 => x"22",
          5646 => x"70",
          5647 => x"56",
          5648 => x"e2",
          5649 => x"14",
          5650 => x"30",
          5651 => x"9f",
          5652 => x"c8",
          5653 => x"19",
          5654 => x"5a",
          5655 => x"81",
          5656 => x"38",
          5657 => x"77",
          5658 => x"82",
          5659 => x"56",
          5660 => x"74",
          5661 => x"ff",
          5662 => x"81",
          5663 => x"55",
          5664 => x"75",
          5665 => x"82",
          5666 => x"c8",
          5667 => x"ff",
          5668 => x"f8",
          5669 => x"2e",
          5670 => x"81",
          5671 => x"8e",
          5672 => x"56",
          5673 => x"09",
          5674 => x"38",
          5675 => x"59",
          5676 => x"77",
          5677 => x"06",
          5678 => x"87",
          5679 => x"39",
          5680 => x"ba",
          5681 => x"55",
          5682 => x"2e",
          5683 => x"15",
          5684 => x"2e",
          5685 => x"83",
          5686 => x"75",
          5687 => x"7e",
          5688 => x"a8",
          5689 => x"c8",
          5690 => x"f8",
          5691 => x"ce",
          5692 => x"16",
          5693 => x"56",
          5694 => x"38",
          5695 => x"19",
          5696 => x"8c",
          5697 => x"7d",
          5698 => x"38",
          5699 => x"0c",
          5700 => x"0c",
          5701 => x"80",
          5702 => x"73",
          5703 => x"98",
          5704 => x"05",
          5705 => x"57",
          5706 => x"26",
          5707 => x"7b",
          5708 => x"0c",
          5709 => x"81",
          5710 => x"84",
          5711 => x"54",
          5712 => x"c8",
          5713 => x"0d",
          5714 => x"0d",
          5715 => x"88",
          5716 => x"05",
          5717 => x"54",
          5718 => x"c5",
          5719 => x"56",
          5720 => x"f8",
          5721 => x"8b",
          5722 => x"f8",
          5723 => x"29",
          5724 => x"05",
          5725 => x"55",
          5726 => x"84",
          5727 => x"34",
          5728 => x"08",
          5729 => x"5f",
          5730 => x"51",
          5731 => x"3f",
          5732 => x"08",
          5733 => x"70",
          5734 => x"57",
          5735 => x"8b",
          5736 => x"82",
          5737 => x"06",
          5738 => x"56",
          5739 => x"38",
          5740 => x"05",
          5741 => x"7e",
          5742 => x"f0",
          5743 => x"c8",
          5744 => x"67",
          5745 => x"2e",
          5746 => x"82",
          5747 => x"8b",
          5748 => x"75",
          5749 => x"80",
          5750 => x"81",
          5751 => x"2e",
          5752 => x"80",
          5753 => x"38",
          5754 => x"0a",
          5755 => x"ff",
          5756 => x"55",
          5757 => x"86",
          5758 => x"8a",
          5759 => x"89",
          5760 => x"2a",
          5761 => x"77",
          5762 => x"59",
          5763 => x"81",
          5764 => x"70",
          5765 => x"07",
          5766 => x"56",
          5767 => x"38",
          5768 => x"05",
          5769 => x"7e",
          5770 => x"80",
          5771 => x"81",
          5772 => x"8a",
          5773 => x"83",
          5774 => x"06",
          5775 => x"08",
          5776 => x"74",
          5777 => x"41",
          5778 => x"56",
          5779 => x"8a",
          5780 => x"61",
          5781 => x"55",
          5782 => x"27",
          5783 => x"93",
          5784 => x"80",
          5785 => x"38",
          5786 => x"70",
          5787 => x"43",
          5788 => x"95",
          5789 => x"06",
          5790 => x"2e",
          5791 => x"77",
          5792 => x"74",
          5793 => x"83",
          5794 => x"06",
          5795 => x"82",
          5796 => x"2e",
          5797 => x"78",
          5798 => x"2e",
          5799 => x"80",
          5800 => x"ae",
          5801 => x"2a",
          5802 => x"81",
          5803 => x"56",
          5804 => x"2e",
          5805 => x"77",
          5806 => x"81",
          5807 => x"79",
          5808 => x"70",
          5809 => x"5a",
          5810 => x"86",
          5811 => x"27",
          5812 => x"52",
          5813 => x"dd",
          5814 => x"f8",
          5815 => x"29",
          5816 => x"70",
          5817 => x"55",
          5818 => x"0b",
          5819 => x"08",
          5820 => x"05",
          5821 => x"ff",
          5822 => x"27",
          5823 => x"88",
          5824 => x"ae",
          5825 => x"2a",
          5826 => x"81",
          5827 => x"56",
          5828 => x"2e",
          5829 => x"77",
          5830 => x"81",
          5831 => x"79",
          5832 => x"70",
          5833 => x"5a",
          5834 => x"86",
          5835 => x"27",
          5836 => x"52",
          5837 => x"dc",
          5838 => x"f8",
          5839 => x"84",
          5840 => x"f8",
          5841 => x"f5",
          5842 => x"81",
          5843 => x"c8",
          5844 => x"f8",
          5845 => x"71",
          5846 => x"83",
          5847 => x"5e",
          5848 => x"89",
          5849 => x"5c",
          5850 => x"1c",
          5851 => x"05",
          5852 => x"ff",
          5853 => x"70",
          5854 => x"31",
          5855 => x"57",
          5856 => x"83",
          5857 => x"06",
          5858 => x"1c",
          5859 => x"5c",
          5860 => x"1d",
          5861 => x"29",
          5862 => x"31",
          5863 => x"55",
          5864 => x"87",
          5865 => x"7c",
          5866 => x"7a",
          5867 => x"31",
          5868 => x"db",
          5869 => x"f8",
          5870 => x"7d",
          5871 => x"81",
          5872 => x"81",
          5873 => x"83",
          5874 => x"80",
          5875 => x"87",
          5876 => x"81",
          5877 => x"fd",
          5878 => x"f8",
          5879 => x"2e",
          5880 => x"80",
          5881 => x"ff",
          5882 => x"f8",
          5883 => x"a0",
          5884 => x"38",
          5885 => x"74",
          5886 => x"86",
          5887 => x"fd",
          5888 => x"81",
          5889 => x"80",
          5890 => x"83",
          5891 => x"39",
          5892 => x"08",
          5893 => x"92",
          5894 => x"b8",
          5895 => x"59",
          5896 => x"27",
          5897 => x"86",
          5898 => x"55",
          5899 => x"09",
          5900 => x"38",
          5901 => x"f5",
          5902 => x"38",
          5903 => x"55",
          5904 => x"86",
          5905 => x"80",
          5906 => x"7a",
          5907 => x"b9",
          5908 => x"81",
          5909 => x"7a",
          5910 => x"8a",
          5911 => x"52",
          5912 => x"ff",
          5913 => x"79",
          5914 => x"7b",
          5915 => x"06",
          5916 => x"51",
          5917 => x"3f",
          5918 => x"1c",
          5919 => x"32",
          5920 => x"96",
          5921 => x"06",
          5922 => x"91",
          5923 => x"a1",
          5924 => x"55",
          5925 => x"ff",
          5926 => x"74",
          5927 => x"06",
          5928 => x"51",
          5929 => x"3f",
          5930 => x"52",
          5931 => x"ff",
          5932 => x"f8",
          5933 => x"34",
          5934 => x"1b",
          5935 => x"d9",
          5936 => x"52",
          5937 => x"ff",
          5938 => x"60",
          5939 => x"51",
          5940 => x"3f",
          5941 => x"09",
          5942 => x"cb",
          5943 => x"b2",
          5944 => x"c3",
          5945 => x"a0",
          5946 => x"52",
          5947 => x"ff",
          5948 => x"82",
          5949 => x"51",
          5950 => x"3f",
          5951 => x"1b",
          5952 => x"95",
          5953 => x"b2",
          5954 => x"a0",
          5955 => x"80",
          5956 => x"1c",
          5957 => x"80",
          5958 => x"93",
          5959 => x"a0",
          5960 => x"1b",
          5961 => x"82",
          5962 => x"52",
          5963 => x"ff",
          5964 => x"7c",
          5965 => x"06",
          5966 => x"51",
          5967 => x"3f",
          5968 => x"a4",
          5969 => x"0b",
          5970 => x"93",
          5971 => x"b4",
          5972 => x"51",
          5973 => x"3f",
          5974 => x"52",
          5975 => x"70",
          5976 => x"9f",
          5977 => x"54",
          5978 => x"52",
          5979 => x"9b",
          5980 => x"56",
          5981 => x"08",
          5982 => x"7d",
          5983 => x"81",
          5984 => x"38",
          5985 => x"86",
          5986 => x"52",
          5987 => x"9b",
          5988 => x"80",
          5989 => x"7a",
          5990 => x"ed",
          5991 => x"85",
          5992 => x"7a",
          5993 => x"8f",
          5994 => x"85",
          5995 => x"83",
          5996 => x"ff",
          5997 => x"ff",
          5998 => x"e8",
          5999 => x"9e",
          6000 => x"52",
          6001 => x"51",
          6002 => x"3f",
          6003 => x"52",
          6004 => x"9e",
          6005 => x"54",
          6006 => x"53",
          6007 => x"51",
          6008 => x"3f",
          6009 => x"16",
          6010 => x"7e",
          6011 => x"d8",
          6012 => x"80",
          6013 => x"ff",
          6014 => x"7f",
          6015 => x"7d",
          6016 => x"81",
          6017 => x"f8",
          6018 => x"ff",
          6019 => x"ff",
          6020 => x"51",
          6021 => x"3f",
          6022 => x"88",
          6023 => x"39",
          6024 => x"f8",
          6025 => x"2e",
          6026 => x"55",
          6027 => x"51",
          6028 => x"3f",
          6029 => x"57",
          6030 => x"83",
          6031 => x"76",
          6032 => x"7a",
          6033 => x"ff",
          6034 => x"81",
          6035 => x"82",
          6036 => x"80",
          6037 => x"c8",
          6038 => x"51",
          6039 => x"3f",
          6040 => x"78",
          6041 => x"74",
          6042 => x"18",
          6043 => x"2e",
          6044 => x"79",
          6045 => x"2e",
          6046 => x"55",
          6047 => x"62",
          6048 => x"74",
          6049 => x"75",
          6050 => x"7e",
          6051 => x"b8",
          6052 => x"c8",
          6053 => x"38",
          6054 => x"78",
          6055 => x"74",
          6056 => x"56",
          6057 => x"93",
          6058 => x"66",
          6059 => x"26",
          6060 => x"56",
          6061 => x"83",
          6062 => x"64",
          6063 => x"77",
          6064 => x"84",
          6065 => x"52",
          6066 => x"9d",
          6067 => x"d4",
          6068 => x"51",
          6069 => x"3f",
          6070 => x"55",
          6071 => x"81",
          6072 => x"34",
          6073 => x"16",
          6074 => x"16",
          6075 => x"16",
          6076 => x"05",
          6077 => x"c1",
          6078 => x"fe",
          6079 => x"fe",
          6080 => x"34",
          6081 => x"08",
          6082 => x"07",
          6083 => x"16",
          6084 => x"c8",
          6085 => x"34",
          6086 => x"c6",
          6087 => x"9c",
          6088 => x"52",
          6089 => x"51",
          6090 => x"3f",
          6091 => x"53",
          6092 => x"51",
          6093 => x"3f",
          6094 => x"f8",
          6095 => x"38",
          6096 => x"52",
          6097 => x"99",
          6098 => x"56",
          6099 => x"08",
          6100 => x"39",
          6101 => x"39",
          6102 => x"39",
          6103 => x"08",
          6104 => x"f8",
          6105 => x"3d",
          6106 => x"3d",
          6107 => x"5b",
          6108 => x"60",
          6109 => x"57",
          6110 => x"25",
          6111 => x"3d",
          6112 => x"55",
          6113 => x"15",
          6114 => x"c9",
          6115 => x"81",
          6116 => x"06",
          6117 => x"3d",
          6118 => x"8d",
          6119 => x"74",
          6120 => x"05",
          6121 => x"17",
          6122 => x"2e",
          6123 => x"c9",
          6124 => x"34",
          6125 => x"83",
          6126 => x"74",
          6127 => x"0c",
          6128 => x"04",
          6129 => x"7b",
          6130 => x"b3",
          6131 => x"57",
          6132 => x"09",
          6133 => x"38",
          6134 => x"51",
          6135 => x"17",
          6136 => x"76",
          6137 => x"88",
          6138 => x"17",
          6139 => x"59",
          6140 => x"81",
          6141 => x"76",
          6142 => x"8b",
          6143 => x"54",
          6144 => x"17",
          6145 => x"51",
          6146 => x"79",
          6147 => x"30",
          6148 => x"9f",
          6149 => x"53",
          6150 => x"75",
          6151 => x"81",
          6152 => x"0c",
          6153 => x"04",
          6154 => x"79",
          6155 => x"56",
          6156 => x"24",
          6157 => x"3d",
          6158 => x"74",
          6159 => x"52",
          6160 => x"cb",
          6161 => x"f8",
          6162 => x"38",
          6163 => x"78",
          6164 => x"06",
          6165 => x"16",
          6166 => x"39",
          6167 => x"81",
          6168 => x"89",
          6169 => x"fd",
          6170 => x"54",
          6171 => x"80",
          6172 => x"ff",
          6173 => x"76",
          6174 => x"3d",
          6175 => x"3d",
          6176 => x"e3",
          6177 => x"53",
          6178 => x"53",
          6179 => x"3f",
          6180 => x"51",
          6181 => x"72",
          6182 => x"3f",
          6183 => x"04",
          6184 => x"7a",
          6185 => x"56",
          6186 => x"80",
          6187 => x"38",
          6188 => x"15",
          6189 => x"16",
          6190 => x"d4",
          6191 => x"54",
          6192 => x"09",
          6193 => x"38",
          6194 => x"f1",
          6195 => x"76",
          6196 => x"f5",
          6197 => x"08",
          6198 => x"da",
          6199 => x"f8",
          6200 => x"f8",
          6201 => x"75",
          6202 => x"52",
          6203 => x"c0",
          6204 => x"c8",
          6205 => x"84",
          6206 => x"73",
          6207 => x"b2",
          6208 => x"70",
          6209 => x"58",
          6210 => x"27",
          6211 => x"54",
          6212 => x"c8",
          6213 => x"0d",
          6214 => x"0d",
          6215 => x"93",
          6216 => x"38",
          6217 => x"81",
          6218 => x"52",
          6219 => x"81",
          6220 => x"81",
          6221 => x"e9",
          6222 => x"f9",
          6223 => x"d4",
          6224 => x"39",
          6225 => x"51",
          6226 => x"81",
          6227 => x"80",
          6228 => x"ea",
          6229 => x"dd",
          6230 => x"9c",
          6231 => x"39",
          6232 => x"51",
          6233 => x"81",
          6234 => x"80",
          6235 => x"ea",
          6236 => x"c1",
          6237 => x"f4",
          6238 => x"81",
          6239 => x"b5",
          6240 => x"a4",
          6241 => x"81",
          6242 => x"a9",
          6243 => x"e4",
          6244 => x"81",
          6245 => x"9d",
          6246 => x"98",
          6247 => x"81",
          6248 => x"91",
          6249 => x"c8",
          6250 => x"81",
          6251 => x"85",
          6252 => x"ec",
          6253 => x"ae",
          6254 => x"0d",
          6255 => x"0d",
          6256 => x"56",
          6257 => x"26",
          6258 => x"52",
          6259 => x"29",
          6260 => x"87",
          6261 => x"51",
          6262 => x"3f",
          6263 => x"08",
          6264 => x"fe",
          6265 => x"81",
          6266 => x"54",
          6267 => x"52",
          6268 => x"51",
          6269 => x"3f",
          6270 => x"04",
          6271 => x"66",
          6272 => x"80",
          6273 => x"5b",
          6274 => x"78",
          6275 => x"07",
          6276 => x"57",
          6277 => x"56",
          6278 => x"26",
          6279 => x"56",
          6280 => x"70",
          6281 => x"51",
          6282 => x"74",
          6283 => x"81",
          6284 => x"8c",
          6285 => x"56",
          6286 => x"3f",
          6287 => x"08",
          6288 => x"c8",
          6289 => x"81",
          6290 => x"87",
          6291 => x"0c",
          6292 => x"08",
          6293 => x"d4",
          6294 => x"80",
          6295 => x"75",
          6296 => x"3f",
          6297 => x"08",
          6298 => x"c8",
          6299 => x"7a",
          6300 => x"2e",
          6301 => x"19",
          6302 => x"59",
          6303 => x"3d",
          6304 => x"cb",
          6305 => x"30",
          6306 => x"80",
          6307 => x"70",
          6308 => x"06",
          6309 => x"56",
          6310 => x"90",
          6311 => x"a0",
          6312 => x"98",
          6313 => x"78",
          6314 => x"3f",
          6315 => x"81",
          6316 => x"96",
          6317 => x"f9",
          6318 => x"02",
          6319 => x"05",
          6320 => x"ff",
          6321 => x"7a",
          6322 => x"fe",
          6323 => x"f8",
          6324 => x"38",
          6325 => x"88",
          6326 => x"2e",
          6327 => x"39",
          6328 => x"54",
          6329 => x"53",
          6330 => x"51",
          6331 => x"f8",
          6332 => x"83",
          6333 => x"76",
          6334 => x"0c",
          6335 => x"04",
          6336 => x"7f",
          6337 => x"8c",
          6338 => x"05",
          6339 => x"15",
          6340 => x"5c",
          6341 => x"5e",
          6342 => x"ed",
          6343 => x"f5",
          6344 => x"ed",
          6345 => x"ef",
          6346 => x"55",
          6347 => x"80",
          6348 => x"90",
          6349 => x"7b",
          6350 => x"38",
          6351 => x"74",
          6352 => x"7a",
          6353 => x"72",
          6354 => x"ed",
          6355 => x"f4",
          6356 => x"39",
          6357 => x"51",
          6358 => x"3f",
          6359 => x"80",
          6360 => x"18",
          6361 => x"27",
          6362 => x"08",
          6363 => x"a8",
          6364 => x"d6",
          6365 => x"81",
          6366 => x"fe",
          6367 => x"84",
          6368 => x"39",
          6369 => x"72",
          6370 => x"38",
          6371 => x"81",
          6372 => x"fe",
          6373 => x"89",
          6374 => x"d0",
          6375 => x"c6",
          6376 => x"55",
          6377 => x"ed",
          6378 => x"80",
          6379 => x"d4",
          6380 => x"b2",
          6381 => x"74",
          6382 => x"38",
          6383 => x"33",
          6384 => x"56",
          6385 => x"83",
          6386 => x"80",
          6387 => x"27",
          6388 => x"53",
          6389 => x"70",
          6390 => x"51",
          6391 => x"2e",
          6392 => x"80",
          6393 => x"38",
          6394 => x"39",
          6395 => x"ed",
          6396 => x"15",
          6397 => x"81",
          6398 => x"fe",
          6399 => x"78",
          6400 => x"5c",
          6401 => x"d7",
          6402 => x"c8",
          6403 => x"70",
          6404 => x"57",
          6405 => x"09",
          6406 => x"38",
          6407 => x"3f",
          6408 => x"08",
          6409 => x"98",
          6410 => x"32",
          6411 => x"9b",
          6412 => x"70",
          6413 => x"75",
          6414 => x"58",
          6415 => x"51",
          6416 => x"24",
          6417 => x"9b",
          6418 => x"06",
          6419 => x"53",
          6420 => x"1e",
          6421 => x"26",
          6422 => x"ff",
          6423 => x"f8",
          6424 => x"3d",
          6425 => x"3d",
          6426 => x"05",
          6427 => x"dc",
          6428 => x"e0",
          6429 => x"f2",
          6430 => x"f3",
          6431 => x"fe",
          6432 => x"81",
          6433 => x"81",
          6434 => x"81",
          6435 => x"52",
          6436 => x"51",
          6437 => x"3f",
          6438 => x"85",
          6439 => x"e3",
          6440 => x"0d",
          6441 => x"0d",
          6442 => x"80",
          6443 => x"e7",
          6444 => x"51",
          6445 => x"3f",
          6446 => x"51",
          6447 => x"3f",
          6448 => x"d9",
          6449 => x"81",
          6450 => x"06",
          6451 => x"80",
          6452 => x"81",
          6453 => x"9b",
          6454 => x"b4",
          6455 => x"93",
          6456 => x"fe",
          6457 => x"72",
          6458 => x"81",
          6459 => x"71",
          6460 => x"38",
          6461 => x"d8",
          6462 => x"ee",
          6463 => x"da",
          6464 => x"51",
          6465 => x"3f",
          6466 => x"70",
          6467 => x"52",
          6468 => x"95",
          6469 => x"fe",
          6470 => x"81",
          6471 => x"fe",
          6472 => x"80",
          6473 => x"cb",
          6474 => x"2a",
          6475 => x"51",
          6476 => x"2e",
          6477 => x"51",
          6478 => x"3f",
          6479 => x"51",
          6480 => x"3f",
          6481 => x"d8",
          6482 => x"85",
          6483 => x"06",
          6484 => x"80",
          6485 => x"81",
          6486 => x"97",
          6487 => x"80",
          6488 => x"8f",
          6489 => x"fe",
          6490 => x"72",
          6491 => x"81",
          6492 => x"71",
          6493 => x"38",
          6494 => x"d7",
          6495 => x"ef",
          6496 => x"d9",
          6497 => x"51",
          6498 => x"3f",
          6499 => x"70",
          6500 => x"52",
          6501 => x"95",
          6502 => x"fe",
          6503 => x"81",
          6504 => x"fe",
          6505 => x"80",
          6506 => x"c7",
          6507 => x"2a",
          6508 => x"51",
          6509 => x"2e",
          6510 => x"51",
          6511 => x"3f",
          6512 => x"51",
          6513 => x"3f",
          6514 => x"d7",
          6515 => x"e5",
          6516 => x"3d",
          6517 => x"3d",
          6518 => x"84",
          6519 => x"33",
          6520 => x"56",
          6521 => x"51",
          6522 => x"3f",
          6523 => x"33",
          6524 => x"38",
          6525 => x"ef",
          6526 => x"8f",
          6527 => x"b8",
          6528 => x"f8",
          6529 => x"70",
          6530 => x"08",
          6531 => x"82",
          6532 => x"51",
          6533 => x"f5",
          6534 => x"f5",
          6535 => x"73",
          6536 => x"81",
          6537 => x"82",
          6538 => x"74",
          6539 => x"f2",
          6540 => x"f8",
          6541 => x"2e",
          6542 => x"f8",
          6543 => x"fe",
          6544 => x"8e",
          6545 => x"e0",
          6546 => x"3f",
          6547 => x"f5",
          6548 => x"f5",
          6549 => x"73",
          6550 => x"81",
          6551 => x"74",
          6552 => x"fe",
          6553 => x"80",
          6554 => x"c8",
          6555 => x"0d",
          6556 => x"0d",
          6557 => x"82",
          6558 => x"5f",
          6559 => x"7c",
          6560 => x"db",
          6561 => x"c8",
          6562 => x"06",
          6563 => x"2e",
          6564 => x"a2",
          6565 => x"8c",
          6566 => x"70",
          6567 => x"ee",
          6568 => x"53",
          6569 => x"fa",
          6570 => x"b5",
          6571 => x"f8",
          6572 => x"2e",
          6573 => x"f0",
          6574 => x"bc",
          6575 => x"5f",
          6576 => x"c8",
          6577 => x"9e",
          6578 => x"70",
          6579 => x"f8",
          6580 => x"fe",
          6581 => x"3d",
          6582 => x"51",
          6583 => x"81",
          6584 => x"90",
          6585 => x"2c",
          6586 => x"80",
          6587 => x"b3",
          6588 => x"c2",
          6589 => x"78",
          6590 => x"d5",
          6591 => x"24",
          6592 => x"80",
          6593 => x"38",
          6594 => x"80",
          6595 => x"e9",
          6596 => x"c0",
          6597 => x"38",
          6598 => x"24",
          6599 => x"78",
          6600 => x"92",
          6601 => x"39",
          6602 => x"2e",
          6603 => x"78",
          6604 => x"92",
          6605 => x"c3",
          6606 => x"38",
          6607 => x"2e",
          6608 => x"8a",
          6609 => x"81",
          6610 => x"99",
          6611 => x"83",
          6612 => x"78",
          6613 => x"89",
          6614 => x"9d",
          6615 => x"85",
          6616 => x"38",
          6617 => x"b4",
          6618 => x"11",
          6619 => x"05",
          6620 => x"cb",
          6621 => x"c8",
          6622 => x"fe",
          6623 => x"3d",
          6624 => x"53",
          6625 => x"51",
          6626 => x"3f",
          6627 => x"08",
          6628 => x"ad",
          6629 => x"fe",
          6630 => x"ff",
          6631 => x"fe",
          6632 => x"81",
          6633 => x"86",
          6634 => x"c8",
          6635 => x"f0",
          6636 => x"e6",
          6637 => x"63",
          6638 => x"7b",
          6639 => x"38",
          6640 => x"7a",
          6641 => x"5c",
          6642 => x"26",
          6643 => x"e1",
          6644 => x"ff",
          6645 => x"ff",
          6646 => x"fe",
          6647 => x"81",
          6648 => x"80",
          6649 => x"38",
          6650 => x"fc",
          6651 => x"84",
          6652 => x"ed",
          6653 => x"f8",
          6654 => x"2e",
          6655 => x"b4",
          6656 => x"11",
          6657 => x"05",
          6658 => x"b3",
          6659 => x"c8",
          6660 => x"fd",
          6661 => x"f0",
          6662 => x"e5",
          6663 => x"5a",
          6664 => x"81",
          6665 => x"59",
          6666 => x"05",
          6667 => x"34",
          6668 => x"42",
          6669 => x"3d",
          6670 => x"53",
          6671 => x"51",
          6672 => x"3f",
          6673 => x"08",
          6674 => x"f5",
          6675 => x"fe",
          6676 => x"ff",
          6677 => x"fe",
          6678 => x"81",
          6679 => x"80",
          6680 => x"38",
          6681 => x"f8",
          6682 => x"84",
          6683 => x"ec",
          6684 => x"f8",
          6685 => x"2e",
          6686 => x"81",
          6687 => x"fe",
          6688 => x"63",
          6689 => x"27",
          6690 => x"70",
          6691 => x"5e",
          6692 => x"7c",
          6693 => x"78",
          6694 => x"79",
          6695 => x"52",
          6696 => x"51",
          6697 => x"3f",
          6698 => x"81",
          6699 => x"d5",
          6700 => x"90",
          6701 => x"39",
          6702 => x"80",
          6703 => x"84",
          6704 => x"eb",
          6705 => x"f8",
          6706 => x"df",
          6707 => x"8c",
          6708 => x"80",
          6709 => x"81",
          6710 => x"44",
          6711 => x"81",
          6712 => x"59",
          6713 => x"88",
          6714 => x"cc",
          6715 => x"39",
          6716 => x"33",
          6717 => x"2e",
          6718 => x"f3",
          6719 => x"ab",
          6720 => x"8f",
          6721 => x"80",
          6722 => x"81",
          6723 => x"44",
          6724 => x"f4",
          6725 => x"78",
          6726 => x"38",
          6727 => x"08",
          6728 => x"81",
          6729 => x"fc",
          6730 => x"b4",
          6731 => x"11",
          6732 => x"05",
          6733 => x"87",
          6734 => x"c8",
          6735 => x"38",
          6736 => x"33",
          6737 => x"2e",
          6738 => x"f3",
          6739 => x"80",
          6740 => x"f4",
          6741 => x"78",
          6742 => x"38",
          6743 => x"08",
          6744 => x"81",
          6745 => x"59",
          6746 => x"88",
          6747 => x"d8",
          6748 => x"39",
          6749 => x"33",
          6750 => x"2e",
          6751 => x"f3",
          6752 => x"99",
          6753 => x"8a",
          6754 => x"80",
          6755 => x"81",
          6756 => x"43",
          6757 => x"f3",
          6758 => x"05",
          6759 => x"fe",
          6760 => x"ff",
          6761 => x"fe",
          6762 => x"81",
          6763 => x"80",
          6764 => x"80",
          6765 => x"7a",
          6766 => x"38",
          6767 => x"90",
          6768 => x"70",
          6769 => x"2a",
          6770 => x"51",
          6771 => x"78",
          6772 => x"38",
          6773 => x"83",
          6774 => x"81",
          6775 => x"fe",
          6776 => x"a0",
          6777 => x"61",
          6778 => x"63",
          6779 => x"3f",
          6780 => x"51",
          6781 => x"3f",
          6782 => x"b4",
          6783 => x"11",
          6784 => x"05",
          6785 => x"b7",
          6786 => x"c8",
          6787 => x"f9",
          6788 => x"3d",
          6789 => x"53",
          6790 => x"51",
          6791 => x"3f",
          6792 => x"08",
          6793 => x"38",
          6794 => x"80",
          6795 => x"79",
          6796 => x"05",
          6797 => x"fe",
          6798 => x"ff",
          6799 => x"fe",
          6800 => x"81",
          6801 => x"e0",
          6802 => x"39",
          6803 => x"54",
          6804 => x"b0",
          6805 => x"f2",
          6806 => x"52",
          6807 => x"e7",
          6808 => x"45",
          6809 => x"78",
          6810 => x"d5",
          6811 => x"27",
          6812 => x"3d",
          6813 => x"53",
          6814 => x"51",
          6815 => x"3f",
          6816 => x"08",
          6817 => x"38",
          6818 => x"80",
          6819 => x"79",
          6820 => x"05",
          6821 => x"39",
          6822 => x"51",
          6823 => x"3f",
          6824 => x"b4",
          6825 => x"11",
          6826 => x"05",
          6827 => x"81",
          6828 => x"c8",
          6829 => x"f8",
          6830 => x"3d",
          6831 => x"53",
          6832 => x"51",
          6833 => x"3f",
          6834 => x"08",
          6835 => x"38",
          6836 => x"be",
          6837 => x"70",
          6838 => x"23",
          6839 => x"3d",
          6840 => x"53",
          6841 => x"51",
          6842 => x"3f",
          6843 => x"08",
          6844 => x"cd",
          6845 => x"22",
          6846 => x"f1",
          6847 => x"e5",
          6848 => x"f8",
          6849 => x"fe",
          6850 => x"79",
          6851 => x"59",
          6852 => x"f7",
          6853 => x"9f",
          6854 => x"60",
          6855 => x"d5",
          6856 => x"fe",
          6857 => x"ff",
          6858 => x"fe",
          6859 => x"81",
          6860 => x"80",
          6861 => x"60",
          6862 => x"05",
          6863 => x"82",
          6864 => x"78",
          6865 => x"39",
          6866 => x"51",
          6867 => x"3f",
          6868 => x"b4",
          6869 => x"11",
          6870 => x"05",
          6871 => x"d1",
          6872 => x"c8",
          6873 => x"f6",
          6874 => x"3d",
          6875 => x"53",
          6876 => x"51",
          6877 => x"3f",
          6878 => x"08",
          6879 => x"38",
          6880 => x"0c",
          6881 => x"05",
          6882 => x"fe",
          6883 => x"ff",
          6884 => x"fe",
          6885 => x"81",
          6886 => x"e4",
          6887 => x"39",
          6888 => x"54",
          6889 => x"d0",
          6890 => x"9e",
          6891 => x"52",
          6892 => x"e4",
          6893 => x"45",
          6894 => x"78",
          6895 => x"81",
          6896 => x"27",
          6897 => x"3d",
          6898 => x"53",
          6899 => x"51",
          6900 => x"3f",
          6901 => x"08",
          6902 => x"38",
          6903 => x"0c",
          6904 => x"05",
          6905 => x"39",
          6906 => x"51",
          6907 => x"3f",
          6908 => x"b4",
          6909 => x"11",
          6910 => x"05",
          6911 => x"bf",
          6912 => x"c8",
          6913 => x"f5",
          6914 => x"52",
          6915 => x"51",
          6916 => x"3f",
          6917 => x"04",
          6918 => x"80",
          6919 => x"84",
          6920 => x"e5",
          6921 => x"f8",
          6922 => x"2e",
          6923 => x"63",
          6924 => x"f8",
          6925 => x"92",
          6926 => x"78",
          6927 => x"c8",
          6928 => x"f4",
          6929 => x"f8",
          6930 => x"81",
          6931 => x"fe",
          6932 => x"f4",
          6933 => x"f2",
          6934 => x"dd",
          6935 => x"ba",
          6936 => x"dd",
          6937 => x"cc",
          6938 => x"fa",
          6939 => x"ff",
          6940 => x"d3",
          6941 => x"c9",
          6942 => x"79",
          6943 => x"80",
          6944 => x"38",
          6945 => x"59",
          6946 => x"81",
          6947 => x"3d",
          6948 => x"51",
          6949 => x"3f",
          6950 => x"08",
          6951 => x"7a",
          6952 => x"38",
          6953 => x"89",
          6954 => x"2e",
          6955 => x"cd",
          6956 => x"2e",
          6957 => x"c5",
          6958 => x"e0",
          6959 => x"81",
          6960 => x"80",
          6961 => x"e8",
          6962 => x"ff",
          6963 => x"fe",
          6964 => x"bb",
          6965 => x"88",
          6966 => x"ff",
          6967 => x"fe",
          6968 => x"ab",
          6969 => x"81",
          6970 => x"80",
          6971 => x"f8",
          6972 => x"ff",
          6973 => x"fe",
          6974 => x"93",
          6975 => x"80",
          6976 => x"84",
          6977 => x"ff",
          6978 => x"fe",
          6979 => x"81",
          6980 => x"81",
          6981 => x"80",
          6982 => x"80",
          6983 => x"80",
          6984 => x"80",
          6985 => x"ff",
          6986 => x"eb",
          6987 => x"f8",
          6988 => x"f8",
          6989 => x"70",
          6990 => x"07",
          6991 => x"5b",
          6992 => x"5a",
          6993 => x"83",
          6994 => x"78",
          6995 => x"78",
          6996 => x"38",
          6997 => x"81",
          6998 => x"59",
          6999 => x"38",
          7000 => x"7d",
          7001 => x"59",
          7002 => x"7e",
          7003 => x"81",
          7004 => x"38",
          7005 => x"51",
          7006 => x"3f",
          7007 => x"fc",
          7008 => x"0b",
          7009 => x"34",
          7010 => x"8c",
          7011 => x"55",
          7012 => x"52",
          7013 => x"b8",
          7014 => x"f8",
          7015 => x"2b",
          7016 => x"53",
          7017 => x"52",
          7018 => x"b8",
          7019 => x"81",
          7020 => x"07",
          7021 => x"c0",
          7022 => x"08",
          7023 => x"84",
          7024 => x"51",
          7025 => x"3f",
          7026 => x"08",
          7027 => x"08",
          7028 => x"84",
          7029 => x"51",
          7030 => x"3f",
          7031 => x"c8",
          7032 => x"0c",
          7033 => x"0b",
          7034 => x"84",
          7035 => x"83",
          7036 => x"94",
          7037 => x"8b",
          7038 => x"dc",
          7039 => x"0b",
          7040 => x"0c",
          7041 => x"3f",
          7042 => x"3f",
          7043 => x"51",
          7044 => x"3f",
          7045 => x"51",
          7046 => x"3f",
          7047 => x"51",
          7048 => x"3f",
          7049 => x"be",
          7050 => x"3f",
          7051 => x"ff",
          7052 => x"00",
          7053 => x"ff",
          7054 => x"ff",
          7055 => x"00",
          7056 => x"00",
          7057 => x"00",
          7058 => x"00",
          7059 => x"00",
          7060 => x"00",
          7061 => x"00",
          7062 => x"00",
          7063 => x"00",
          7064 => x"00",
          7065 => x"00",
          7066 => x"00",
          7067 => x"00",
          7068 => x"00",
          7069 => x"00",
          7070 => x"00",
          7071 => x"00",
          7072 => x"00",
          7073 => x"00",
          7074 => x"00",
          7075 => x"00",
          7076 => x"00",
          7077 => x"00",
          7078 => x"00",
          7079 => x"00",
          7080 => x"00",
          7081 => x"00",
          7082 => x"00",
          7083 => x"00",
          7084 => x"00",
          7085 => x"00",
          7086 => x"00",
          7087 => x"00",
          7088 => x"00",
          7089 => x"00",
          7090 => x"00",
          7091 => x"00",
          7092 => x"64",
          7093 => x"2f",
          7094 => x"25",
          7095 => x"64",
          7096 => x"2e",
          7097 => x"64",
          7098 => x"6f",
          7099 => x"6f",
          7100 => x"67",
          7101 => x"74",
          7102 => x"00",
          7103 => x"28",
          7104 => x"6d",
          7105 => x"43",
          7106 => x"6e",
          7107 => x"29",
          7108 => x"0a",
          7109 => x"69",
          7110 => x"20",
          7111 => x"6c",
          7112 => x"6e",
          7113 => x"3a",
          7114 => x"20",
          7115 => x"42",
          7116 => x"52",
          7117 => x"20",
          7118 => x"38",
          7119 => x"30",
          7120 => x"2e",
          7121 => x"20",
          7122 => x"44",
          7123 => x"20",
          7124 => x"20",
          7125 => x"38",
          7126 => x"30",
          7127 => x"2e",
          7128 => x"20",
          7129 => x"4e",
          7130 => x"42",
          7131 => x"20",
          7132 => x"38",
          7133 => x"30",
          7134 => x"2e",
          7135 => x"20",
          7136 => x"52",
          7137 => x"20",
          7138 => x"20",
          7139 => x"38",
          7140 => x"30",
          7141 => x"2e",
          7142 => x"20",
          7143 => x"41",
          7144 => x"20",
          7145 => x"20",
          7146 => x"38",
          7147 => x"30",
          7148 => x"2e",
          7149 => x"20",
          7150 => x"44",
          7151 => x"52",
          7152 => x"20",
          7153 => x"76",
          7154 => x"73",
          7155 => x"30",
          7156 => x"2e",
          7157 => x"20",
          7158 => x"49",
          7159 => x"31",
          7160 => x"20",
          7161 => x"6d",
          7162 => x"20",
          7163 => x"30",
          7164 => x"2e",
          7165 => x"20",
          7166 => x"4e",
          7167 => x"43",
          7168 => x"20",
          7169 => x"61",
          7170 => x"6c",
          7171 => x"30",
          7172 => x"2e",
          7173 => x"20",
          7174 => x"49",
          7175 => x"4f",
          7176 => x"42",
          7177 => x"00",
          7178 => x"20",
          7179 => x"42",
          7180 => x"43",
          7181 => x"20",
          7182 => x"4f",
          7183 => x"0a",
          7184 => x"20",
          7185 => x"53",
          7186 => x"00",
          7187 => x"20",
          7188 => x"50",
          7189 => x"00",
          7190 => x"64",
          7191 => x"73",
          7192 => x"3a",
          7193 => x"20",
          7194 => x"50",
          7195 => x"65",
          7196 => x"20",
          7197 => x"74",
          7198 => x"41",
          7199 => x"65",
          7200 => x"3d",
          7201 => x"38",
          7202 => x"00",
          7203 => x"20",
          7204 => x"50",
          7205 => x"65",
          7206 => x"79",
          7207 => x"61",
          7208 => x"41",
          7209 => x"65",
          7210 => x"3d",
          7211 => x"38",
          7212 => x"00",
          7213 => x"20",
          7214 => x"74",
          7215 => x"20",
          7216 => x"72",
          7217 => x"64",
          7218 => x"73",
          7219 => x"20",
          7220 => x"3d",
          7221 => x"38",
          7222 => x"00",
          7223 => x"69",
          7224 => x"0a",
          7225 => x"20",
          7226 => x"50",
          7227 => x"64",
          7228 => x"20",
          7229 => x"20",
          7230 => x"20",
          7231 => x"20",
          7232 => x"3d",
          7233 => x"34",
          7234 => x"00",
          7235 => x"20",
          7236 => x"79",
          7237 => x"6d",
          7238 => x"6f",
          7239 => x"46",
          7240 => x"20",
          7241 => x"20",
          7242 => x"3d",
          7243 => x"2e",
          7244 => x"64",
          7245 => x"0a",
          7246 => x"20",
          7247 => x"44",
          7248 => x"20",
          7249 => x"63",
          7250 => x"72",
          7251 => x"20",
          7252 => x"20",
          7253 => x"3d",
          7254 => x"2e",
          7255 => x"64",
          7256 => x"0a",
          7257 => x"20",
          7258 => x"69",
          7259 => x"6f",
          7260 => x"53",
          7261 => x"4d",
          7262 => x"6f",
          7263 => x"46",
          7264 => x"3d",
          7265 => x"2e",
          7266 => x"64",
          7267 => x"0a",
          7268 => x"6d",
          7269 => x"00",
          7270 => x"65",
          7271 => x"6d",
          7272 => x"6c",
          7273 => x"00",
          7274 => x"56",
          7275 => x"56",
          7276 => x"6e",
          7277 => x"6e",
          7278 => x"77",
          7279 => x"69",
          7280 => x"72",
          7281 => x"78",
          7282 => x"69",
          7283 => x"72",
          7284 => x"69",
          7285 => x"00",
          7286 => x"00",
          7287 => x"30",
          7288 => x"20",
          7289 => x"00",
          7290 => x"61",
          7291 => x"64",
          7292 => x"20",
          7293 => x"65",
          7294 => x"68",
          7295 => x"69",
          7296 => x"72",
          7297 => x"69",
          7298 => x"74",
          7299 => x"4f",
          7300 => x"00",
          7301 => x"61",
          7302 => x"74",
          7303 => x"65",
          7304 => x"72",
          7305 => x"65",
          7306 => x"73",
          7307 => x"79",
          7308 => x"6c",
          7309 => x"64",
          7310 => x"62",
          7311 => x"67",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"5b",
          7347 => x"5b",
          7348 => x"5b",
          7349 => x"5b",
          7350 => x"5b",
          7351 => x"5b",
          7352 => x"5b",
          7353 => x"5b",
          7354 => x"5b",
          7355 => x"00",
          7356 => x"00",
          7357 => x"44",
          7358 => x"2a",
          7359 => x"3b",
          7360 => x"3f",
          7361 => x"7f",
          7362 => x"41",
          7363 => x"41",
          7364 => x"00",
          7365 => x"fe",
          7366 => x"44",
          7367 => x"2e",
          7368 => x"4f",
          7369 => x"4d",
          7370 => x"20",
          7371 => x"54",
          7372 => x"20",
          7373 => x"4f",
          7374 => x"4d",
          7375 => x"20",
          7376 => x"54",
          7377 => x"20",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"9a",
          7383 => x"41",
          7384 => x"45",
          7385 => x"49",
          7386 => x"92",
          7387 => x"4f",
          7388 => x"99",
          7389 => x"9d",
          7390 => x"49",
          7391 => x"a5",
          7392 => x"a9",
          7393 => x"ad",
          7394 => x"b1",
          7395 => x"b5",
          7396 => x"b9",
          7397 => x"bd",
          7398 => x"c1",
          7399 => x"c5",
          7400 => x"c9",
          7401 => x"cd",
          7402 => x"d1",
          7403 => x"d5",
          7404 => x"d9",
          7405 => x"dd",
          7406 => x"e1",
          7407 => x"e5",
          7408 => x"e9",
          7409 => x"ed",
          7410 => x"f1",
          7411 => x"f5",
          7412 => x"f9",
          7413 => x"fd",
          7414 => x"2e",
          7415 => x"5b",
          7416 => x"22",
          7417 => x"3e",
          7418 => x"00",
          7419 => x"01",
          7420 => x"10",
          7421 => x"00",
          7422 => x"00",
          7423 => x"01",
          7424 => x"04",
          7425 => x"10",
          7426 => x"00",
          7427 => x"69",
          7428 => x"00",
          7429 => x"69",
          7430 => x"6c",
          7431 => x"69",
          7432 => x"00",
          7433 => x"6c",
          7434 => x"00",
          7435 => x"65",
          7436 => x"00",
          7437 => x"63",
          7438 => x"72",
          7439 => x"63",
          7440 => x"00",
          7441 => x"64",
          7442 => x"00",
          7443 => x"64",
          7444 => x"00",
          7445 => x"65",
          7446 => x"65",
          7447 => x"65",
          7448 => x"69",
          7449 => x"69",
          7450 => x"66",
          7451 => x"66",
          7452 => x"61",
          7453 => x"00",
          7454 => x"6d",
          7455 => x"65",
          7456 => x"72",
          7457 => x"65",
          7458 => x"00",
          7459 => x"6e",
          7460 => x"00",
          7461 => x"65",
          7462 => x"00",
          7463 => x"62",
          7464 => x"63",
          7465 => x"62",
          7466 => x"63",
          7467 => x"69",
          7468 => x"00",
          7469 => x"69",
          7470 => x"45",
          7471 => x"72",
          7472 => x"6e",
          7473 => x"6e",
          7474 => x"65",
          7475 => x"72",
          7476 => x"00",
          7477 => x"69",
          7478 => x"6e",
          7479 => x"72",
          7480 => x"79",
          7481 => x"00",
          7482 => x"6f",
          7483 => x"6c",
          7484 => x"6f",
          7485 => x"2e",
          7486 => x"6f",
          7487 => x"74",
          7488 => x"6f",
          7489 => x"2e",
          7490 => x"6e",
          7491 => x"69",
          7492 => x"69",
          7493 => x"61",
          7494 => x"0a",
          7495 => x"63",
          7496 => x"73",
          7497 => x"6e",
          7498 => x"2e",
          7499 => x"69",
          7500 => x"61",
          7501 => x"61",
          7502 => x"65",
          7503 => x"74",
          7504 => x"00",
          7505 => x"69",
          7506 => x"68",
          7507 => x"6c",
          7508 => x"6e",
          7509 => x"69",
          7510 => x"00",
          7511 => x"44",
          7512 => x"20",
          7513 => x"74",
          7514 => x"72",
          7515 => x"63",
          7516 => x"2e",
          7517 => x"72",
          7518 => x"20",
          7519 => x"62",
          7520 => x"69",
          7521 => x"6e",
          7522 => x"69",
          7523 => x"00",
          7524 => x"69",
          7525 => x"6e",
          7526 => x"65",
          7527 => x"6c",
          7528 => x"0a",
          7529 => x"6f",
          7530 => x"6d",
          7531 => x"69",
          7532 => x"20",
          7533 => x"65",
          7534 => x"74",
          7535 => x"66",
          7536 => x"64",
          7537 => x"20",
          7538 => x"6b",
          7539 => x"00",
          7540 => x"6f",
          7541 => x"74",
          7542 => x"6f",
          7543 => x"64",
          7544 => x"00",
          7545 => x"69",
          7546 => x"75",
          7547 => x"6f",
          7548 => x"61",
          7549 => x"6e",
          7550 => x"6e",
          7551 => x"6c",
          7552 => x"0a",
          7553 => x"69",
          7554 => x"69",
          7555 => x"6f",
          7556 => x"64",
          7557 => x"00",
          7558 => x"6e",
          7559 => x"66",
          7560 => x"65",
          7561 => x"6d",
          7562 => x"72",
          7563 => x"00",
          7564 => x"6f",
          7565 => x"61",
          7566 => x"6f",
          7567 => x"20",
          7568 => x"65",
          7569 => x"00",
          7570 => x"61",
          7571 => x"65",
          7572 => x"73",
          7573 => x"63",
          7574 => x"65",
          7575 => x"0a",
          7576 => x"75",
          7577 => x"73",
          7578 => x"00",
          7579 => x"6e",
          7580 => x"77",
          7581 => x"72",
          7582 => x"2e",
          7583 => x"25",
          7584 => x"62",
          7585 => x"73",
          7586 => x"20",
          7587 => x"25",
          7588 => x"62",
          7589 => x"73",
          7590 => x"63",
          7591 => x"00",
          7592 => x"65",
          7593 => x"00",
          7594 => x"30",
          7595 => x"00",
          7596 => x"20",
          7597 => x"30",
          7598 => x"00",
          7599 => x"20",
          7600 => x"20",
          7601 => x"00",
          7602 => x"30",
          7603 => x"00",
          7604 => x"20",
          7605 => x"7c",
          7606 => x"0d",
          7607 => x"4f",
          7608 => x"2a",
          7609 => x"73",
          7610 => x"00",
          7611 => x"37",
          7612 => x"2f",
          7613 => x"30",
          7614 => x"31",
          7615 => x"00",
          7616 => x"5a",
          7617 => x"20",
          7618 => x"20",
          7619 => x"78",
          7620 => x"73",
          7621 => x"20",
          7622 => x"0a",
          7623 => x"50",
          7624 => x"6e",
          7625 => x"72",
          7626 => x"20",
          7627 => x"64",
          7628 => x"0a",
          7629 => x"69",
          7630 => x"20",
          7631 => x"65",
          7632 => x"70",
          7633 => x"00",
          7634 => x"53",
          7635 => x"6e",
          7636 => x"72",
          7637 => x"0a",
          7638 => x"4f",
          7639 => x"20",
          7640 => x"69",
          7641 => x"72",
          7642 => x"74",
          7643 => x"4f",
          7644 => x"20",
          7645 => x"69",
          7646 => x"72",
          7647 => x"74",
          7648 => x"41",
          7649 => x"20",
          7650 => x"69",
          7651 => x"72",
          7652 => x"74",
          7653 => x"41",
          7654 => x"20",
          7655 => x"69",
          7656 => x"72",
          7657 => x"74",
          7658 => x"41",
          7659 => x"20",
          7660 => x"69",
          7661 => x"72",
          7662 => x"74",
          7663 => x"41",
          7664 => x"20",
          7665 => x"69",
          7666 => x"72",
          7667 => x"74",
          7668 => x"65",
          7669 => x"6e",
          7670 => x"70",
          7671 => x"6d",
          7672 => x"2e",
          7673 => x"00",
          7674 => x"6e",
          7675 => x"69",
          7676 => x"74",
          7677 => x"72",
          7678 => x"0a",
          7679 => x"75",
          7680 => x"78",
          7681 => x"62",
          7682 => x"00",
          7683 => x"3a",
          7684 => x"61",
          7685 => x"64",
          7686 => x"20",
          7687 => x"74",
          7688 => x"69",
          7689 => x"73",
          7690 => x"61",
          7691 => x"30",
          7692 => x"6c",
          7693 => x"65",
          7694 => x"69",
          7695 => x"61",
          7696 => x"6c",
          7697 => x"0a",
          7698 => x"20",
          7699 => x"6c",
          7700 => x"69",
          7701 => x"2e",
          7702 => x"00",
          7703 => x"6f",
          7704 => x"6e",
          7705 => x"2e",
          7706 => x"6f",
          7707 => x"72",
          7708 => x"2e",
          7709 => x"00",
          7710 => x"30",
          7711 => x"28",
          7712 => x"78",
          7713 => x"25",
          7714 => x"78",
          7715 => x"38",
          7716 => x"00",
          7717 => x"75",
          7718 => x"4d",
          7719 => x"72",
          7720 => x"00",
          7721 => x"43",
          7722 => x"6c",
          7723 => x"2e",
          7724 => x"30",
          7725 => x"25",
          7726 => x"2d",
          7727 => x"3f",
          7728 => x"00",
          7729 => x"30",
          7730 => x"25",
          7731 => x"2d",
          7732 => x"30",
          7733 => x"25",
          7734 => x"2d",
          7735 => x"78",
          7736 => x"74",
          7737 => x"20",
          7738 => x"65",
          7739 => x"25",
          7740 => x"20",
          7741 => x"0a",
          7742 => x"61",
          7743 => x"6e",
          7744 => x"6f",
          7745 => x"40",
          7746 => x"38",
          7747 => x"2e",
          7748 => x"00",
          7749 => x"61",
          7750 => x"72",
          7751 => x"72",
          7752 => x"20",
          7753 => x"65",
          7754 => x"64",
          7755 => x"00",
          7756 => x"65",
          7757 => x"72",
          7758 => x"67",
          7759 => x"70",
          7760 => x"61",
          7761 => x"6e",
          7762 => x"0a",
          7763 => x"6f",
          7764 => x"72",
          7765 => x"6f",
          7766 => x"67",
          7767 => x"0a",
          7768 => x"50",
          7769 => x"69",
          7770 => x"64",
          7771 => x"73",
          7772 => x"2e",
          7773 => x"00",
          7774 => x"64",
          7775 => x"73",
          7776 => x"00",
          7777 => x"64",
          7778 => x"73",
          7779 => x"61",
          7780 => x"6f",
          7781 => x"6e",
          7782 => x"00",
          7783 => x"75",
          7784 => x"6e",
          7785 => x"2e",
          7786 => x"6e",
          7787 => x"69",
          7788 => x"69",
          7789 => x"72",
          7790 => x"74",
          7791 => x"2e",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"01",
          7798 => x"00",
          7799 => x"01",
          7800 => x"81",
          7801 => x"00",
          7802 => x"7f",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"f5",
          7808 => x"f5",
          7809 => x"f5",
          7810 => x"00",
          7811 => x"01",
          7812 => x"01",
          7813 => x"01",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"00",
          7848 => x"00",
          7849 => x"00",
          7850 => x"00",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"00",
          7855 => x"02",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"04",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"14",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"2b",
          7868 => x"00",
          7869 => x"00",
          7870 => x"00",
          7871 => x"30",
          7872 => x"00",
          7873 => x"00",
          7874 => x"00",
          7875 => x"3c",
          7876 => x"00",
          7877 => x"00",
          7878 => x"00",
          7879 => x"3d",
          7880 => x"00",
          7881 => x"00",
          7882 => x"00",
          7883 => x"3f",
          7884 => x"00",
          7885 => x"00",
          7886 => x"00",
          7887 => x"40",
          7888 => x"00",
          7889 => x"00",
          7890 => x"00",
          7891 => x"41",
          7892 => x"00",
          7893 => x"00",
          7894 => x"00",
          7895 => x"42",
          7896 => x"00",
          7897 => x"00",
          7898 => x"00",
          7899 => x"43",
          7900 => x"00",
          7901 => x"00",
          7902 => x"00",
          7903 => x"50",
          7904 => x"00",
          7905 => x"00",
          7906 => x"00",
          7907 => x"51",
          7908 => x"00",
          7909 => x"00",
          7910 => x"00",
          7911 => x"54",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"55",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"79",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"78",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"82",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"83",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"85",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"87",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"8c",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"8d",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"8e",
          7952 => x"00",
          7953 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"8c",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"f0",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"ac",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"91",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"fd",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b2",
           272 => x"0b",
           273 => x"0b",
           274 => x"d0",
           275 => x"0b",
           276 => x"0b",
           277 => x"ee",
           278 => x"0b",
           279 => x"0b",
           280 => x"8c",
           281 => x"0b",
           282 => x"0b",
           283 => x"aa",
           284 => x"0b",
           285 => x"0b",
           286 => x"c8",
           287 => x"0b",
           288 => x"0b",
           289 => x"e6",
           290 => x"0b",
           291 => x"0b",
           292 => x"84",
           293 => x"0b",
           294 => x"0b",
           295 => x"a3",
           296 => x"0b",
           297 => x"0b",
           298 => x"c3",
           299 => x"0b",
           300 => x"0b",
           301 => x"e3",
           302 => x"0b",
           303 => x"0b",
           304 => x"83",
           305 => x"0b",
           306 => x"0b",
           307 => x"a3",
           308 => x"0b",
           309 => x"0b",
           310 => x"c3",
           311 => x"0b",
           312 => x"0b",
           313 => x"e3",
           314 => x"0b",
           315 => x"0b",
           316 => x"83",
           317 => x"0b",
           318 => x"0b",
           319 => x"a3",
           320 => x"0b",
           321 => x"0b",
           322 => x"c3",
           323 => x"0b",
           324 => x"0b",
           325 => x"e3",
           326 => x"0b",
           327 => x"0b",
           328 => x"83",
           329 => x"0b",
           330 => x"0b",
           331 => x"a3",
           332 => x"0b",
           333 => x"0b",
           334 => x"c3",
           335 => x"0b",
           336 => x"0b",
           337 => x"e3",
           338 => x"0b",
           339 => x"0b",
           340 => x"82",
           341 => x"0b",
           342 => x"0b",
           343 => x"a0",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"81",
           388 => x"83",
           389 => x"81",
           390 => x"b5",
           391 => x"f8",
           392 => x"80",
           393 => x"f8",
           394 => x"c6",
           395 => x"d4",
           396 => x"90",
           397 => x"d4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"81",
           403 => x"83",
           404 => x"81",
           405 => x"bd",
           406 => x"f8",
           407 => x"80",
           408 => x"f8",
           409 => x"87",
           410 => x"d4",
           411 => x"90",
           412 => x"d4",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"81",
           418 => x"83",
           419 => x"81",
           420 => x"bb",
           421 => x"f8",
           422 => x"80",
           423 => x"f8",
           424 => x"b9",
           425 => x"d4",
           426 => x"90",
           427 => x"d4",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"81",
           433 => x"83",
           434 => x"81",
           435 => x"a6",
           436 => x"f8",
           437 => x"80",
           438 => x"f8",
           439 => x"dd",
           440 => x"d4",
           441 => x"90",
           442 => x"d4",
           443 => x"2d",
           444 => x"08",
           445 => x"04",
           446 => x"0c",
           447 => x"81",
           448 => x"83",
           449 => x"81",
           450 => x"a1",
           451 => x"f8",
           452 => x"80",
           453 => x"f8",
           454 => x"84",
           455 => x"f8",
           456 => x"80",
           457 => x"f8",
           458 => x"90",
           459 => x"f8",
           460 => x"80",
           461 => x"f8",
           462 => x"88",
           463 => x"f8",
           464 => x"80",
           465 => x"f8",
           466 => x"8b",
           467 => x"f8",
           468 => x"80",
           469 => x"f8",
           470 => x"96",
           471 => x"f8",
           472 => x"80",
           473 => x"f8",
           474 => x"9e",
           475 => x"f8",
           476 => x"80",
           477 => x"f8",
           478 => x"8f",
           479 => x"f8",
           480 => x"80",
           481 => x"f8",
           482 => x"99",
           483 => x"f8",
           484 => x"80",
           485 => x"f8",
           486 => x"9a",
           487 => x"f8",
           488 => x"80",
           489 => x"f8",
           490 => x"9a",
           491 => x"f8",
           492 => x"80",
           493 => x"f8",
           494 => x"a2",
           495 => x"f8",
           496 => x"80",
           497 => x"f8",
           498 => x"a0",
           499 => x"f8",
           500 => x"80",
           501 => x"f8",
           502 => x"a5",
           503 => x"f8",
           504 => x"80",
           505 => x"f8",
           506 => x"9b",
           507 => x"f8",
           508 => x"80",
           509 => x"f8",
           510 => x"a8",
           511 => x"f8",
           512 => x"80",
           513 => x"f8",
           514 => x"a9",
           515 => x"f8",
           516 => x"80",
           517 => x"f8",
           518 => x"91",
           519 => x"f8",
           520 => x"80",
           521 => x"f8",
           522 => x"91",
           523 => x"f8",
           524 => x"80",
           525 => x"f8",
           526 => x"92",
           527 => x"f8",
           528 => x"80",
           529 => x"f8",
           530 => x"9c",
           531 => x"f8",
           532 => x"80",
           533 => x"f8",
           534 => x"aa",
           535 => x"f8",
           536 => x"80",
           537 => x"f8",
           538 => x"ac",
           539 => x"f8",
           540 => x"80",
           541 => x"f8",
           542 => x"af",
           543 => x"f8",
           544 => x"80",
           545 => x"f8",
           546 => x"83",
           547 => x"f8",
           548 => x"80",
           549 => x"f8",
           550 => x"b2",
           551 => x"f8",
           552 => x"80",
           553 => x"f8",
           554 => x"c0",
           555 => x"f8",
           556 => x"80",
           557 => x"f8",
           558 => x"be",
           559 => x"f8",
           560 => x"80",
           561 => x"f8",
           562 => x"d4",
           563 => x"f8",
           564 => x"80",
           565 => x"f8",
           566 => x"d6",
           567 => x"f8",
           568 => x"80",
           569 => x"f8",
           570 => x"d8",
           571 => x"f8",
           572 => x"80",
           573 => x"f8",
           574 => x"a2",
           575 => x"d4",
           576 => x"90",
           577 => x"d4",
           578 => x"2d",
           579 => x"08",
           580 => x"04",
           581 => x"0c",
           582 => x"81",
           583 => x"83",
           584 => x"81",
           585 => x"81",
           586 => x"81",
           587 => x"83",
           588 => x"3c",
           589 => x"10",
           590 => x"10",
           591 => x"10",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"51",
           598 => x"73",
           599 => x"73",
           600 => x"81",
           601 => x"10",
           602 => x"07",
           603 => x"0c",
           604 => x"72",
           605 => x"81",
           606 => x"09",
           607 => x"71",
           608 => x"0a",
           609 => x"72",
           610 => x"51",
           611 => x"81",
           612 => x"82",
           613 => x"8e",
           614 => x"70",
           615 => x"0c",
           616 => x"93",
           617 => x"81",
           618 => x"fd",
           619 => x"f8",
           620 => x"81",
           621 => x"fd",
           622 => x"53",
           623 => x"08",
           624 => x"52",
           625 => x"08",
           626 => x"51",
           627 => x"81",
           628 => x"70",
           629 => x"0c",
           630 => x"0d",
           631 => x"0c",
           632 => x"d4",
           633 => x"f8",
           634 => x"3d",
           635 => x"81",
           636 => x"8c",
           637 => x"81",
           638 => x"88",
           639 => x"83",
           640 => x"f8",
           641 => x"81",
           642 => x"54",
           643 => x"81",
           644 => x"04",
           645 => x"08",
           646 => x"d4",
           647 => x"0d",
           648 => x"f8",
           649 => x"05",
           650 => x"d4",
           651 => x"08",
           652 => x"38",
           653 => x"08",
           654 => x"30",
           655 => x"08",
           656 => x"80",
           657 => x"d4",
           658 => x"0c",
           659 => x"08",
           660 => x"8a",
           661 => x"81",
           662 => x"f4",
           663 => x"f8",
           664 => x"05",
           665 => x"d4",
           666 => x"0c",
           667 => x"08",
           668 => x"80",
           669 => x"81",
           670 => x"8c",
           671 => x"81",
           672 => x"8c",
           673 => x"0b",
           674 => x"08",
           675 => x"81",
           676 => x"fc",
           677 => x"38",
           678 => x"f8",
           679 => x"05",
           680 => x"d4",
           681 => x"08",
           682 => x"08",
           683 => x"80",
           684 => x"d4",
           685 => x"08",
           686 => x"d4",
           687 => x"08",
           688 => x"3f",
           689 => x"08",
           690 => x"d4",
           691 => x"0c",
           692 => x"d4",
           693 => x"08",
           694 => x"38",
           695 => x"08",
           696 => x"30",
           697 => x"08",
           698 => x"81",
           699 => x"f8",
           700 => x"81",
           701 => x"54",
           702 => x"81",
           703 => x"04",
           704 => x"08",
           705 => x"d4",
           706 => x"0d",
           707 => x"f8",
           708 => x"05",
           709 => x"d4",
           710 => x"08",
           711 => x"38",
           712 => x"08",
           713 => x"30",
           714 => x"08",
           715 => x"81",
           716 => x"d4",
           717 => x"0c",
           718 => x"08",
           719 => x"80",
           720 => x"81",
           721 => x"8c",
           722 => x"81",
           723 => x"8c",
           724 => x"53",
           725 => x"08",
           726 => x"52",
           727 => x"08",
           728 => x"51",
           729 => x"f8",
           730 => x"81",
           731 => x"f8",
           732 => x"81",
           733 => x"fc",
           734 => x"2e",
           735 => x"f8",
           736 => x"05",
           737 => x"f8",
           738 => x"05",
           739 => x"d4",
           740 => x"08",
           741 => x"c8",
           742 => x"3d",
           743 => x"d4",
           744 => x"f8",
           745 => x"81",
           746 => x"fd",
           747 => x"0b",
           748 => x"08",
           749 => x"80",
           750 => x"d4",
           751 => x"0c",
           752 => x"08",
           753 => x"81",
           754 => x"88",
           755 => x"b9",
           756 => x"d4",
           757 => x"08",
           758 => x"38",
           759 => x"f8",
           760 => x"05",
           761 => x"38",
           762 => x"08",
           763 => x"10",
           764 => x"08",
           765 => x"81",
           766 => x"fc",
           767 => x"81",
           768 => x"fc",
           769 => x"b8",
           770 => x"d4",
           771 => x"08",
           772 => x"e1",
           773 => x"d4",
           774 => x"08",
           775 => x"08",
           776 => x"26",
           777 => x"f8",
           778 => x"05",
           779 => x"d4",
           780 => x"08",
           781 => x"d4",
           782 => x"0c",
           783 => x"08",
           784 => x"81",
           785 => x"fc",
           786 => x"81",
           787 => x"f8",
           788 => x"f8",
           789 => x"05",
           790 => x"81",
           791 => x"fc",
           792 => x"f8",
           793 => x"05",
           794 => x"81",
           795 => x"8c",
           796 => x"95",
           797 => x"d4",
           798 => x"08",
           799 => x"38",
           800 => x"08",
           801 => x"70",
           802 => x"08",
           803 => x"51",
           804 => x"f8",
           805 => x"05",
           806 => x"f8",
           807 => x"05",
           808 => x"f8",
           809 => x"05",
           810 => x"c8",
           811 => x"0d",
           812 => x"0c",
           813 => x"0d",
           814 => x"7b",
           815 => x"55",
           816 => x"8c",
           817 => x"07",
           818 => x"70",
           819 => x"38",
           820 => x"71",
           821 => x"38",
           822 => x"05",
           823 => x"70",
           824 => x"34",
           825 => x"71",
           826 => x"81",
           827 => x"74",
           828 => x"0c",
           829 => x"04",
           830 => x"70",
           831 => x"08",
           832 => x"05",
           833 => x"70",
           834 => x"08",
           835 => x"05",
           836 => x"70",
           837 => x"08",
           838 => x"05",
           839 => x"70",
           840 => x"08",
           841 => x"05",
           842 => x"12",
           843 => x"26",
           844 => x"72",
           845 => x"72",
           846 => x"54",
           847 => x"84",
           848 => x"fc",
           849 => x"83",
           850 => x"70",
           851 => x"39",
           852 => x"76",
           853 => x"8c",
           854 => x"33",
           855 => x"55",
           856 => x"8a",
           857 => x"06",
           858 => x"2e",
           859 => x"12",
           860 => x"2e",
           861 => x"73",
           862 => x"55",
           863 => x"52",
           864 => x"09",
           865 => x"38",
           866 => x"c8",
           867 => x"0d",
           868 => x"88",
           869 => x"70",
           870 => x"07",
           871 => x"8f",
           872 => x"38",
           873 => x"84",
           874 => x"72",
           875 => x"05",
           876 => x"71",
           877 => x"53",
           878 => x"70",
           879 => x"0c",
           880 => x"71",
           881 => x"38",
           882 => x"90",
           883 => x"70",
           884 => x"0c",
           885 => x"71",
           886 => x"38",
           887 => x"8e",
           888 => x"0d",
           889 => x"70",
           890 => x"06",
           891 => x"55",
           892 => x"38",
           893 => x"70",
           894 => x"fb",
           895 => x"06",
           896 => x"82",
           897 => x"51",
           898 => x"54",
           899 => x"84",
           900 => x"70",
           901 => x"0c",
           902 => x"09",
           903 => x"fd",
           904 => x"70",
           905 => x"81",
           906 => x"51",
           907 => x"70",
           908 => x"38",
           909 => x"70",
           910 => x"33",
           911 => x"70",
           912 => x"34",
           913 => x"74",
           914 => x"0c",
           915 => x"04",
           916 => x"75",
           917 => x"06",
           918 => x"70",
           919 => x"70",
           920 => x"f7",
           921 => x"12",
           922 => x"84",
           923 => x"06",
           924 => x"53",
           925 => x"84",
           926 => x"70",
           927 => x"fd",
           928 => x"70",
           929 => x"81",
           930 => x"51",
           931 => x"80",
           932 => x"72",
           933 => x"51",
           934 => x"8a",
           935 => x"70",
           936 => x"70",
           937 => x"74",
           938 => x"c8",
           939 => x"0d",
           940 => x"0d",
           941 => x"70",
           942 => x"52",
           943 => x"80",
           944 => x"74",
           945 => x"51",
           946 => x"80",
           947 => x"13",
           948 => x"2e",
           949 => x"33",
           950 => x"51",
           951 => x"09",
           952 => x"38",
           953 => x"81",
           954 => x"81",
           955 => x"70",
           956 => x"fe",
           957 => x"81",
           958 => x"55",
           959 => x"ff",
           960 => x"06",
           961 => x"33",
           962 => x"51",
           963 => x"06",
           964 => x"06",
           965 => x"51",
           966 => x"81",
           967 => x"88",
           968 => x"71",
           969 => x"83",
           970 => x"38",
           971 => x"08",
           972 => x"74",
           973 => x"ff",
           974 => x"13",
           975 => x"2e",
           976 => x"08",
           977 => x"fb",
           978 => x"06",
           979 => x"82",
           980 => x"51",
           981 => x"9a",
           982 => x"84",
           983 => x"83",
           984 => x"38",
           985 => x"08",
           986 => x"74",
           987 => x"fe",
           988 => x"0b",
           989 => x"0c",
           990 => x"04",
           991 => x"80",
           992 => x"71",
           993 => x"87",
           994 => x"f8",
           995 => x"ff",
           996 => x"ff",
           997 => x"72",
           998 => x"38",
           999 => x"c8",
          1000 => x"0d",
          1001 => x"0d",
          1002 => x"70",
          1003 => x"71",
          1004 => x"ca",
          1005 => x"51",
          1006 => x"09",
          1007 => x"38",
          1008 => x"f1",
          1009 => x"84",
          1010 => x"53",
          1011 => x"70",
          1012 => x"53",
          1013 => x"a0",
          1014 => x"81",
          1015 => x"2e",
          1016 => x"e5",
          1017 => x"ff",
          1018 => x"a0",
          1019 => x"06",
          1020 => x"73",
          1021 => x"55",
          1022 => x"0c",
          1023 => x"81",
          1024 => x"87",
          1025 => x"fc",
          1026 => x"53",
          1027 => x"2e",
          1028 => x"3d",
          1029 => x"72",
          1030 => x"3f",
          1031 => x"08",
          1032 => x"53",
          1033 => x"53",
          1034 => x"c8",
          1035 => x"0d",
          1036 => x"0d",
          1037 => x"33",
          1038 => x"53",
          1039 => x"8b",
          1040 => x"38",
          1041 => x"ff",
          1042 => x"52",
          1043 => x"81",
          1044 => x"13",
          1045 => x"52",
          1046 => x"80",
          1047 => x"13",
          1048 => x"52",
          1049 => x"80",
          1050 => x"13",
          1051 => x"52",
          1052 => x"80",
          1053 => x"13",
          1054 => x"52",
          1055 => x"26",
          1056 => x"8a",
          1057 => x"87",
          1058 => x"e7",
          1059 => x"38",
          1060 => x"c0",
          1061 => x"72",
          1062 => x"98",
          1063 => x"13",
          1064 => x"98",
          1065 => x"13",
          1066 => x"98",
          1067 => x"13",
          1068 => x"98",
          1069 => x"13",
          1070 => x"98",
          1071 => x"13",
          1072 => x"98",
          1073 => x"87",
          1074 => x"0c",
          1075 => x"98",
          1076 => x"0b",
          1077 => x"9c",
          1078 => x"71",
          1079 => x"0c",
          1080 => x"04",
          1081 => x"7f",
          1082 => x"98",
          1083 => x"7d",
          1084 => x"98",
          1085 => x"7d",
          1086 => x"c0",
          1087 => x"5a",
          1088 => x"34",
          1089 => x"b4",
          1090 => x"83",
          1091 => x"c0",
          1092 => x"5a",
          1093 => x"34",
          1094 => x"ac",
          1095 => x"85",
          1096 => x"c0",
          1097 => x"5a",
          1098 => x"34",
          1099 => x"a4",
          1100 => x"88",
          1101 => x"c0",
          1102 => x"5a",
          1103 => x"23",
          1104 => x"79",
          1105 => x"06",
          1106 => x"ff",
          1107 => x"86",
          1108 => x"85",
          1109 => x"84",
          1110 => x"83",
          1111 => x"82",
          1112 => x"7d",
          1113 => x"06",
          1114 => x"d0",
          1115 => x"3f",
          1116 => x"04",
          1117 => x"02",
          1118 => x"70",
          1119 => x"2a",
          1120 => x"70",
          1121 => x"f3",
          1122 => x"3d",
          1123 => x"3d",
          1124 => x"0b",
          1125 => x"33",
          1126 => x"06",
          1127 => x"87",
          1128 => x"51",
          1129 => x"86",
          1130 => x"94",
          1131 => x"08",
          1132 => x"70",
          1133 => x"54",
          1134 => x"2e",
          1135 => x"91",
          1136 => x"06",
          1137 => x"d7",
          1138 => x"32",
          1139 => x"51",
          1140 => x"2e",
          1141 => x"93",
          1142 => x"06",
          1143 => x"ff",
          1144 => x"81",
          1145 => x"87",
          1146 => x"52",
          1147 => x"86",
          1148 => x"94",
          1149 => x"72",
          1150 => x"f8",
          1151 => x"3d",
          1152 => x"3d",
          1153 => x"05",
          1154 => x"81",
          1155 => x"70",
          1156 => x"57",
          1157 => x"c0",
          1158 => x"74",
          1159 => x"38",
          1160 => x"94",
          1161 => x"70",
          1162 => x"81",
          1163 => x"52",
          1164 => x"8c",
          1165 => x"2a",
          1166 => x"51",
          1167 => x"38",
          1168 => x"70",
          1169 => x"51",
          1170 => x"8d",
          1171 => x"2a",
          1172 => x"51",
          1173 => x"be",
          1174 => x"ff",
          1175 => x"c0",
          1176 => x"70",
          1177 => x"38",
          1178 => x"90",
          1179 => x"0c",
          1180 => x"04",
          1181 => x"79",
          1182 => x"33",
          1183 => x"06",
          1184 => x"70",
          1185 => x"fe",
          1186 => x"ff",
          1187 => x"0b",
          1188 => x"c0",
          1189 => x"ff",
          1190 => x"55",
          1191 => x"94",
          1192 => x"80",
          1193 => x"87",
          1194 => x"51",
          1195 => x"96",
          1196 => x"06",
          1197 => x"70",
          1198 => x"38",
          1199 => x"70",
          1200 => x"51",
          1201 => x"72",
          1202 => x"81",
          1203 => x"70",
          1204 => x"38",
          1205 => x"70",
          1206 => x"51",
          1207 => x"38",
          1208 => x"06",
          1209 => x"94",
          1210 => x"80",
          1211 => x"87",
          1212 => x"52",
          1213 => x"81",
          1214 => x"70",
          1215 => x"53",
          1216 => x"ff",
          1217 => x"81",
          1218 => x"89",
          1219 => x"fe",
          1220 => x"0b",
          1221 => x"33",
          1222 => x"06",
          1223 => x"c0",
          1224 => x"72",
          1225 => x"38",
          1226 => x"94",
          1227 => x"70",
          1228 => x"81",
          1229 => x"51",
          1230 => x"e2",
          1231 => x"ff",
          1232 => x"c0",
          1233 => x"70",
          1234 => x"38",
          1235 => x"90",
          1236 => x"70",
          1237 => x"81",
          1238 => x"51",
          1239 => x"04",
          1240 => x"0b",
          1241 => x"c0",
          1242 => x"ff",
          1243 => x"87",
          1244 => x"52",
          1245 => x"86",
          1246 => x"94",
          1247 => x"08",
          1248 => x"70",
          1249 => x"51",
          1250 => x"70",
          1251 => x"38",
          1252 => x"06",
          1253 => x"94",
          1254 => x"80",
          1255 => x"87",
          1256 => x"52",
          1257 => x"98",
          1258 => x"2c",
          1259 => x"71",
          1260 => x"0c",
          1261 => x"04",
          1262 => x"87",
          1263 => x"08",
          1264 => x"8a",
          1265 => x"70",
          1266 => x"b4",
          1267 => x"9e",
          1268 => x"f3",
          1269 => x"c0",
          1270 => x"81",
          1271 => x"87",
          1272 => x"08",
          1273 => x"0c",
          1274 => x"98",
          1275 => x"d0",
          1276 => x"9e",
          1277 => x"f3",
          1278 => x"c0",
          1279 => x"81",
          1280 => x"87",
          1281 => x"08",
          1282 => x"0c",
          1283 => x"b0",
          1284 => x"e0",
          1285 => x"9e",
          1286 => x"f3",
          1287 => x"c0",
          1288 => x"81",
          1289 => x"87",
          1290 => x"08",
          1291 => x"0c",
          1292 => x"c0",
          1293 => x"f0",
          1294 => x"9e",
          1295 => x"f3",
          1296 => x"c0",
          1297 => x"51",
          1298 => x"f8",
          1299 => x"9e",
          1300 => x"f3",
          1301 => x"c0",
          1302 => x"81",
          1303 => x"87",
          1304 => x"08",
          1305 => x"0c",
          1306 => x"f4",
          1307 => x"0b",
          1308 => x"90",
          1309 => x"80",
          1310 => x"52",
          1311 => x"2e",
          1312 => x"52",
          1313 => x"89",
          1314 => x"87",
          1315 => x"08",
          1316 => x"0a",
          1317 => x"52",
          1318 => x"83",
          1319 => x"71",
          1320 => x"34",
          1321 => x"c0",
          1322 => x"70",
          1323 => x"06",
          1324 => x"70",
          1325 => x"38",
          1326 => x"81",
          1327 => x"80",
          1328 => x"9e",
          1329 => x"88",
          1330 => x"51",
          1331 => x"80",
          1332 => x"81",
          1333 => x"f4",
          1334 => x"0b",
          1335 => x"90",
          1336 => x"80",
          1337 => x"52",
          1338 => x"2e",
          1339 => x"52",
          1340 => x"8d",
          1341 => x"87",
          1342 => x"08",
          1343 => x"80",
          1344 => x"52",
          1345 => x"83",
          1346 => x"71",
          1347 => x"34",
          1348 => x"c0",
          1349 => x"70",
          1350 => x"06",
          1351 => x"70",
          1352 => x"38",
          1353 => x"81",
          1354 => x"80",
          1355 => x"9e",
          1356 => x"82",
          1357 => x"51",
          1358 => x"80",
          1359 => x"81",
          1360 => x"f4",
          1361 => x"0b",
          1362 => x"90",
          1363 => x"80",
          1364 => x"52",
          1365 => x"2e",
          1366 => x"52",
          1367 => x"91",
          1368 => x"87",
          1369 => x"08",
          1370 => x"80",
          1371 => x"52",
          1372 => x"83",
          1373 => x"71",
          1374 => x"34",
          1375 => x"c0",
          1376 => x"70",
          1377 => x"51",
          1378 => x"80",
          1379 => x"81",
          1380 => x"f4",
          1381 => x"c0",
          1382 => x"70",
          1383 => x"70",
          1384 => x"51",
          1385 => x"f4",
          1386 => x"0b",
          1387 => x"90",
          1388 => x"80",
          1389 => x"52",
          1390 => x"83",
          1391 => x"71",
          1392 => x"34",
          1393 => x"90",
          1394 => x"f0",
          1395 => x"2a",
          1396 => x"70",
          1397 => x"34",
          1398 => x"c0",
          1399 => x"70",
          1400 => x"52",
          1401 => x"2e",
          1402 => x"52",
          1403 => x"97",
          1404 => x"9e",
          1405 => x"87",
          1406 => x"70",
          1407 => x"34",
          1408 => x"04",
          1409 => x"81",
          1410 => x"89",
          1411 => x"f4",
          1412 => x"73",
          1413 => x"38",
          1414 => x"51",
          1415 => x"81",
          1416 => x"89",
          1417 => x"f4",
          1418 => x"73",
          1419 => x"38",
          1420 => x"08",
          1421 => x"08",
          1422 => x"81",
          1423 => x"8f",
          1424 => x"f4",
          1425 => x"73",
          1426 => x"38",
          1427 => x"08",
          1428 => x"08",
          1429 => x"81",
          1430 => x"8e",
          1431 => x"f4",
          1432 => x"73",
          1433 => x"38",
          1434 => x"08",
          1435 => x"08",
          1436 => x"81",
          1437 => x"8e",
          1438 => x"f4",
          1439 => x"73",
          1440 => x"38",
          1441 => x"08",
          1442 => x"08",
          1443 => x"81",
          1444 => x"8e",
          1445 => x"f4",
          1446 => x"73",
          1447 => x"38",
          1448 => x"08",
          1449 => x"08",
          1450 => x"81",
          1451 => x"8e",
          1452 => x"f4",
          1453 => x"73",
          1454 => x"38",
          1455 => x"33",
          1456 => x"b4",
          1457 => x"3f",
          1458 => x"33",
          1459 => x"2e",
          1460 => x"f4",
          1461 => x"81",
          1462 => x"8d",
          1463 => x"f4",
          1464 => x"73",
          1465 => x"38",
          1466 => x"33",
          1467 => x"f4",
          1468 => x"3f",
          1469 => x"33",
          1470 => x"2e",
          1471 => x"e0",
          1472 => x"e3",
          1473 => x"8b",
          1474 => x"80",
          1475 => x"81",
          1476 => x"87",
          1477 => x"f4",
          1478 => x"73",
          1479 => x"38",
          1480 => x"51",
          1481 => x"81",
          1482 => x"54",
          1483 => x"88",
          1484 => x"c0",
          1485 => x"3f",
          1486 => x"33",
          1487 => x"2e",
          1488 => x"e0",
          1489 => x"9f",
          1490 => x"d8",
          1491 => x"3f",
          1492 => x"08",
          1493 => x"e4",
          1494 => x"3f",
          1495 => x"08",
          1496 => x"8c",
          1497 => x"3f",
          1498 => x"08",
          1499 => x"b4",
          1500 => x"3f",
          1501 => x"51",
          1502 => x"81",
          1503 => x"52",
          1504 => x"51",
          1505 => x"81",
          1506 => x"56",
          1507 => x"52",
          1508 => x"9a",
          1509 => x"c8",
          1510 => x"c0",
          1511 => x"31",
          1512 => x"f8",
          1513 => x"81",
          1514 => x"8c",
          1515 => x"f4",
          1516 => x"73",
          1517 => x"38",
          1518 => x"08",
          1519 => x"c0",
          1520 => x"e3",
          1521 => x"f8",
          1522 => x"84",
          1523 => x"71",
          1524 => x"81",
          1525 => x"52",
          1526 => x"51",
          1527 => x"81",
          1528 => x"54",
          1529 => x"a8",
          1530 => x"84",
          1531 => x"84",
          1532 => x"51",
          1533 => x"81",
          1534 => x"bd",
          1535 => x"76",
          1536 => x"54",
          1537 => x"08",
          1538 => x"e4",
          1539 => x"3f",
          1540 => x"51",
          1541 => x"87",
          1542 => x"fe",
          1543 => x"92",
          1544 => x"05",
          1545 => x"26",
          1546 => x"84",
          1547 => x"bc",
          1548 => x"08",
          1549 => x"90",
          1550 => x"81",
          1551 => x"97",
          1552 => x"a0",
          1553 => x"81",
          1554 => x"8b",
          1555 => x"ac",
          1556 => x"81",
          1557 => x"85",
          1558 => x"3d",
          1559 => x"88",
          1560 => x"80",
          1561 => x"96",
          1562 => x"81",
          1563 => x"87",
          1564 => x"0c",
          1565 => x"0d",
          1566 => x"08",
          1567 => x"90",
          1568 => x"f8",
          1569 => x"f8",
          1570 => x"11",
          1571 => x"53",
          1572 => x"f8",
          1573 => x"70",
          1574 => x"0c",
          1575 => x"81",
          1576 => x"84",
          1577 => x"f9",
          1578 => x"7b",
          1579 => x"a0",
          1580 => x"08",
          1581 => x"90",
          1582 => x"58",
          1583 => x"53",
          1584 => x"ba",
          1585 => x"88",
          1586 => x"51",
          1587 => x"76",
          1588 => x"12",
          1589 => x"0c",
          1590 => x"0c",
          1591 => x"0c",
          1592 => x"0c",
          1593 => x"0c",
          1594 => x"0c",
          1595 => x"0c",
          1596 => x"0c",
          1597 => x"0c",
          1598 => x"0c",
          1599 => x"73",
          1600 => x"16",
          1601 => x"15",
          1602 => x"f8",
          1603 => x"3d",
          1604 => x"3d",
          1605 => x"11",
          1606 => x"08",
          1607 => x"71",
          1608 => x"09",
          1609 => x"38",
          1610 => x"70",
          1611 => x"70",
          1612 => x"81",
          1613 => x"84",
          1614 => x"84",
          1615 => x"88",
          1616 => x"8c",
          1617 => x"53",
          1618 => x"73",
          1619 => x"b0",
          1620 => x"0c",
          1621 => x"0b",
          1622 => x"72",
          1623 => x"0c",
          1624 => x"73",
          1625 => x"51",
          1626 => x"2e",
          1627 => x"b3",
          1628 => x"08",
          1629 => x"52",
          1630 => x"09",
          1631 => x"38",
          1632 => x"12",
          1633 => x"94",
          1634 => x"15",
          1635 => x"13",
          1636 => x"12",
          1637 => x"08",
          1638 => x"70",
          1639 => x"52",
          1640 => x"72",
          1641 => x"0c",
          1642 => x"04",
          1643 => x"79",
          1644 => x"76",
          1645 => x"b5",
          1646 => x"f0",
          1647 => x"b0",
          1648 => x"75",
          1649 => x"8f",
          1650 => x"08",
          1651 => x"c7",
          1652 => x"08",
          1653 => x"83",
          1654 => x"fc",
          1655 => x"70",
          1656 => x"91",
          1657 => x"c8",
          1658 => x"c8",
          1659 => x"81",
          1660 => x"07",
          1661 => x"f8",
          1662 => x"70",
          1663 => x"07",
          1664 => x"07",
          1665 => x"51",
          1666 => x"54",
          1667 => x"09",
          1668 => x"d9",
          1669 => x"76",
          1670 => x"80",
          1671 => x"0b",
          1672 => x"08",
          1673 => x"f8",
          1674 => x"05",
          1675 => x"ac",
          1676 => x"08",
          1677 => x"38",
          1678 => x"87",
          1679 => x"08",
          1680 => x"88",
          1681 => x"17",
          1682 => x"17",
          1683 => x"14",
          1684 => x"08",
          1685 => x"0c",
          1686 => x"fd",
          1687 => x"52",
          1688 => x"08",
          1689 => x"3f",
          1690 => x"08",
          1691 => x"f8",
          1692 => x"3d",
          1693 => x"3d",
          1694 => x"71",
          1695 => x"38",
          1696 => x"fd",
          1697 => x"3d",
          1698 => x"3d",
          1699 => x"05",
          1700 => x"8a",
          1701 => x"06",
          1702 => x"51",
          1703 => x"f8",
          1704 => x"71",
          1705 => x"38",
          1706 => x"81",
          1707 => x"81",
          1708 => x"e4",
          1709 => x"81",
          1710 => x"52",
          1711 => x"85",
          1712 => x"71",
          1713 => x"0d",
          1714 => x"0d",
          1715 => x"33",
          1716 => x"08",
          1717 => x"dc",
          1718 => x"ff",
          1719 => x"81",
          1720 => x"84",
          1721 => x"fd",
          1722 => x"54",
          1723 => x"81",
          1724 => x"53",
          1725 => x"8e",
          1726 => x"ff",
          1727 => x"14",
          1728 => x"3f",
          1729 => x"3d",
          1730 => x"3d",
          1731 => x"f8",
          1732 => x"81",
          1733 => x"56",
          1734 => x"70",
          1735 => x"53",
          1736 => x"2e",
          1737 => x"81",
          1738 => x"81",
          1739 => x"da",
          1740 => x"74",
          1741 => x"0c",
          1742 => x"04",
          1743 => x"66",
          1744 => x"78",
          1745 => x"5a",
          1746 => x"80",
          1747 => x"38",
          1748 => x"09",
          1749 => x"de",
          1750 => x"7a",
          1751 => x"5c",
          1752 => x"5b",
          1753 => x"09",
          1754 => x"38",
          1755 => x"39",
          1756 => x"09",
          1757 => x"38",
          1758 => x"70",
          1759 => x"33",
          1760 => x"2e",
          1761 => x"92",
          1762 => x"19",
          1763 => x"70",
          1764 => x"33",
          1765 => x"53",
          1766 => x"16",
          1767 => x"26",
          1768 => x"88",
          1769 => x"05",
          1770 => x"05",
          1771 => x"05",
          1772 => x"5b",
          1773 => x"80",
          1774 => x"30",
          1775 => x"80",
          1776 => x"cc",
          1777 => x"70",
          1778 => x"25",
          1779 => x"54",
          1780 => x"53",
          1781 => x"8c",
          1782 => x"07",
          1783 => x"05",
          1784 => x"5a",
          1785 => x"83",
          1786 => x"54",
          1787 => x"27",
          1788 => x"16",
          1789 => x"06",
          1790 => x"80",
          1791 => x"aa",
          1792 => x"cf",
          1793 => x"73",
          1794 => x"81",
          1795 => x"80",
          1796 => x"38",
          1797 => x"2e",
          1798 => x"81",
          1799 => x"80",
          1800 => x"8a",
          1801 => x"39",
          1802 => x"2e",
          1803 => x"73",
          1804 => x"8a",
          1805 => x"d3",
          1806 => x"80",
          1807 => x"80",
          1808 => x"ee",
          1809 => x"39",
          1810 => x"71",
          1811 => x"53",
          1812 => x"54",
          1813 => x"2e",
          1814 => x"15",
          1815 => x"33",
          1816 => x"72",
          1817 => x"81",
          1818 => x"39",
          1819 => x"56",
          1820 => x"27",
          1821 => x"51",
          1822 => x"75",
          1823 => x"72",
          1824 => x"38",
          1825 => x"df",
          1826 => x"16",
          1827 => x"7b",
          1828 => x"38",
          1829 => x"f2",
          1830 => x"77",
          1831 => x"12",
          1832 => x"53",
          1833 => x"5c",
          1834 => x"5c",
          1835 => x"5c",
          1836 => x"5c",
          1837 => x"51",
          1838 => x"fd",
          1839 => x"82",
          1840 => x"06",
          1841 => x"80",
          1842 => x"77",
          1843 => x"53",
          1844 => x"18",
          1845 => x"72",
          1846 => x"c4",
          1847 => x"70",
          1848 => x"25",
          1849 => x"55",
          1850 => x"8d",
          1851 => x"2e",
          1852 => x"30",
          1853 => x"5b",
          1854 => x"8f",
          1855 => x"7b",
          1856 => x"d9",
          1857 => x"f8",
          1858 => x"ff",
          1859 => x"75",
          1860 => x"9a",
          1861 => x"c8",
          1862 => x"74",
          1863 => x"a7",
          1864 => x"80",
          1865 => x"38",
          1866 => x"72",
          1867 => x"54",
          1868 => x"72",
          1869 => x"05",
          1870 => x"17",
          1871 => x"77",
          1872 => x"51",
          1873 => x"9f",
          1874 => x"72",
          1875 => x"79",
          1876 => x"81",
          1877 => x"72",
          1878 => x"38",
          1879 => x"05",
          1880 => x"ad",
          1881 => x"17",
          1882 => x"81",
          1883 => x"b0",
          1884 => x"38",
          1885 => x"81",
          1886 => x"06",
          1887 => x"9f",
          1888 => x"55",
          1889 => x"97",
          1890 => x"f9",
          1891 => x"81",
          1892 => x"8b",
          1893 => x"16",
          1894 => x"73",
          1895 => x"96",
          1896 => x"e0",
          1897 => x"17",
          1898 => x"33",
          1899 => x"f9",
          1900 => x"f2",
          1901 => x"16",
          1902 => x"7b",
          1903 => x"38",
          1904 => x"c6",
          1905 => x"96",
          1906 => x"fd",
          1907 => x"3d",
          1908 => x"05",
          1909 => x"52",
          1910 => x"e0",
          1911 => x"0d",
          1912 => x"0d",
          1913 => x"e4",
          1914 => x"88",
          1915 => x"51",
          1916 => x"81",
          1917 => x"53",
          1918 => x"80",
          1919 => x"e4",
          1920 => x"0d",
          1921 => x"0d",
          1922 => x"08",
          1923 => x"dc",
          1924 => x"88",
          1925 => x"52",
          1926 => x"3f",
          1927 => x"dc",
          1928 => x"0d",
          1929 => x"0d",
          1930 => x"f8",
          1931 => x"56",
          1932 => x"80",
          1933 => x"2e",
          1934 => x"81",
          1935 => x"52",
          1936 => x"f8",
          1937 => x"ff",
          1938 => x"80",
          1939 => x"38",
          1940 => x"b9",
          1941 => x"32",
          1942 => x"80",
          1943 => x"52",
          1944 => x"8b",
          1945 => x"2e",
          1946 => x"14",
          1947 => x"9f",
          1948 => x"38",
          1949 => x"73",
          1950 => x"38",
          1951 => x"72",
          1952 => x"14",
          1953 => x"f8",
          1954 => x"af",
          1955 => x"52",
          1956 => x"8a",
          1957 => x"3f",
          1958 => x"81",
          1959 => x"87",
          1960 => x"fe",
          1961 => x"f8",
          1962 => x"81",
          1963 => x"77",
          1964 => x"53",
          1965 => x"72",
          1966 => x"0c",
          1967 => x"04",
          1968 => x"7a",
          1969 => x"80",
          1970 => x"58",
          1971 => x"33",
          1972 => x"a0",
          1973 => x"06",
          1974 => x"13",
          1975 => x"39",
          1976 => x"09",
          1977 => x"38",
          1978 => x"11",
          1979 => x"08",
          1980 => x"54",
          1981 => x"2e",
          1982 => x"80",
          1983 => x"08",
          1984 => x"0c",
          1985 => x"33",
          1986 => x"80",
          1987 => x"38",
          1988 => x"80",
          1989 => x"38",
          1990 => x"57",
          1991 => x"0c",
          1992 => x"33",
          1993 => x"39",
          1994 => x"74",
          1995 => x"38",
          1996 => x"80",
          1997 => x"89",
          1998 => x"38",
          1999 => x"d0",
          2000 => x"55",
          2001 => x"80",
          2002 => x"39",
          2003 => x"d9",
          2004 => x"80",
          2005 => x"27",
          2006 => x"80",
          2007 => x"89",
          2008 => x"70",
          2009 => x"55",
          2010 => x"70",
          2011 => x"55",
          2012 => x"27",
          2013 => x"14",
          2014 => x"06",
          2015 => x"74",
          2016 => x"73",
          2017 => x"38",
          2018 => x"14",
          2019 => x"05",
          2020 => x"08",
          2021 => x"54",
          2022 => x"39",
          2023 => x"84",
          2024 => x"55",
          2025 => x"81",
          2026 => x"f8",
          2027 => x"3d",
          2028 => x"3d",
          2029 => x"5a",
          2030 => x"7a",
          2031 => x"08",
          2032 => x"53",
          2033 => x"09",
          2034 => x"38",
          2035 => x"0c",
          2036 => x"ad",
          2037 => x"06",
          2038 => x"76",
          2039 => x"0c",
          2040 => x"33",
          2041 => x"73",
          2042 => x"81",
          2043 => x"38",
          2044 => x"05",
          2045 => x"08",
          2046 => x"53",
          2047 => x"2e",
          2048 => x"57",
          2049 => x"2e",
          2050 => x"39",
          2051 => x"13",
          2052 => x"08",
          2053 => x"53",
          2054 => x"55",
          2055 => x"80",
          2056 => x"14",
          2057 => x"88",
          2058 => x"27",
          2059 => x"eb",
          2060 => x"53",
          2061 => x"89",
          2062 => x"38",
          2063 => x"55",
          2064 => x"8a",
          2065 => x"a0",
          2066 => x"c2",
          2067 => x"74",
          2068 => x"e0",
          2069 => x"ff",
          2070 => x"d0",
          2071 => x"ff",
          2072 => x"90",
          2073 => x"38",
          2074 => x"81",
          2075 => x"53",
          2076 => x"ca",
          2077 => x"27",
          2078 => x"77",
          2079 => x"08",
          2080 => x"0c",
          2081 => x"33",
          2082 => x"ff",
          2083 => x"80",
          2084 => x"74",
          2085 => x"79",
          2086 => x"74",
          2087 => x"0c",
          2088 => x"04",
          2089 => x"76",
          2090 => x"98",
          2091 => x"2b",
          2092 => x"72",
          2093 => x"82",
          2094 => x"51",
          2095 => x"80",
          2096 => x"c8",
          2097 => x"53",
          2098 => x"9c",
          2099 => x"c4",
          2100 => x"02",
          2101 => x"05",
          2102 => x"52",
          2103 => x"72",
          2104 => x"06",
          2105 => x"53",
          2106 => x"c8",
          2107 => x"0d",
          2108 => x"0d",
          2109 => x"05",
          2110 => x"71",
          2111 => x"53",
          2112 => x"9f",
          2113 => x"f3",
          2114 => x"51",
          2115 => x"88",
          2116 => x"3f",
          2117 => x"05",
          2118 => x"34",
          2119 => x"06",
          2120 => x"76",
          2121 => x"3f",
          2122 => x"86",
          2123 => x"f6",
          2124 => x"02",
          2125 => x"05",
          2126 => x"05",
          2127 => x"81",
          2128 => x"70",
          2129 => x"f4",
          2130 => x"08",
          2131 => x"5a",
          2132 => x"80",
          2133 => x"74",
          2134 => x"3f",
          2135 => x"33",
          2136 => x"81",
          2137 => x"81",
          2138 => x"58",
          2139 => x"bc",
          2140 => x"c8",
          2141 => x"81",
          2142 => x"70",
          2143 => x"f4",
          2144 => x"08",
          2145 => x"74",
          2146 => x"38",
          2147 => x"52",
          2148 => x"a1",
          2149 => x"94",
          2150 => x"55",
          2151 => x"94",
          2152 => x"ff",
          2153 => x"75",
          2154 => x"80",
          2155 => x"94",
          2156 => x"2e",
          2157 => x"f5",
          2158 => x"75",
          2159 => x"38",
          2160 => x"33",
          2161 => x"38",
          2162 => x"05",
          2163 => x"78",
          2164 => x"80",
          2165 => x"81",
          2166 => x"52",
          2167 => x"fd",
          2168 => x"f5",
          2169 => x"80",
          2170 => x"8c",
          2171 => x"dc",
          2172 => x"57",
          2173 => x"f5",
          2174 => x"80",
          2175 => x"81",
          2176 => x"80",
          2177 => x"f5",
          2178 => x"80",
          2179 => x"3d",
          2180 => x"80",
          2181 => x"81",
          2182 => x"80",
          2183 => x"75",
          2184 => x"3f",
          2185 => x"08",
          2186 => x"81",
          2187 => x"25",
          2188 => x"f8",
          2189 => x"05",
          2190 => x"55",
          2191 => x"75",
          2192 => x"81",
          2193 => x"dc",
          2194 => x"ff",
          2195 => x"2e",
          2196 => x"ff",
          2197 => x"3d",
          2198 => x"3d",
          2199 => x"08",
          2200 => x"5a",
          2201 => x"58",
          2202 => x"81",
          2203 => x"51",
          2204 => x"3f",
          2205 => x"08",
          2206 => x"ff",
          2207 => x"90",
          2208 => x"80",
          2209 => x"3d",
          2210 => x"80",
          2211 => x"81",
          2212 => x"80",
          2213 => x"75",
          2214 => x"3f",
          2215 => x"08",
          2216 => x"55",
          2217 => x"f8",
          2218 => x"8e",
          2219 => x"c8",
          2220 => x"70",
          2221 => x"80",
          2222 => x"09",
          2223 => x"72",
          2224 => x"51",
          2225 => x"77",
          2226 => x"73",
          2227 => x"81",
          2228 => x"8c",
          2229 => x"51",
          2230 => x"3f",
          2231 => x"08",
          2232 => x"38",
          2233 => x"51",
          2234 => x"78",
          2235 => x"81",
          2236 => x"75",
          2237 => x"d5",
          2238 => x"51",
          2239 => x"ab",
          2240 => x"81",
          2241 => x"74",
          2242 => x"77",
          2243 => x"0c",
          2244 => x"04",
          2245 => x"7c",
          2246 => x"71",
          2247 => x"59",
          2248 => x"a0",
          2249 => x"06",
          2250 => x"33",
          2251 => x"77",
          2252 => x"38",
          2253 => x"5b",
          2254 => x"56",
          2255 => x"a0",
          2256 => x"06",
          2257 => x"75",
          2258 => x"80",
          2259 => x"29",
          2260 => x"05",
          2261 => x"55",
          2262 => x"81",
          2263 => x"53",
          2264 => x"08",
          2265 => x"3f",
          2266 => x"08",
          2267 => x"84",
          2268 => x"74",
          2269 => x"38",
          2270 => x"88",
          2271 => x"fc",
          2272 => x"39",
          2273 => x"8c",
          2274 => x"53",
          2275 => x"f6",
          2276 => x"f8",
          2277 => x"2e",
          2278 => x"53",
          2279 => x"51",
          2280 => x"81",
          2281 => x"81",
          2282 => x"74",
          2283 => x"54",
          2284 => x"14",
          2285 => x"06",
          2286 => x"74",
          2287 => x"38",
          2288 => x"81",
          2289 => x"8c",
          2290 => x"d3",
          2291 => x"3d",
          2292 => x"05",
          2293 => x"33",
          2294 => x"0b",
          2295 => x"81",
          2296 => x"5b",
          2297 => x"08",
          2298 => x"81",
          2299 => x"54",
          2300 => x"38",
          2301 => x"b4",
          2302 => x"c8",
          2303 => x"90",
          2304 => x"c8",
          2305 => x"80",
          2306 => x"53",
          2307 => x"08",
          2308 => x"c8",
          2309 => x"ed",
          2310 => x"c8",
          2311 => x"8b",
          2312 => x"94",
          2313 => x"3f",
          2314 => x"81",
          2315 => x"53",
          2316 => x"90",
          2317 => x"54",
          2318 => x"3f",
          2319 => x"08",
          2320 => x"c8",
          2321 => x"09",
          2322 => x"c1",
          2323 => x"c8",
          2324 => x"fc",
          2325 => x"c8",
          2326 => x"0b",
          2327 => x"08",
          2328 => x"81",
          2329 => x"ff",
          2330 => x"55",
          2331 => x"34",
          2332 => x"81",
          2333 => x"75",
          2334 => x"3f",
          2335 => x"09",
          2336 => x"a7",
          2337 => x"81",
          2338 => x"8c",
          2339 => x"5d",
          2340 => x"81",
          2341 => x"98",
          2342 => x"2c",
          2343 => x"ff",
          2344 => x"78",
          2345 => x"81",
          2346 => x"70",
          2347 => x"98",
          2348 => x"e8",
          2349 => x"2b",
          2350 => x"71",
          2351 => x"70",
          2352 => x"e4",
          2353 => x"08",
          2354 => x"51",
          2355 => x"59",
          2356 => x"5d",
          2357 => x"73",
          2358 => x"e9",
          2359 => x"27",
          2360 => x"81",
          2361 => x"81",
          2362 => x"70",
          2363 => x"55",
          2364 => x"80",
          2365 => x"53",
          2366 => x"51",
          2367 => x"81",
          2368 => x"81",
          2369 => x"73",
          2370 => x"38",
          2371 => x"e8",
          2372 => x"b1",
          2373 => x"80",
          2374 => x"80",
          2375 => x"98",
          2376 => x"ff",
          2377 => x"55",
          2378 => x"97",
          2379 => x"74",
          2380 => x"f6",
          2381 => x"f8",
          2382 => x"ff",
          2383 => x"cc",
          2384 => x"80",
          2385 => x"2e",
          2386 => x"81",
          2387 => x"81",
          2388 => x"74",
          2389 => x"98",
          2390 => x"e8",
          2391 => x"2b",
          2392 => x"70",
          2393 => x"82",
          2394 => x"c8",
          2395 => x"51",
          2396 => x"58",
          2397 => x"77",
          2398 => x"06",
          2399 => x"81",
          2400 => x"08",
          2401 => x"0b",
          2402 => x"34",
          2403 => x"f8",
          2404 => x"39",
          2405 => x"ec",
          2406 => x"f8",
          2407 => x"af",
          2408 => x"7d",
          2409 => x"73",
          2410 => x"e1",
          2411 => x"29",
          2412 => x"05",
          2413 => x"04",
          2414 => x"33",
          2415 => x"2e",
          2416 => x"81",
          2417 => x"55",
          2418 => x"ab",
          2419 => x"2b",
          2420 => x"51",
          2421 => x"24",
          2422 => x"1a",
          2423 => x"81",
          2424 => x"81",
          2425 => x"81",
          2426 => x"70",
          2427 => x"f8",
          2428 => x"51",
          2429 => x"81",
          2430 => x"81",
          2431 => x"74",
          2432 => x"34",
          2433 => x"ae",
          2434 => x"34",
          2435 => x"33",
          2436 => x"27",
          2437 => x"14",
          2438 => x"f8",
          2439 => x"f8",
          2440 => x"81",
          2441 => x"81",
          2442 => x"70",
          2443 => x"f8",
          2444 => x"51",
          2445 => x"77",
          2446 => x"74",
          2447 => x"52",
          2448 => x"3f",
          2449 => x"0a",
          2450 => x"0a",
          2451 => x"2c",
          2452 => x"33",
          2453 => x"73",
          2454 => x"38",
          2455 => x"33",
          2456 => x"70",
          2457 => x"f8",
          2458 => x"51",
          2459 => x"77",
          2460 => x"38",
          2461 => x"92",
          2462 => x"80",
          2463 => x"80",
          2464 => x"98",
          2465 => x"f0",
          2466 => x"55",
          2467 => x"e4",
          2468 => x"39",
          2469 => x"33",
          2470 => x"06",
          2471 => x"80",
          2472 => x"38",
          2473 => x"33",
          2474 => x"73",
          2475 => x"34",
          2476 => x"73",
          2477 => x"34",
          2478 => x"ce",
          2479 => x"f4",
          2480 => x"2b",
          2481 => x"81",
          2482 => x"57",
          2483 => x"74",
          2484 => x"38",
          2485 => x"81",
          2486 => x"34",
          2487 => x"e7",
          2488 => x"81",
          2489 => x"81",
          2490 => x"70",
          2491 => x"f8",
          2492 => x"51",
          2493 => x"24",
          2494 => x"51",
          2495 => x"81",
          2496 => x"70",
          2497 => x"98",
          2498 => x"f0",
          2499 => x"56",
          2500 => x"24",
          2501 => x"88",
          2502 => x"3f",
          2503 => x"0a",
          2504 => x"0a",
          2505 => x"2c",
          2506 => x"33",
          2507 => x"75",
          2508 => x"38",
          2509 => x"81",
          2510 => x"7a",
          2511 => x"74",
          2512 => x"e6",
          2513 => x"f8",
          2514 => x"51",
          2515 => x"81",
          2516 => x"81",
          2517 => x"73",
          2518 => x"f8",
          2519 => x"73",
          2520 => x"c9",
          2521 => x"73",
          2522 => x"f3",
          2523 => x"bd",
          2524 => x"34",
          2525 => x"81",
          2526 => x"54",
          2527 => x"fa",
          2528 => x"51",
          2529 => x"81",
          2530 => x"ff",
          2531 => x"81",
          2532 => x"73",
          2533 => x"54",
          2534 => x"f8",
          2535 => x"f8",
          2536 => x"55",
          2537 => x"f9",
          2538 => x"14",
          2539 => x"f8",
          2540 => x"98",
          2541 => x"2c",
          2542 => x"06",
          2543 => x"74",
          2544 => x"38",
          2545 => x"81",
          2546 => x"34",
          2547 => x"e5",
          2548 => x"81",
          2549 => x"81",
          2550 => x"70",
          2551 => x"f8",
          2552 => x"51",
          2553 => x"24",
          2554 => x"51",
          2555 => x"81",
          2556 => x"70",
          2557 => x"98",
          2558 => x"f0",
          2559 => x"56",
          2560 => x"24",
          2561 => x"88",
          2562 => x"3f",
          2563 => x"0a",
          2564 => x"0a",
          2565 => x"2c",
          2566 => x"33",
          2567 => x"75",
          2568 => x"38",
          2569 => x"81",
          2570 => x"70",
          2571 => x"81",
          2572 => x"59",
          2573 => x"77",
          2574 => x"38",
          2575 => x"73",
          2576 => x"34",
          2577 => x"33",
          2578 => x"be",
          2579 => x"f4",
          2580 => x"ff",
          2581 => x"f0",
          2582 => x"54",
          2583 => x"dc",
          2584 => x"39",
          2585 => x"81",
          2586 => x"55",
          2587 => x"a4",
          2588 => x"cb",
          2589 => x"f8",
          2590 => x"f8",
          2591 => x"f8",
          2592 => x"ff",
          2593 => x"53",
          2594 => x"51",
          2595 => x"93",
          2596 => x"39",
          2597 => x"81",
          2598 => x"fc",
          2599 => x"54",
          2600 => x"a5",
          2601 => x"cb",
          2602 => x"f8",
          2603 => x"f8",
          2604 => x"f8",
          2605 => x"ff",
          2606 => x"53",
          2607 => x"51",
          2608 => x"ff",
          2609 => x"de",
          2610 => x"55",
          2611 => x"f7",
          2612 => x"51",
          2613 => x"80",
          2614 => x"93",
          2615 => x"06",
          2616 => x"f4",
          2617 => x"74",
          2618 => x"38",
          2619 => x"e0",
          2620 => x"39",
          2621 => x"81",
          2622 => x"84",
          2623 => x"54",
          2624 => x"a9",
          2625 => x"ca",
          2626 => x"f8",
          2627 => x"f8",
          2628 => x"f8",
          2629 => x"ff",
          2630 => x"53",
          2631 => x"51",
          2632 => x"81",
          2633 => x"81",
          2634 => x"a8",
          2635 => x"55",
          2636 => x"f6",
          2637 => x"51",
          2638 => x"81",
          2639 => x"81",
          2640 => x"81",
          2641 => x"81",
          2642 => x"05",
          2643 => x"79",
          2644 => x"3f",
          2645 => x"53",
          2646 => x"33",
          2647 => x"ef",
          2648 => x"a9",
          2649 => x"f4",
          2650 => x"ff",
          2651 => x"f0",
          2652 => x"54",
          2653 => x"f6",
          2654 => x"14",
          2655 => x"f8",
          2656 => x"1a",
          2657 => x"54",
          2658 => x"f6",
          2659 => x"f8",
          2660 => x"73",
          2661 => x"f5",
          2662 => x"e1",
          2663 => x"f8",
          2664 => x"05",
          2665 => x"f8",
          2666 => x"e1",
          2667 => x"81",
          2668 => x"80",
          2669 => x"f0",
          2670 => x"f8",
          2671 => x"3d",
          2672 => x"3d",
          2673 => x"05",
          2674 => x"52",
          2675 => x"87",
          2676 => x"b0",
          2677 => x"71",
          2678 => x"0c",
          2679 => x"04",
          2680 => x"02",
          2681 => x"02",
          2682 => x"05",
          2683 => x"83",
          2684 => x"26",
          2685 => x"72",
          2686 => x"c0",
          2687 => x"53",
          2688 => x"74",
          2689 => x"38",
          2690 => x"73",
          2691 => x"c0",
          2692 => x"51",
          2693 => x"85",
          2694 => x"98",
          2695 => x"52",
          2696 => x"82",
          2697 => x"70",
          2698 => x"38",
          2699 => x"8c",
          2700 => x"ec",
          2701 => x"fc",
          2702 => x"52",
          2703 => x"87",
          2704 => x"08",
          2705 => x"2e",
          2706 => x"81",
          2707 => x"34",
          2708 => x"13",
          2709 => x"81",
          2710 => x"86",
          2711 => x"f3",
          2712 => x"62",
          2713 => x"05",
          2714 => x"57",
          2715 => x"83",
          2716 => x"fe",
          2717 => x"f8",
          2718 => x"06",
          2719 => x"71",
          2720 => x"71",
          2721 => x"2b",
          2722 => x"80",
          2723 => x"92",
          2724 => x"c0",
          2725 => x"41",
          2726 => x"5a",
          2727 => x"87",
          2728 => x"0c",
          2729 => x"84",
          2730 => x"08",
          2731 => x"70",
          2732 => x"53",
          2733 => x"2e",
          2734 => x"08",
          2735 => x"70",
          2736 => x"34",
          2737 => x"80",
          2738 => x"53",
          2739 => x"2e",
          2740 => x"53",
          2741 => x"26",
          2742 => x"80",
          2743 => x"87",
          2744 => x"08",
          2745 => x"38",
          2746 => x"8c",
          2747 => x"80",
          2748 => x"78",
          2749 => x"99",
          2750 => x"0c",
          2751 => x"8c",
          2752 => x"08",
          2753 => x"51",
          2754 => x"38",
          2755 => x"8d",
          2756 => x"17",
          2757 => x"81",
          2758 => x"53",
          2759 => x"2e",
          2760 => x"fc",
          2761 => x"52",
          2762 => x"7d",
          2763 => x"ed",
          2764 => x"80",
          2765 => x"71",
          2766 => x"38",
          2767 => x"53",
          2768 => x"c8",
          2769 => x"0d",
          2770 => x"0d",
          2771 => x"02",
          2772 => x"05",
          2773 => x"58",
          2774 => x"80",
          2775 => x"fc",
          2776 => x"f8",
          2777 => x"06",
          2778 => x"71",
          2779 => x"81",
          2780 => x"38",
          2781 => x"2b",
          2782 => x"80",
          2783 => x"92",
          2784 => x"c0",
          2785 => x"40",
          2786 => x"5a",
          2787 => x"c0",
          2788 => x"76",
          2789 => x"76",
          2790 => x"75",
          2791 => x"2a",
          2792 => x"51",
          2793 => x"80",
          2794 => x"7a",
          2795 => x"5c",
          2796 => x"81",
          2797 => x"81",
          2798 => x"06",
          2799 => x"80",
          2800 => x"87",
          2801 => x"08",
          2802 => x"38",
          2803 => x"8c",
          2804 => x"80",
          2805 => x"77",
          2806 => x"99",
          2807 => x"0c",
          2808 => x"8c",
          2809 => x"08",
          2810 => x"51",
          2811 => x"38",
          2812 => x"8d",
          2813 => x"70",
          2814 => x"84",
          2815 => x"5b",
          2816 => x"2e",
          2817 => x"fc",
          2818 => x"52",
          2819 => x"7d",
          2820 => x"f8",
          2821 => x"80",
          2822 => x"71",
          2823 => x"38",
          2824 => x"53",
          2825 => x"c8",
          2826 => x"0d",
          2827 => x"0d",
          2828 => x"05",
          2829 => x"02",
          2830 => x"05",
          2831 => x"54",
          2832 => x"fe",
          2833 => x"c8",
          2834 => x"53",
          2835 => x"80",
          2836 => x"0b",
          2837 => x"8c",
          2838 => x"71",
          2839 => x"dc",
          2840 => x"24",
          2841 => x"84",
          2842 => x"92",
          2843 => x"54",
          2844 => x"8d",
          2845 => x"39",
          2846 => x"80",
          2847 => x"cb",
          2848 => x"70",
          2849 => x"81",
          2850 => x"52",
          2851 => x"8a",
          2852 => x"98",
          2853 => x"71",
          2854 => x"c0",
          2855 => x"52",
          2856 => x"81",
          2857 => x"c0",
          2858 => x"53",
          2859 => x"82",
          2860 => x"71",
          2861 => x"39",
          2862 => x"39",
          2863 => x"77",
          2864 => x"81",
          2865 => x"72",
          2866 => x"84",
          2867 => x"73",
          2868 => x"0c",
          2869 => x"04",
          2870 => x"74",
          2871 => x"71",
          2872 => x"2b",
          2873 => x"c8",
          2874 => x"84",
          2875 => x"fd",
          2876 => x"83",
          2877 => x"12",
          2878 => x"2b",
          2879 => x"07",
          2880 => x"70",
          2881 => x"2b",
          2882 => x"07",
          2883 => x"0c",
          2884 => x"56",
          2885 => x"3d",
          2886 => x"3d",
          2887 => x"84",
          2888 => x"22",
          2889 => x"72",
          2890 => x"54",
          2891 => x"2a",
          2892 => x"34",
          2893 => x"04",
          2894 => x"73",
          2895 => x"70",
          2896 => x"05",
          2897 => x"88",
          2898 => x"72",
          2899 => x"54",
          2900 => x"2a",
          2901 => x"70",
          2902 => x"34",
          2903 => x"51",
          2904 => x"83",
          2905 => x"fe",
          2906 => x"75",
          2907 => x"51",
          2908 => x"92",
          2909 => x"81",
          2910 => x"73",
          2911 => x"55",
          2912 => x"51",
          2913 => x"3d",
          2914 => x"3d",
          2915 => x"76",
          2916 => x"72",
          2917 => x"05",
          2918 => x"11",
          2919 => x"38",
          2920 => x"04",
          2921 => x"78",
          2922 => x"56",
          2923 => x"81",
          2924 => x"74",
          2925 => x"56",
          2926 => x"31",
          2927 => x"52",
          2928 => x"80",
          2929 => x"71",
          2930 => x"38",
          2931 => x"c8",
          2932 => x"0d",
          2933 => x"0d",
          2934 => x"51",
          2935 => x"73",
          2936 => x"81",
          2937 => x"33",
          2938 => x"38",
          2939 => x"f8",
          2940 => x"3d",
          2941 => x"0b",
          2942 => x"0c",
          2943 => x"81",
          2944 => x"04",
          2945 => x"7b",
          2946 => x"83",
          2947 => x"5a",
          2948 => x"80",
          2949 => x"54",
          2950 => x"53",
          2951 => x"53",
          2952 => x"52",
          2953 => x"3f",
          2954 => x"08",
          2955 => x"81",
          2956 => x"81",
          2957 => x"83",
          2958 => x"16",
          2959 => x"18",
          2960 => x"18",
          2961 => x"58",
          2962 => x"9f",
          2963 => x"33",
          2964 => x"2e",
          2965 => x"93",
          2966 => x"76",
          2967 => x"52",
          2968 => x"51",
          2969 => x"83",
          2970 => x"79",
          2971 => x"0c",
          2972 => x"04",
          2973 => x"78",
          2974 => x"80",
          2975 => x"17",
          2976 => x"38",
          2977 => x"fc",
          2978 => x"c8",
          2979 => x"f8",
          2980 => x"38",
          2981 => x"53",
          2982 => x"81",
          2983 => x"f7",
          2984 => x"f8",
          2985 => x"2e",
          2986 => x"55",
          2987 => x"b0",
          2988 => x"81",
          2989 => x"88",
          2990 => x"f8",
          2991 => x"70",
          2992 => x"c0",
          2993 => x"c8",
          2994 => x"f8",
          2995 => x"91",
          2996 => x"55",
          2997 => x"09",
          2998 => x"f0",
          2999 => x"33",
          3000 => x"2e",
          3001 => x"80",
          3002 => x"80",
          3003 => x"c8",
          3004 => x"17",
          3005 => x"fd",
          3006 => x"d4",
          3007 => x"b2",
          3008 => x"96",
          3009 => x"85",
          3010 => x"75",
          3011 => x"3f",
          3012 => x"e4",
          3013 => x"98",
          3014 => x"9c",
          3015 => x"08",
          3016 => x"17",
          3017 => x"3f",
          3018 => x"52",
          3019 => x"51",
          3020 => x"a0",
          3021 => x"05",
          3022 => x"0c",
          3023 => x"75",
          3024 => x"33",
          3025 => x"3f",
          3026 => x"34",
          3027 => x"52",
          3028 => x"51",
          3029 => x"81",
          3030 => x"80",
          3031 => x"81",
          3032 => x"f8",
          3033 => x"3d",
          3034 => x"3d",
          3035 => x"1a",
          3036 => x"fe",
          3037 => x"54",
          3038 => x"73",
          3039 => x"8a",
          3040 => x"71",
          3041 => x"08",
          3042 => x"75",
          3043 => x"0c",
          3044 => x"04",
          3045 => x"7a",
          3046 => x"56",
          3047 => x"77",
          3048 => x"38",
          3049 => x"08",
          3050 => x"38",
          3051 => x"54",
          3052 => x"2e",
          3053 => x"72",
          3054 => x"38",
          3055 => x"8d",
          3056 => x"39",
          3057 => x"81",
          3058 => x"b6",
          3059 => x"2a",
          3060 => x"2a",
          3061 => x"05",
          3062 => x"55",
          3063 => x"81",
          3064 => x"81",
          3065 => x"83",
          3066 => x"b4",
          3067 => x"17",
          3068 => x"a4",
          3069 => x"55",
          3070 => x"57",
          3071 => x"3f",
          3072 => x"08",
          3073 => x"74",
          3074 => x"14",
          3075 => x"70",
          3076 => x"07",
          3077 => x"71",
          3078 => x"52",
          3079 => x"72",
          3080 => x"75",
          3081 => x"58",
          3082 => x"76",
          3083 => x"15",
          3084 => x"73",
          3085 => x"3f",
          3086 => x"08",
          3087 => x"76",
          3088 => x"06",
          3089 => x"05",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"06",
          3093 => x"76",
          3094 => x"15",
          3095 => x"73",
          3096 => x"3f",
          3097 => x"08",
          3098 => x"82",
          3099 => x"06",
          3100 => x"05",
          3101 => x"3f",
          3102 => x"08",
          3103 => x"58",
          3104 => x"58",
          3105 => x"c8",
          3106 => x"0d",
          3107 => x"0d",
          3108 => x"5a",
          3109 => x"59",
          3110 => x"82",
          3111 => x"98",
          3112 => x"82",
          3113 => x"33",
          3114 => x"2e",
          3115 => x"72",
          3116 => x"38",
          3117 => x"8d",
          3118 => x"39",
          3119 => x"81",
          3120 => x"f7",
          3121 => x"2a",
          3122 => x"2a",
          3123 => x"05",
          3124 => x"55",
          3125 => x"81",
          3126 => x"59",
          3127 => x"08",
          3128 => x"74",
          3129 => x"16",
          3130 => x"16",
          3131 => x"59",
          3132 => x"53",
          3133 => x"8f",
          3134 => x"2b",
          3135 => x"74",
          3136 => x"71",
          3137 => x"72",
          3138 => x"0b",
          3139 => x"74",
          3140 => x"17",
          3141 => x"75",
          3142 => x"3f",
          3143 => x"08",
          3144 => x"c8",
          3145 => x"38",
          3146 => x"06",
          3147 => x"78",
          3148 => x"54",
          3149 => x"77",
          3150 => x"33",
          3151 => x"71",
          3152 => x"51",
          3153 => x"34",
          3154 => x"76",
          3155 => x"17",
          3156 => x"75",
          3157 => x"3f",
          3158 => x"08",
          3159 => x"c8",
          3160 => x"38",
          3161 => x"ff",
          3162 => x"10",
          3163 => x"76",
          3164 => x"51",
          3165 => x"be",
          3166 => x"2a",
          3167 => x"05",
          3168 => x"f9",
          3169 => x"f8",
          3170 => x"81",
          3171 => x"ab",
          3172 => x"0a",
          3173 => x"2b",
          3174 => x"70",
          3175 => x"70",
          3176 => x"54",
          3177 => x"81",
          3178 => x"8f",
          3179 => x"07",
          3180 => x"f7",
          3181 => x"0b",
          3182 => x"78",
          3183 => x"0c",
          3184 => x"04",
          3185 => x"7a",
          3186 => x"08",
          3187 => x"59",
          3188 => x"a4",
          3189 => x"17",
          3190 => x"38",
          3191 => x"aa",
          3192 => x"73",
          3193 => x"fd",
          3194 => x"f8",
          3195 => x"81",
          3196 => x"80",
          3197 => x"39",
          3198 => x"eb",
          3199 => x"80",
          3200 => x"f8",
          3201 => x"80",
          3202 => x"52",
          3203 => x"84",
          3204 => x"c8",
          3205 => x"f8",
          3206 => x"2e",
          3207 => x"81",
          3208 => x"81",
          3209 => x"81",
          3210 => x"ff",
          3211 => x"80",
          3212 => x"75",
          3213 => x"3f",
          3214 => x"08",
          3215 => x"16",
          3216 => x"90",
          3217 => x"55",
          3218 => x"27",
          3219 => x"15",
          3220 => x"84",
          3221 => x"07",
          3222 => x"17",
          3223 => x"76",
          3224 => x"a6",
          3225 => x"73",
          3226 => x"0c",
          3227 => x"04",
          3228 => x"7c",
          3229 => x"59",
          3230 => x"95",
          3231 => x"08",
          3232 => x"2e",
          3233 => x"17",
          3234 => x"b2",
          3235 => x"ae",
          3236 => x"7a",
          3237 => x"3f",
          3238 => x"81",
          3239 => x"27",
          3240 => x"81",
          3241 => x"55",
          3242 => x"08",
          3243 => x"d2",
          3244 => x"08",
          3245 => x"08",
          3246 => x"38",
          3247 => x"17",
          3248 => x"54",
          3249 => x"82",
          3250 => x"7a",
          3251 => x"06",
          3252 => x"81",
          3253 => x"17",
          3254 => x"83",
          3255 => x"75",
          3256 => x"f9",
          3257 => x"59",
          3258 => x"08",
          3259 => x"81",
          3260 => x"81",
          3261 => x"59",
          3262 => x"08",
          3263 => x"70",
          3264 => x"25",
          3265 => x"81",
          3266 => x"54",
          3267 => x"55",
          3268 => x"38",
          3269 => x"08",
          3270 => x"38",
          3271 => x"54",
          3272 => x"90",
          3273 => x"18",
          3274 => x"38",
          3275 => x"39",
          3276 => x"38",
          3277 => x"16",
          3278 => x"08",
          3279 => x"38",
          3280 => x"78",
          3281 => x"38",
          3282 => x"51",
          3283 => x"81",
          3284 => x"80",
          3285 => x"80",
          3286 => x"c8",
          3287 => x"09",
          3288 => x"38",
          3289 => x"08",
          3290 => x"c8",
          3291 => x"30",
          3292 => x"80",
          3293 => x"07",
          3294 => x"55",
          3295 => x"38",
          3296 => x"09",
          3297 => x"ae",
          3298 => x"80",
          3299 => x"53",
          3300 => x"51",
          3301 => x"81",
          3302 => x"81",
          3303 => x"30",
          3304 => x"c8",
          3305 => x"25",
          3306 => x"79",
          3307 => x"38",
          3308 => x"8f",
          3309 => x"79",
          3310 => x"f9",
          3311 => x"f8",
          3312 => x"74",
          3313 => x"8c",
          3314 => x"17",
          3315 => x"90",
          3316 => x"54",
          3317 => x"86",
          3318 => x"90",
          3319 => x"17",
          3320 => x"54",
          3321 => x"34",
          3322 => x"56",
          3323 => x"90",
          3324 => x"80",
          3325 => x"81",
          3326 => x"55",
          3327 => x"56",
          3328 => x"81",
          3329 => x"8c",
          3330 => x"f8",
          3331 => x"70",
          3332 => x"f0",
          3333 => x"c8",
          3334 => x"56",
          3335 => x"08",
          3336 => x"7b",
          3337 => x"f6",
          3338 => x"f8",
          3339 => x"f8",
          3340 => x"17",
          3341 => x"80",
          3342 => x"b4",
          3343 => x"57",
          3344 => x"77",
          3345 => x"81",
          3346 => x"15",
          3347 => x"78",
          3348 => x"81",
          3349 => x"53",
          3350 => x"15",
          3351 => x"e9",
          3352 => x"c8",
          3353 => x"df",
          3354 => x"22",
          3355 => x"30",
          3356 => x"70",
          3357 => x"51",
          3358 => x"81",
          3359 => x"8a",
          3360 => x"f8",
          3361 => x"7c",
          3362 => x"56",
          3363 => x"80",
          3364 => x"f1",
          3365 => x"06",
          3366 => x"e9",
          3367 => x"18",
          3368 => x"08",
          3369 => x"38",
          3370 => x"82",
          3371 => x"38",
          3372 => x"54",
          3373 => x"74",
          3374 => x"82",
          3375 => x"22",
          3376 => x"79",
          3377 => x"38",
          3378 => x"98",
          3379 => x"cd",
          3380 => x"22",
          3381 => x"54",
          3382 => x"26",
          3383 => x"52",
          3384 => x"b0",
          3385 => x"c8",
          3386 => x"f8",
          3387 => x"2e",
          3388 => x"0b",
          3389 => x"08",
          3390 => x"98",
          3391 => x"f8",
          3392 => x"85",
          3393 => x"bd",
          3394 => x"31",
          3395 => x"73",
          3396 => x"f4",
          3397 => x"f8",
          3398 => x"18",
          3399 => x"18",
          3400 => x"08",
          3401 => x"72",
          3402 => x"38",
          3403 => x"58",
          3404 => x"89",
          3405 => x"18",
          3406 => x"ff",
          3407 => x"05",
          3408 => x"80",
          3409 => x"f8",
          3410 => x"3d",
          3411 => x"3d",
          3412 => x"08",
          3413 => x"a0",
          3414 => x"54",
          3415 => x"77",
          3416 => x"80",
          3417 => x"0c",
          3418 => x"53",
          3419 => x"80",
          3420 => x"38",
          3421 => x"06",
          3422 => x"b5",
          3423 => x"98",
          3424 => x"14",
          3425 => x"92",
          3426 => x"2a",
          3427 => x"56",
          3428 => x"26",
          3429 => x"80",
          3430 => x"16",
          3431 => x"77",
          3432 => x"53",
          3433 => x"38",
          3434 => x"51",
          3435 => x"81",
          3436 => x"53",
          3437 => x"0b",
          3438 => x"08",
          3439 => x"38",
          3440 => x"f8",
          3441 => x"2e",
          3442 => x"98",
          3443 => x"f8",
          3444 => x"80",
          3445 => x"8a",
          3446 => x"15",
          3447 => x"80",
          3448 => x"14",
          3449 => x"51",
          3450 => x"81",
          3451 => x"53",
          3452 => x"f8",
          3453 => x"2e",
          3454 => x"82",
          3455 => x"c8",
          3456 => x"ba",
          3457 => x"81",
          3458 => x"ff",
          3459 => x"81",
          3460 => x"52",
          3461 => x"f3",
          3462 => x"c8",
          3463 => x"72",
          3464 => x"72",
          3465 => x"f2",
          3466 => x"f8",
          3467 => x"15",
          3468 => x"15",
          3469 => x"b4",
          3470 => x"0c",
          3471 => x"81",
          3472 => x"8a",
          3473 => x"f7",
          3474 => x"7d",
          3475 => x"5b",
          3476 => x"76",
          3477 => x"3f",
          3478 => x"08",
          3479 => x"c8",
          3480 => x"38",
          3481 => x"08",
          3482 => x"08",
          3483 => x"f0",
          3484 => x"f8",
          3485 => x"81",
          3486 => x"80",
          3487 => x"f8",
          3488 => x"18",
          3489 => x"51",
          3490 => x"81",
          3491 => x"81",
          3492 => x"81",
          3493 => x"c8",
          3494 => x"83",
          3495 => x"77",
          3496 => x"72",
          3497 => x"38",
          3498 => x"75",
          3499 => x"81",
          3500 => x"a5",
          3501 => x"c8",
          3502 => x"52",
          3503 => x"8e",
          3504 => x"c8",
          3505 => x"f8",
          3506 => x"2e",
          3507 => x"73",
          3508 => x"81",
          3509 => x"87",
          3510 => x"f8",
          3511 => x"3d",
          3512 => x"3d",
          3513 => x"11",
          3514 => x"ec",
          3515 => x"c8",
          3516 => x"ff",
          3517 => x"33",
          3518 => x"71",
          3519 => x"81",
          3520 => x"94",
          3521 => x"d0",
          3522 => x"c8",
          3523 => x"73",
          3524 => x"81",
          3525 => x"85",
          3526 => x"fc",
          3527 => x"79",
          3528 => x"ff",
          3529 => x"12",
          3530 => x"eb",
          3531 => x"70",
          3532 => x"72",
          3533 => x"81",
          3534 => x"73",
          3535 => x"94",
          3536 => x"d6",
          3537 => x"0d",
          3538 => x"0d",
          3539 => x"55",
          3540 => x"5a",
          3541 => x"08",
          3542 => x"8a",
          3543 => x"08",
          3544 => x"ee",
          3545 => x"f8",
          3546 => x"81",
          3547 => x"80",
          3548 => x"15",
          3549 => x"55",
          3550 => x"38",
          3551 => x"e6",
          3552 => x"33",
          3553 => x"70",
          3554 => x"58",
          3555 => x"86",
          3556 => x"f8",
          3557 => x"73",
          3558 => x"83",
          3559 => x"73",
          3560 => x"38",
          3561 => x"06",
          3562 => x"80",
          3563 => x"75",
          3564 => x"38",
          3565 => x"08",
          3566 => x"54",
          3567 => x"2e",
          3568 => x"83",
          3569 => x"73",
          3570 => x"38",
          3571 => x"51",
          3572 => x"81",
          3573 => x"58",
          3574 => x"08",
          3575 => x"15",
          3576 => x"38",
          3577 => x"0b",
          3578 => x"77",
          3579 => x"0c",
          3580 => x"04",
          3581 => x"77",
          3582 => x"54",
          3583 => x"51",
          3584 => x"81",
          3585 => x"55",
          3586 => x"08",
          3587 => x"14",
          3588 => x"51",
          3589 => x"81",
          3590 => x"55",
          3591 => x"08",
          3592 => x"53",
          3593 => x"08",
          3594 => x"08",
          3595 => x"3f",
          3596 => x"14",
          3597 => x"08",
          3598 => x"3f",
          3599 => x"17",
          3600 => x"f8",
          3601 => x"3d",
          3602 => x"3d",
          3603 => x"08",
          3604 => x"54",
          3605 => x"53",
          3606 => x"81",
          3607 => x"8d",
          3608 => x"08",
          3609 => x"34",
          3610 => x"15",
          3611 => x"0d",
          3612 => x"0d",
          3613 => x"57",
          3614 => x"17",
          3615 => x"08",
          3616 => x"82",
          3617 => x"89",
          3618 => x"55",
          3619 => x"14",
          3620 => x"16",
          3621 => x"71",
          3622 => x"38",
          3623 => x"09",
          3624 => x"38",
          3625 => x"73",
          3626 => x"81",
          3627 => x"ae",
          3628 => x"05",
          3629 => x"15",
          3630 => x"70",
          3631 => x"34",
          3632 => x"8a",
          3633 => x"38",
          3634 => x"05",
          3635 => x"81",
          3636 => x"17",
          3637 => x"12",
          3638 => x"34",
          3639 => x"9c",
          3640 => x"e8",
          3641 => x"f8",
          3642 => x"0c",
          3643 => x"e7",
          3644 => x"f8",
          3645 => x"17",
          3646 => x"51",
          3647 => x"81",
          3648 => x"84",
          3649 => x"3d",
          3650 => x"3d",
          3651 => x"08",
          3652 => x"61",
          3653 => x"55",
          3654 => x"2e",
          3655 => x"55",
          3656 => x"2e",
          3657 => x"80",
          3658 => x"94",
          3659 => x"1c",
          3660 => x"81",
          3661 => x"61",
          3662 => x"56",
          3663 => x"2e",
          3664 => x"83",
          3665 => x"73",
          3666 => x"70",
          3667 => x"25",
          3668 => x"51",
          3669 => x"38",
          3670 => x"0c",
          3671 => x"51",
          3672 => x"26",
          3673 => x"80",
          3674 => x"34",
          3675 => x"51",
          3676 => x"81",
          3677 => x"55",
          3678 => x"91",
          3679 => x"1d",
          3680 => x"8b",
          3681 => x"79",
          3682 => x"3f",
          3683 => x"57",
          3684 => x"55",
          3685 => x"2e",
          3686 => x"80",
          3687 => x"18",
          3688 => x"1a",
          3689 => x"70",
          3690 => x"2a",
          3691 => x"07",
          3692 => x"5a",
          3693 => x"8c",
          3694 => x"54",
          3695 => x"81",
          3696 => x"39",
          3697 => x"70",
          3698 => x"2a",
          3699 => x"75",
          3700 => x"8c",
          3701 => x"2e",
          3702 => x"a0",
          3703 => x"38",
          3704 => x"0c",
          3705 => x"76",
          3706 => x"38",
          3707 => x"b8",
          3708 => x"70",
          3709 => x"5a",
          3710 => x"76",
          3711 => x"38",
          3712 => x"70",
          3713 => x"dc",
          3714 => x"72",
          3715 => x"80",
          3716 => x"51",
          3717 => x"73",
          3718 => x"38",
          3719 => x"18",
          3720 => x"1a",
          3721 => x"55",
          3722 => x"2e",
          3723 => x"83",
          3724 => x"73",
          3725 => x"70",
          3726 => x"25",
          3727 => x"51",
          3728 => x"38",
          3729 => x"75",
          3730 => x"81",
          3731 => x"81",
          3732 => x"27",
          3733 => x"73",
          3734 => x"38",
          3735 => x"70",
          3736 => x"32",
          3737 => x"80",
          3738 => x"2a",
          3739 => x"56",
          3740 => x"81",
          3741 => x"57",
          3742 => x"f5",
          3743 => x"2b",
          3744 => x"25",
          3745 => x"80",
          3746 => x"e6",
          3747 => x"57",
          3748 => x"e6",
          3749 => x"f8",
          3750 => x"2e",
          3751 => x"18",
          3752 => x"1a",
          3753 => x"56",
          3754 => x"3f",
          3755 => x"08",
          3756 => x"e8",
          3757 => x"54",
          3758 => x"80",
          3759 => x"17",
          3760 => x"34",
          3761 => x"11",
          3762 => x"74",
          3763 => x"75",
          3764 => x"f8",
          3765 => x"3f",
          3766 => x"08",
          3767 => x"9f",
          3768 => x"99",
          3769 => x"e0",
          3770 => x"ff",
          3771 => x"79",
          3772 => x"74",
          3773 => x"57",
          3774 => x"77",
          3775 => x"76",
          3776 => x"38",
          3777 => x"73",
          3778 => x"09",
          3779 => x"38",
          3780 => x"84",
          3781 => x"27",
          3782 => x"39",
          3783 => x"f2",
          3784 => x"80",
          3785 => x"54",
          3786 => x"34",
          3787 => x"58",
          3788 => x"f2",
          3789 => x"f8",
          3790 => x"81",
          3791 => x"80",
          3792 => x"1b",
          3793 => x"51",
          3794 => x"81",
          3795 => x"56",
          3796 => x"08",
          3797 => x"9c",
          3798 => x"33",
          3799 => x"80",
          3800 => x"38",
          3801 => x"bf",
          3802 => x"86",
          3803 => x"15",
          3804 => x"2a",
          3805 => x"51",
          3806 => x"92",
          3807 => x"79",
          3808 => x"e4",
          3809 => x"f8",
          3810 => x"2e",
          3811 => x"52",
          3812 => x"ba",
          3813 => x"39",
          3814 => x"33",
          3815 => x"80",
          3816 => x"74",
          3817 => x"81",
          3818 => x"38",
          3819 => x"70",
          3820 => x"82",
          3821 => x"54",
          3822 => x"96",
          3823 => x"06",
          3824 => x"2e",
          3825 => x"ff",
          3826 => x"1c",
          3827 => x"80",
          3828 => x"81",
          3829 => x"ba",
          3830 => x"b6",
          3831 => x"2a",
          3832 => x"51",
          3833 => x"38",
          3834 => x"70",
          3835 => x"81",
          3836 => x"55",
          3837 => x"e1",
          3838 => x"08",
          3839 => x"1d",
          3840 => x"7c",
          3841 => x"3f",
          3842 => x"08",
          3843 => x"fa",
          3844 => x"81",
          3845 => x"8f",
          3846 => x"f6",
          3847 => x"5b",
          3848 => x"70",
          3849 => x"59",
          3850 => x"73",
          3851 => x"c6",
          3852 => x"81",
          3853 => x"70",
          3854 => x"52",
          3855 => x"8d",
          3856 => x"38",
          3857 => x"09",
          3858 => x"a5",
          3859 => x"d0",
          3860 => x"ff",
          3861 => x"53",
          3862 => x"91",
          3863 => x"73",
          3864 => x"d0",
          3865 => x"71",
          3866 => x"f7",
          3867 => x"81",
          3868 => x"55",
          3869 => x"55",
          3870 => x"81",
          3871 => x"74",
          3872 => x"56",
          3873 => x"12",
          3874 => x"70",
          3875 => x"38",
          3876 => x"81",
          3877 => x"51",
          3878 => x"51",
          3879 => x"89",
          3880 => x"70",
          3881 => x"53",
          3882 => x"70",
          3883 => x"51",
          3884 => x"09",
          3885 => x"38",
          3886 => x"38",
          3887 => x"77",
          3888 => x"70",
          3889 => x"2a",
          3890 => x"07",
          3891 => x"51",
          3892 => x"8f",
          3893 => x"84",
          3894 => x"83",
          3895 => x"94",
          3896 => x"74",
          3897 => x"38",
          3898 => x"0c",
          3899 => x"86",
          3900 => x"8c",
          3901 => x"81",
          3902 => x"8c",
          3903 => x"fa",
          3904 => x"56",
          3905 => x"17",
          3906 => x"b0",
          3907 => x"52",
          3908 => x"e0",
          3909 => x"81",
          3910 => x"81",
          3911 => x"b2",
          3912 => x"b4",
          3913 => x"c8",
          3914 => x"ff",
          3915 => x"55",
          3916 => x"d5",
          3917 => x"06",
          3918 => x"80",
          3919 => x"33",
          3920 => x"81",
          3921 => x"81",
          3922 => x"81",
          3923 => x"eb",
          3924 => x"70",
          3925 => x"07",
          3926 => x"73",
          3927 => x"81",
          3928 => x"81",
          3929 => x"83",
          3930 => x"88",
          3931 => x"16",
          3932 => x"3f",
          3933 => x"08",
          3934 => x"c8",
          3935 => x"9d",
          3936 => x"81",
          3937 => x"81",
          3938 => x"e0",
          3939 => x"f8",
          3940 => x"81",
          3941 => x"80",
          3942 => x"82",
          3943 => x"f8",
          3944 => x"3d",
          3945 => x"3d",
          3946 => x"84",
          3947 => x"05",
          3948 => x"80",
          3949 => x"51",
          3950 => x"81",
          3951 => x"58",
          3952 => x"0b",
          3953 => x"08",
          3954 => x"38",
          3955 => x"08",
          3956 => x"f8",
          3957 => x"08",
          3958 => x"56",
          3959 => x"86",
          3960 => x"75",
          3961 => x"fe",
          3962 => x"54",
          3963 => x"2e",
          3964 => x"14",
          3965 => x"ca",
          3966 => x"c8",
          3967 => x"06",
          3968 => x"54",
          3969 => x"38",
          3970 => x"86",
          3971 => x"82",
          3972 => x"06",
          3973 => x"56",
          3974 => x"38",
          3975 => x"80",
          3976 => x"81",
          3977 => x"52",
          3978 => x"51",
          3979 => x"81",
          3980 => x"81",
          3981 => x"81",
          3982 => x"83",
          3983 => x"87",
          3984 => x"2e",
          3985 => x"82",
          3986 => x"06",
          3987 => x"56",
          3988 => x"38",
          3989 => x"74",
          3990 => x"a3",
          3991 => x"c8",
          3992 => x"06",
          3993 => x"2e",
          3994 => x"80",
          3995 => x"3d",
          3996 => x"83",
          3997 => x"15",
          3998 => x"53",
          3999 => x"8d",
          4000 => x"15",
          4001 => x"3f",
          4002 => x"08",
          4003 => x"70",
          4004 => x"0c",
          4005 => x"16",
          4006 => x"80",
          4007 => x"80",
          4008 => x"54",
          4009 => x"84",
          4010 => x"5b",
          4011 => x"80",
          4012 => x"7a",
          4013 => x"fc",
          4014 => x"f8",
          4015 => x"ff",
          4016 => x"77",
          4017 => x"81",
          4018 => x"76",
          4019 => x"81",
          4020 => x"2e",
          4021 => x"8d",
          4022 => x"26",
          4023 => x"bf",
          4024 => x"f4",
          4025 => x"c8",
          4026 => x"ff",
          4027 => x"84",
          4028 => x"81",
          4029 => x"38",
          4030 => x"51",
          4031 => x"81",
          4032 => x"83",
          4033 => x"58",
          4034 => x"80",
          4035 => x"db",
          4036 => x"f8",
          4037 => x"77",
          4038 => x"80",
          4039 => x"82",
          4040 => x"c4",
          4041 => x"11",
          4042 => x"06",
          4043 => x"8d",
          4044 => x"26",
          4045 => x"74",
          4046 => x"78",
          4047 => x"c1",
          4048 => x"59",
          4049 => x"15",
          4050 => x"2e",
          4051 => x"13",
          4052 => x"72",
          4053 => x"38",
          4054 => x"eb",
          4055 => x"14",
          4056 => x"3f",
          4057 => x"08",
          4058 => x"c8",
          4059 => x"23",
          4060 => x"57",
          4061 => x"83",
          4062 => x"c7",
          4063 => x"d8",
          4064 => x"c8",
          4065 => x"ff",
          4066 => x"8d",
          4067 => x"14",
          4068 => x"3f",
          4069 => x"08",
          4070 => x"14",
          4071 => x"3f",
          4072 => x"08",
          4073 => x"06",
          4074 => x"72",
          4075 => x"97",
          4076 => x"22",
          4077 => x"84",
          4078 => x"5a",
          4079 => x"83",
          4080 => x"14",
          4081 => x"79",
          4082 => x"93",
          4083 => x"f8",
          4084 => x"81",
          4085 => x"80",
          4086 => x"38",
          4087 => x"08",
          4088 => x"ff",
          4089 => x"38",
          4090 => x"83",
          4091 => x"83",
          4092 => x"74",
          4093 => x"85",
          4094 => x"89",
          4095 => x"76",
          4096 => x"c3",
          4097 => x"70",
          4098 => x"7b",
          4099 => x"73",
          4100 => x"17",
          4101 => x"ac",
          4102 => x"55",
          4103 => x"09",
          4104 => x"38",
          4105 => x"51",
          4106 => x"81",
          4107 => x"83",
          4108 => x"53",
          4109 => x"82",
          4110 => x"82",
          4111 => x"e0",
          4112 => x"ab",
          4113 => x"c8",
          4114 => x"0c",
          4115 => x"53",
          4116 => x"56",
          4117 => x"81",
          4118 => x"13",
          4119 => x"74",
          4120 => x"82",
          4121 => x"74",
          4122 => x"81",
          4123 => x"06",
          4124 => x"83",
          4125 => x"2a",
          4126 => x"72",
          4127 => x"26",
          4128 => x"ff",
          4129 => x"0c",
          4130 => x"15",
          4131 => x"0b",
          4132 => x"76",
          4133 => x"81",
          4134 => x"38",
          4135 => x"51",
          4136 => x"81",
          4137 => x"83",
          4138 => x"53",
          4139 => x"09",
          4140 => x"f9",
          4141 => x"52",
          4142 => x"b8",
          4143 => x"c8",
          4144 => x"38",
          4145 => x"08",
          4146 => x"84",
          4147 => x"d8",
          4148 => x"f8",
          4149 => x"ff",
          4150 => x"72",
          4151 => x"2e",
          4152 => x"80",
          4153 => x"14",
          4154 => x"3f",
          4155 => x"08",
          4156 => x"a4",
          4157 => x"81",
          4158 => x"84",
          4159 => x"d7",
          4160 => x"f8",
          4161 => x"8a",
          4162 => x"2e",
          4163 => x"9d",
          4164 => x"14",
          4165 => x"3f",
          4166 => x"08",
          4167 => x"84",
          4168 => x"d7",
          4169 => x"f8",
          4170 => x"15",
          4171 => x"34",
          4172 => x"22",
          4173 => x"72",
          4174 => x"23",
          4175 => x"23",
          4176 => x"15",
          4177 => x"75",
          4178 => x"0c",
          4179 => x"04",
          4180 => x"77",
          4181 => x"73",
          4182 => x"38",
          4183 => x"72",
          4184 => x"38",
          4185 => x"71",
          4186 => x"38",
          4187 => x"84",
          4188 => x"52",
          4189 => x"09",
          4190 => x"38",
          4191 => x"51",
          4192 => x"81",
          4193 => x"81",
          4194 => x"88",
          4195 => x"08",
          4196 => x"39",
          4197 => x"73",
          4198 => x"74",
          4199 => x"0c",
          4200 => x"04",
          4201 => x"02",
          4202 => x"7a",
          4203 => x"fc",
          4204 => x"f4",
          4205 => x"54",
          4206 => x"f8",
          4207 => x"bc",
          4208 => x"c8",
          4209 => x"81",
          4210 => x"70",
          4211 => x"73",
          4212 => x"38",
          4213 => x"78",
          4214 => x"2e",
          4215 => x"74",
          4216 => x"0c",
          4217 => x"80",
          4218 => x"80",
          4219 => x"70",
          4220 => x"51",
          4221 => x"81",
          4222 => x"54",
          4223 => x"c8",
          4224 => x"0d",
          4225 => x"0d",
          4226 => x"05",
          4227 => x"33",
          4228 => x"54",
          4229 => x"84",
          4230 => x"bf",
          4231 => x"98",
          4232 => x"53",
          4233 => x"05",
          4234 => x"fa",
          4235 => x"c8",
          4236 => x"f8",
          4237 => x"a4",
          4238 => x"68",
          4239 => x"70",
          4240 => x"c6",
          4241 => x"c8",
          4242 => x"f8",
          4243 => x"38",
          4244 => x"05",
          4245 => x"2b",
          4246 => x"80",
          4247 => x"86",
          4248 => x"06",
          4249 => x"2e",
          4250 => x"74",
          4251 => x"38",
          4252 => x"09",
          4253 => x"38",
          4254 => x"f8",
          4255 => x"c8",
          4256 => x"39",
          4257 => x"33",
          4258 => x"73",
          4259 => x"77",
          4260 => x"81",
          4261 => x"73",
          4262 => x"38",
          4263 => x"bc",
          4264 => x"07",
          4265 => x"b4",
          4266 => x"2a",
          4267 => x"51",
          4268 => x"2e",
          4269 => x"62",
          4270 => x"e8",
          4271 => x"f8",
          4272 => x"82",
          4273 => x"52",
          4274 => x"51",
          4275 => x"62",
          4276 => x"8b",
          4277 => x"53",
          4278 => x"51",
          4279 => x"80",
          4280 => x"05",
          4281 => x"3f",
          4282 => x"0b",
          4283 => x"75",
          4284 => x"f1",
          4285 => x"11",
          4286 => x"80",
          4287 => x"97",
          4288 => x"51",
          4289 => x"81",
          4290 => x"55",
          4291 => x"08",
          4292 => x"b7",
          4293 => x"c4",
          4294 => x"05",
          4295 => x"2a",
          4296 => x"51",
          4297 => x"80",
          4298 => x"84",
          4299 => x"39",
          4300 => x"70",
          4301 => x"54",
          4302 => x"a9",
          4303 => x"06",
          4304 => x"2e",
          4305 => x"55",
          4306 => x"73",
          4307 => x"d6",
          4308 => x"f8",
          4309 => x"ff",
          4310 => x"0c",
          4311 => x"f8",
          4312 => x"f8",
          4313 => x"2a",
          4314 => x"51",
          4315 => x"2e",
          4316 => x"80",
          4317 => x"7a",
          4318 => x"a0",
          4319 => x"a4",
          4320 => x"53",
          4321 => x"e6",
          4322 => x"f8",
          4323 => x"f8",
          4324 => x"1b",
          4325 => x"05",
          4326 => x"d3",
          4327 => x"c8",
          4328 => x"c8",
          4329 => x"0c",
          4330 => x"56",
          4331 => x"84",
          4332 => x"90",
          4333 => x"0b",
          4334 => x"80",
          4335 => x"0c",
          4336 => x"1a",
          4337 => x"2a",
          4338 => x"51",
          4339 => x"2e",
          4340 => x"81",
          4341 => x"80",
          4342 => x"38",
          4343 => x"08",
          4344 => x"8a",
          4345 => x"89",
          4346 => x"59",
          4347 => x"76",
          4348 => x"d7",
          4349 => x"f8",
          4350 => x"81",
          4351 => x"81",
          4352 => x"82",
          4353 => x"c8",
          4354 => x"09",
          4355 => x"38",
          4356 => x"78",
          4357 => x"30",
          4358 => x"80",
          4359 => x"77",
          4360 => x"38",
          4361 => x"06",
          4362 => x"c3",
          4363 => x"1a",
          4364 => x"38",
          4365 => x"06",
          4366 => x"2e",
          4367 => x"52",
          4368 => x"a6",
          4369 => x"c8",
          4370 => x"82",
          4371 => x"75",
          4372 => x"f8",
          4373 => x"9c",
          4374 => x"39",
          4375 => x"74",
          4376 => x"f8",
          4377 => x"3d",
          4378 => x"3d",
          4379 => x"65",
          4380 => x"5d",
          4381 => x"0c",
          4382 => x"05",
          4383 => x"f9",
          4384 => x"f8",
          4385 => x"81",
          4386 => x"8a",
          4387 => x"33",
          4388 => x"2e",
          4389 => x"56",
          4390 => x"90",
          4391 => x"06",
          4392 => x"74",
          4393 => x"b6",
          4394 => x"82",
          4395 => x"34",
          4396 => x"aa",
          4397 => x"91",
          4398 => x"56",
          4399 => x"8c",
          4400 => x"1a",
          4401 => x"74",
          4402 => x"38",
          4403 => x"80",
          4404 => x"38",
          4405 => x"70",
          4406 => x"56",
          4407 => x"b2",
          4408 => x"11",
          4409 => x"77",
          4410 => x"5b",
          4411 => x"38",
          4412 => x"88",
          4413 => x"8f",
          4414 => x"08",
          4415 => x"d5",
          4416 => x"f8",
          4417 => x"81",
          4418 => x"9f",
          4419 => x"2e",
          4420 => x"74",
          4421 => x"98",
          4422 => x"7e",
          4423 => x"3f",
          4424 => x"08",
          4425 => x"83",
          4426 => x"c8",
          4427 => x"89",
          4428 => x"77",
          4429 => x"d6",
          4430 => x"7f",
          4431 => x"58",
          4432 => x"75",
          4433 => x"75",
          4434 => x"77",
          4435 => x"7c",
          4436 => x"33",
          4437 => x"3f",
          4438 => x"08",
          4439 => x"7e",
          4440 => x"56",
          4441 => x"2e",
          4442 => x"16",
          4443 => x"55",
          4444 => x"94",
          4445 => x"53",
          4446 => x"b0",
          4447 => x"31",
          4448 => x"05",
          4449 => x"3f",
          4450 => x"56",
          4451 => x"9c",
          4452 => x"19",
          4453 => x"06",
          4454 => x"31",
          4455 => x"76",
          4456 => x"7b",
          4457 => x"08",
          4458 => x"d1",
          4459 => x"f8",
          4460 => x"81",
          4461 => x"94",
          4462 => x"ff",
          4463 => x"05",
          4464 => x"cf",
          4465 => x"76",
          4466 => x"17",
          4467 => x"1e",
          4468 => x"18",
          4469 => x"5e",
          4470 => x"39",
          4471 => x"81",
          4472 => x"90",
          4473 => x"f2",
          4474 => x"63",
          4475 => x"40",
          4476 => x"7e",
          4477 => x"fc",
          4478 => x"51",
          4479 => x"81",
          4480 => x"55",
          4481 => x"08",
          4482 => x"18",
          4483 => x"80",
          4484 => x"74",
          4485 => x"39",
          4486 => x"70",
          4487 => x"81",
          4488 => x"56",
          4489 => x"80",
          4490 => x"38",
          4491 => x"0b",
          4492 => x"82",
          4493 => x"39",
          4494 => x"19",
          4495 => x"83",
          4496 => x"18",
          4497 => x"56",
          4498 => x"27",
          4499 => x"09",
          4500 => x"2e",
          4501 => x"94",
          4502 => x"83",
          4503 => x"56",
          4504 => x"38",
          4505 => x"22",
          4506 => x"89",
          4507 => x"55",
          4508 => x"75",
          4509 => x"18",
          4510 => x"9c",
          4511 => x"85",
          4512 => x"08",
          4513 => x"d7",
          4514 => x"f8",
          4515 => x"81",
          4516 => x"80",
          4517 => x"38",
          4518 => x"ff",
          4519 => x"ff",
          4520 => x"38",
          4521 => x"0c",
          4522 => x"85",
          4523 => x"19",
          4524 => x"b0",
          4525 => x"19",
          4526 => x"81",
          4527 => x"74",
          4528 => x"3f",
          4529 => x"08",
          4530 => x"98",
          4531 => x"7e",
          4532 => x"3f",
          4533 => x"08",
          4534 => x"d2",
          4535 => x"c8",
          4536 => x"89",
          4537 => x"78",
          4538 => x"d5",
          4539 => x"7f",
          4540 => x"58",
          4541 => x"75",
          4542 => x"75",
          4543 => x"78",
          4544 => x"7c",
          4545 => x"33",
          4546 => x"3f",
          4547 => x"08",
          4548 => x"7e",
          4549 => x"78",
          4550 => x"74",
          4551 => x"38",
          4552 => x"b0",
          4553 => x"31",
          4554 => x"05",
          4555 => x"51",
          4556 => x"7e",
          4557 => x"83",
          4558 => x"89",
          4559 => x"db",
          4560 => x"08",
          4561 => x"26",
          4562 => x"51",
          4563 => x"81",
          4564 => x"fd",
          4565 => x"77",
          4566 => x"55",
          4567 => x"0c",
          4568 => x"83",
          4569 => x"80",
          4570 => x"55",
          4571 => x"83",
          4572 => x"9c",
          4573 => x"7e",
          4574 => x"3f",
          4575 => x"08",
          4576 => x"75",
          4577 => x"94",
          4578 => x"ff",
          4579 => x"05",
          4580 => x"3f",
          4581 => x"0b",
          4582 => x"7b",
          4583 => x"08",
          4584 => x"76",
          4585 => x"08",
          4586 => x"1c",
          4587 => x"08",
          4588 => x"5c",
          4589 => x"83",
          4590 => x"74",
          4591 => x"fd",
          4592 => x"18",
          4593 => x"07",
          4594 => x"19",
          4595 => x"75",
          4596 => x"0c",
          4597 => x"04",
          4598 => x"7a",
          4599 => x"05",
          4600 => x"56",
          4601 => x"81",
          4602 => x"57",
          4603 => x"08",
          4604 => x"90",
          4605 => x"86",
          4606 => x"06",
          4607 => x"73",
          4608 => x"e9",
          4609 => x"08",
          4610 => x"cc",
          4611 => x"f8",
          4612 => x"81",
          4613 => x"80",
          4614 => x"16",
          4615 => x"33",
          4616 => x"55",
          4617 => x"34",
          4618 => x"53",
          4619 => x"08",
          4620 => x"3f",
          4621 => x"52",
          4622 => x"c9",
          4623 => x"88",
          4624 => x"96",
          4625 => x"f0",
          4626 => x"92",
          4627 => x"ca",
          4628 => x"81",
          4629 => x"34",
          4630 => x"df",
          4631 => x"c8",
          4632 => x"33",
          4633 => x"55",
          4634 => x"17",
          4635 => x"f8",
          4636 => x"3d",
          4637 => x"3d",
          4638 => x"52",
          4639 => x"3f",
          4640 => x"08",
          4641 => x"c8",
          4642 => x"86",
          4643 => x"52",
          4644 => x"bc",
          4645 => x"c8",
          4646 => x"f8",
          4647 => x"38",
          4648 => x"08",
          4649 => x"81",
          4650 => x"86",
          4651 => x"ff",
          4652 => x"3d",
          4653 => x"3f",
          4654 => x"0b",
          4655 => x"08",
          4656 => x"81",
          4657 => x"81",
          4658 => x"80",
          4659 => x"f8",
          4660 => x"3d",
          4661 => x"3d",
          4662 => x"93",
          4663 => x"52",
          4664 => x"e9",
          4665 => x"f8",
          4666 => x"81",
          4667 => x"80",
          4668 => x"58",
          4669 => x"3d",
          4670 => x"e0",
          4671 => x"f8",
          4672 => x"81",
          4673 => x"bc",
          4674 => x"c7",
          4675 => x"98",
          4676 => x"73",
          4677 => x"38",
          4678 => x"12",
          4679 => x"39",
          4680 => x"33",
          4681 => x"70",
          4682 => x"55",
          4683 => x"2e",
          4684 => x"7f",
          4685 => x"54",
          4686 => x"81",
          4687 => x"94",
          4688 => x"39",
          4689 => x"08",
          4690 => x"81",
          4691 => x"85",
          4692 => x"f8",
          4693 => x"3d",
          4694 => x"3d",
          4695 => x"5b",
          4696 => x"34",
          4697 => x"3d",
          4698 => x"52",
          4699 => x"e8",
          4700 => x"f8",
          4701 => x"81",
          4702 => x"82",
          4703 => x"43",
          4704 => x"11",
          4705 => x"58",
          4706 => x"80",
          4707 => x"38",
          4708 => x"3d",
          4709 => x"d5",
          4710 => x"f8",
          4711 => x"81",
          4712 => x"82",
          4713 => x"52",
          4714 => x"c8",
          4715 => x"c8",
          4716 => x"f8",
          4717 => x"c1",
          4718 => x"7b",
          4719 => x"3f",
          4720 => x"08",
          4721 => x"74",
          4722 => x"3f",
          4723 => x"08",
          4724 => x"c8",
          4725 => x"38",
          4726 => x"51",
          4727 => x"81",
          4728 => x"57",
          4729 => x"08",
          4730 => x"52",
          4731 => x"f2",
          4732 => x"f8",
          4733 => x"a6",
          4734 => x"74",
          4735 => x"3f",
          4736 => x"08",
          4737 => x"c8",
          4738 => x"cc",
          4739 => x"2e",
          4740 => x"86",
          4741 => x"81",
          4742 => x"81",
          4743 => x"3d",
          4744 => x"52",
          4745 => x"c9",
          4746 => x"3d",
          4747 => x"11",
          4748 => x"5a",
          4749 => x"2e",
          4750 => x"b9",
          4751 => x"16",
          4752 => x"33",
          4753 => x"73",
          4754 => x"16",
          4755 => x"26",
          4756 => x"75",
          4757 => x"38",
          4758 => x"05",
          4759 => x"6f",
          4760 => x"ff",
          4761 => x"55",
          4762 => x"74",
          4763 => x"38",
          4764 => x"11",
          4765 => x"74",
          4766 => x"39",
          4767 => x"09",
          4768 => x"38",
          4769 => x"11",
          4770 => x"74",
          4771 => x"81",
          4772 => x"70",
          4773 => x"e6",
          4774 => x"08",
          4775 => x"5c",
          4776 => x"73",
          4777 => x"38",
          4778 => x"1a",
          4779 => x"55",
          4780 => x"38",
          4781 => x"73",
          4782 => x"38",
          4783 => x"76",
          4784 => x"74",
          4785 => x"33",
          4786 => x"05",
          4787 => x"15",
          4788 => x"ba",
          4789 => x"05",
          4790 => x"ff",
          4791 => x"06",
          4792 => x"57",
          4793 => x"18",
          4794 => x"54",
          4795 => x"70",
          4796 => x"34",
          4797 => x"ee",
          4798 => x"34",
          4799 => x"c8",
          4800 => x"0d",
          4801 => x"0d",
          4802 => x"3d",
          4803 => x"71",
          4804 => x"ec",
          4805 => x"f8",
          4806 => x"81",
          4807 => x"82",
          4808 => x"15",
          4809 => x"82",
          4810 => x"15",
          4811 => x"76",
          4812 => x"90",
          4813 => x"81",
          4814 => x"06",
          4815 => x"72",
          4816 => x"56",
          4817 => x"54",
          4818 => x"17",
          4819 => x"78",
          4820 => x"38",
          4821 => x"22",
          4822 => x"59",
          4823 => x"78",
          4824 => x"76",
          4825 => x"51",
          4826 => x"3f",
          4827 => x"08",
          4828 => x"54",
          4829 => x"53",
          4830 => x"3f",
          4831 => x"08",
          4832 => x"38",
          4833 => x"75",
          4834 => x"18",
          4835 => x"31",
          4836 => x"57",
          4837 => x"b1",
          4838 => x"08",
          4839 => x"38",
          4840 => x"51",
          4841 => x"81",
          4842 => x"54",
          4843 => x"08",
          4844 => x"9a",
          4845 => x"c8",
          4846 => x"81",
          4847 => x"f8",
          4848 => x"16",
          4849 => x"16",
          4850 => x"2e",
          4851 => x"76",
          4852 => x"dc",
          4853 => x"31",
          4854 => x"18",
          4855 => x"90",
          4856 => x"81",
          4857 => x"06",
          4858 => x"56",
          4859 => x"9a",
          4860 => x"74",
          4861 => x"3f",
          4862 => x"08",
          4863 => x"c8",
          4864 => x"81",
          4865 => x"56",
          4866 => x"52",
          4867 => x"84",
          4868 => x"c8",
          4869 => x"ff",
          4870 => x"81",
          4871 => x"38",
          4872 => x"98",
          4873 => x"a6",
          4874 => x"16",
          4875 => x"39",
          4876 => x"16",
          4877 => x"75",
          4878 => x"53",
          4879 => x"aa",
          4880 => x"79",
          4881 => x"3f",
          4882 => x"08",
          4883 => x"0b",
          4884 => x"82",
          4885 => x"39",
          4886 => x"16",
          4887 => x"bb",
          4888 => x"2a",
          4889 => x"08",
          4890 => x"15",
          4891 => x"15",
          4892 => x"90",
          4893 => x"16",
          4894 => x"33",
          4895 => x"53",
          4896 => x"34",
          4897 => x"06",
          4898 => x"2e",
          4899 => x"9c",
          4900 => x"85",
          4901 => x"16",
          4902 => x"72",
          4903 => x"0c",
          4904 => x"04",
          4905 => x"79",
          4906 => x"75",
          4907 => x"8a",
          4908 => x"89",
          4909 => x"52",
          4910 => x"05",
          4911 => x"3f",
          4912 => x"08",
          4913 => x"c8",
          4914 => x"38",
          4915 => x"7a",
          4916 => x"d8",
          4917 => x"f8",
          4918 => x"81",
          4919 => x"80",
          4920 => x"16",
          4921 => x"2b",
          4922 => x"74",
          4923 => x"86",
          4924 => x"84",
          4925 => x"06",
          4926 => x"73",
          4927 => x"38",
          4928 => x"52",
          4929 => x"da",
          4930 => x"c8",
          4931 => x"0c",
          4932 => x"14",
          4933 => x"23",
          4934 => x"51",
          4935 => x"81",
          4936 => x"55",
          4937 => x"09",
          4938 => x"38",
          4939 => x"39",
          4940 => x"84",
          4941 => x"0c",
          4942 => x"81",
          4943 => x"89",
          4944 => x"fc",
          4945 => x"87",
          4946 => x"53",
          4947 => x"e7",
          4948 => x"f8",
          4949 => x"38",
          4950 => x"08",
          4951 => x"3d",
          4952 => x"3d",
          4953 => x"89",
          4954 => x"54",
          4955 => x"54",
          4956 => x"81",
          4957 => x"53",
          4958 => x"08",
          4959 => x"74",
          4960 => x"f8",
          4961 => x"73",
          4962 => x"3f",
          4963 => x"08",
          4964 => x"39",
          4965 => x"08",
          4966 => x"d3",
          4967 => x"f8",
          4968 => x"81",
          4969 => x"84",
          4970 => x"06",
          4971 => x"53",
          4972 => x"f8",
          4973 => x"38",
          4974 => x"51",
          4975 => x"72",
          4976 => x"cf",
          4977 => x"f8",
          4978 => x"32",
          4979 => x"72",
          4980 => x"70",
          4981 => x"08",
          4982 => x"54",
          4983 => x"f8",
          4984 => x"3d",
          4985 => x"3d",
          4986 => x"80",
          4987 => x"70",
          4988 => x"52",
          4989 => x"3f",
          4990 => x"08",
          4991 => x"c8",
          4992 => x"64",
          4993 => x"d6",
          4994 => x"f8",
          4995 => x"81",
          4996 => x"a0",
          4997 => x"cb",
          4998 => x"98",
          4999 => x"73",
          5000 => x"38",
          5001 => x"39",
          5002 => x"88",
          5003 => x"75",
          5004 => x"3f",
          5005 => x"c8",
          5006 => x"0d",
          5007 => x"0d",
          5008 => x"5c",
          5009 => x"3d",
          5010 => x"93",
          5011 => x"d6",
          5012 => x"c8",
          5013 => x"f8",
          5014 => x"80",
          5015 => x"0c",
          5016 => x"11",
          5017 => x"90",
          5018 => x"56",
          5019 => x"74",
          5020 => x"75",
          5021 => x"e4",
          5022 => x"81",
          5023 => x"5b",
          5024 => x"81",
          5025 => x"75",
          5026 => x"73",
          5027 => x"81",
          5028 => x"82",
          5029 => x"76",
          5030 => x"f0",
          5031 => x"f4",
          5032 => x"c8",
          5033 => x"d1",
          5034 => x"c8",
          5035 => x"ce",
          5036 => x"c8",
          5037 => x"81",
          5038 => x"07",
          5039 => x"05",
          5040 => x"53",
          5041 => x"98",
          5042 => x"26",
          5043 => x"f9",
          5044 => x"08",
          5045 => x"08",
          5046 => x"98",
          5047 => x"81",
          5048 => x"58",
          5049 => x"3f",
          5050 => x"08",
          5051 => x"c8",
          5052 => x"38",
          5053 => x"77",
          5054 => x"5d",
          5055 => x"74",
          5056 => x"81",
          5057 => x"b4",
          5058 => x"bb",
          5059 => x"f8",
          5060 => x"ff",
          5061 => x"30",
          5062 => x"1b",
          5063 => x"5b",
          5064 => x"39",
          5065 => x"ff",
          5066 => x"81",
          5067 => x"f0",
          5068 => x"30",
          5069 => x"1b",
          5070 => x"5b",
          5071 => x"83",
          5072 => x"58",
          5073 => x"92",
          5074 => x"0c",
          5075 => x"12",
          5076 => x"33",
          5077 => x"54",
          5078 => x"34",
          5079 => x"c8",
          5080 => x"0d",
          5081 => x"0d",
          5082 => x"fc",
          5083 => x"52",
          5084 => x"3f",
          5085 => x"08",
          5086 => x"c8",
          5087 => x"38",
          5088 => x"56",
          5089 => x"38",
          5090 => x"70",
          5091 => x"81",
          5092 => x"55",
          5093 => x"80",
          5094 => x"38",
          5095 => x"54",
          5096 => x"08",
          5097 => x"38",
          5098 => x"81",
          5099 => x"53",
          5100 => x"52",
          5101 => x"8c",
          5102 => x"c8",
          5103 => x"19",
          5104 => x"c9",
          5105 => x"08",
          5106 => x"ff",
          5107 => x"81",
          5108 => x"ff",
          5109 => x"06",
          5110 => x"56",
          5111 => x"08",
          5112 => x"81",
          5113 => x"82",
          5114 => x"75",
          5115 => x"54",
          5116 => x"08",
          5117 => x"27",
          5118 => x"17",
          5119 => x"f8",
          5120 => x"76",
          5121 => x"3f",
          5122 => x"08",
          5123 => x"08",
          5124 => x"90",
          5125 => x"c0",
          5126 => x"90",
          5127 => x"80",
          5128 => x"75",
          5129 => x"75",
          5130 => x"f8",
          5131 => x"3d",
          5132 => x"3d",
          5133 => x"a0",
          5134 => x"05",
          5135 => x"51",
          5136 => x"81",
          5137 => x"55",
          5138 => x"08",
          5139 => x"78",
          5140 => x"08",
          5141 => x"70",
          5142 => x"ae",
          5143 => x"c8",
          5144 => x"f8",
          5145 => x"db",
          5146 => x"fb",
          5147 => x"85",
          5148 => x"06",
          5149 => x"86",
          5150 => x"c7",
          5151 => x"2b",
          5152 => x"24",
          5153 => x"02",
          5154 => x"33",
          5155 => x"58",
          5156 => x"76",
          5157 => x"6b",
          5158 => x"cc",
          5159 => x"f8",
          5160 => x"84",
          5161 => x"06",
          5162 => x"73",
          5163 => x"d4",
          5164 => x"81",
          5165 => x"94",
          5166 => x"81",
          5167 => x"5a",
          5168 => x"08",
          5169 => x"8a",
          5170 => x"54",
          5171 => x"81",
          5172 => x"55",
          5173 => x"08",
          5174 => x"81",
          5175 => x"52",
          5176 => x"e5",
          5177 => x"c8",
          5178 => x"f8",
          5179 => x"38",
          5180 => x"cf",
          5181 => x"c8",
          5182 => x"88",
          5183 => x"c8",
          5184 => x"38",
          5185 => x"c2",
          5186 => x"c8",
          5187 => x"c8",
          5188 => x"81",
          5189 => x"07",
          5190 => x"55",
          5191 => x"2e",
          5192 => x"80",
          5193 => x"80",
          5194 => x"77",
          5195 => x"3f",
          5196 => x"08",
          5197 => x"38",
          5198 => x"ba",
          5199 => x"f8",
          5200 => x"74",
          5201 => x"0c",
          5202 => x"04",
          5203 => x"82",
          5204 => x"c0",
          5205 => x"3d",
          5206 => x"3f",
          5207 => x"08",
          5208 => x"c8",
          5209 => x"38",
          5210 => x"52",
          5211 => x"52",
          5212 => x"3f",
          5213 => x"08",
          5214 => x"c8",
          5215 => x"88",
          5216 => x"39",
          5217 => x"08",
          5218 => x"81",
          5219 => x"38",
          5220 => x"05",
          5221 => x"2a",
          5222 => x"55",
          5223 => x"81",
          5224 => x"5a",
          5225 => x"3d",
          5226 => x"c1",
          5227 => x"f8",
          5228 => x"55",
          5229 => x"c8",
          5230 => x"87",
          5231 => x"c8",
          5232 => x"09",
          5233 => x"38",
          5234 => x"f8",
          5235 => x"2e",
          5236 => x"86",
          5237 => x"81",
          5238 => x"81",
          5239 => x"f8",
          5240 => x"78",
          5241 => x"3f",
          5242 => x"08",
          5243 => x"c8",
          5244 => x"38",
          5245 => x"52",
          5246 => x"ff",
          5247 => x"78",
          5248 => x"b4",
          5249 => x"54",
          5250 => x"15",
          5251 => x"b2",
          5252 => x"ca",
          5253 => x"b6",
          5254 => x"53",
          5255 => x"53",
          5256 => x"3f",
          5257 => x"b4",
          5258 => x"d4",
          5259 => x"b6",
          5260 => x"54",
          5261 => x"d5",
          5262 => x"53",
          5263 => x"11",
          5264 => x"d7",
          5265 => x"81",
          5266 => x"34",
          5267 => x"a4",
          5268 => x"c8",
          5269 => x"f8",
          5270 => x"38",
          5271 => x"0a",
          5272 => x"05",
          5273 => x"d0",
          5274 => x"64",
          5275 => x"c9",
          5276 => x"54",
          5277 => x"15",
          5278 => x"81",
          5279 => x"34",
          5280 => x"b8",
          5281 => x"f8",
          5282 => x"8b",
          5283 => x"75",
          5284 => x"ff",
          5285 => x"73",
          5286 => x"0c",
          5287 => x"04",
          5288 => x"a9",
          5289 => x"51",
          5290 => x"82",
          5291 => x"ff",
          5292 => x"a9",
          5293 => x"ee",
          5294 => x"c8",
          5295 => x"f8",
          5296 => x"d3",
          5297 => x"a9",
          5298 => x"9d",
          5299 => x"58",
          5300 => x"81",
          5301 => x"55",
          5302 => x"08",
          5303 => x"02",
          5304 => x"33",
          5305 => x"54",
          5306 => x"82",
          5307 => x"53",
          5308 => x"52",
          5309 => x"88",
          5310 => x"b4",
          5311 => x"53",
          5312 => x"3d",
          5313 => x"ff",
          5314 => x"aa",
          5315 => x"73",
          5316 => x"3f",
          5317 => x"08",
          5318 => x"c8",
          5319 => x"63",
          5320 => x"81",
          5321 => x"65",
          5322 => x"2e",
          5323 => x"55",
          5324 => x"81",
          5325 => x"84",
          5326 => x"06",
          5327 => x"73",
          5328 => x"3f",
          5329 => x"08",
          5330 => x"c8",
          5331 => x"38",
          5332 => x"53",
          5333 => x"95",
          5334 => x"16",
          5335 => x"87",
          5336 => x"05",
          5337 => x"34",
          5338 => x"70",
          5339 => x"81",
          5340 => x"55",
          5341 => x"74",
          5342 => x"73",
          5343 => x"78",
          5344 => x"83",
          5345 => x"16",
          5346 => x"2a",
          5347 => x"51",
          5348 => x"80",
          5349 => x"38",
          5350 => x"80",
          5351 => x"52",
          5352 => x"be",
          5353 => x"c8",
          5354 => x"51",
          5355 => x"3f",
          5356 => x"f8",
          5357 => x"2e",
          5358 => x"81",
          5359 => x"52",
          5360 => x"b5",
          5361 => x"f8",
          5362 => x"80",
          5363 => x"58",
          5364 => x"c8",
          5365 => x"38",
          5366 => x"54",
          5367 => x"09",
          5368 => x"38",
          5369 => x"52",
          5370 => x"af",
          5371 => x"81",
          5372 => x"34",
          5373 => x"f8",
          5374 => x"38",
          5375 => x"ca",
          5376 => x"c8",
          5377 => x"f8",
          5378 => x"38",
          5379 => x"b5",
          5380 => x"f8",
          5381 => x"74",
          5382 => x"0c",
          5383 => x"04",
          5384 => x"02",
          5385 => x"33",
          5386 => x"80",
          5387 => x"57",
          5388 => x"95",
          5389 => x"52",
          5390 => x"d2",
          5391 => x"f8",
          5392 => x"81",
          5393 => x"80",
          5394 => x"5a",
          5395 => x"3d",
          5396 => x"c9",
          5397 => x"f8",
          5398 => x"81",
          5399 => x"b8",
          5400 => x"cf",
          5401 => x"a0",
          5402 => x"55",
          5403 => x"75",
          5404 => x"71",
          5405 => x"33",
          5406 => x"74",
          5407 => x"57",
          5408 => x"8b",
          5409 => x"54",
          5410 => x"15",
          5411 => x"ff",
          5412 => x"81",
          5413 => x"55",
          5414 => x"c8",
          5415 => x"0d",
          5416 => x"0d",
          5417 => x"53",
          5418 => x"05",
          5419 => x"51",
          5420 => x"81",
          5421 => x"55",
          5422 => x"08",
          5423 => x"76",
          5424 => x"93",
          5425 => x"51",
          5426 => x"81",
          5427 => x"55",
          5428 => x"08",
          5429 => x"80",
          5430 => x"81",
          5431 => x"86",
          5432 => x"38",
          5433 => x"86",
          5434 => x"90",
          5435 => x"54",
          5436 => x"ff",
          5437 => x"76",
          5438 => x"83",
          5439 => x"51",
          5440 => x"3f",
          5441 => x"08",
          5442 => x"f8",
          5443 => x"3d",
          5444 => x"3d",
          5445 => x"5c",
          5446 => x"98",
          5447 => x"52",
          5448 => x"d1",
          5449 => x"f8",
          5450 => x"f8",
          5451 => x"70",
          5452 => x"08",
          5453 => x"51",
          5454 => x"80",
          5455 => x"38",
          5456 => x"06",
          5457 => x"80",
          5458 => x"38",
          5459 => x"5f",
          5460 => x"3d",
          5461 => x"ff",
          5462 => x"81",
          5463 => x"57",
          5464 => x"08",
          5465 => x"74",
          5466 => x"c3",
          5467 => x"f8",
          5468 => x"81",
          5469 => x"bf",
          5470 => x"c8",
          5471 => x"c8",
          5472 => x"59",
          5473 => x"81",
          5474 => x"56",
          5475 => x"33",
          5476 => x"16",
          5477 => x"27",
          5478 => x"56",
          5479 => x"80",
          5480 => x"80",
          5481 => x"ff",
          5482 => x"70",
          5483 => x"56",
          5484 => x"e8",
          5485 => x"76",
          5486 => x"81",
          5487 => x"80",
          5488 => x"57",
          5489 => x"78",
          5490 => x"51",
          5491 => x"2e",
          5492 => x"73",
          5493 => x"38",
          5494 => x"08",
          5495 => x"b1",
          5496 => x"f8",
          5497 => x"81",
          5498 => x"a7",
          5499 => x"33",
          5500 => x"c3",
          5501 => x"2e",
          5502 => x"e4",
          5503 => x"2e",
          5504 => x"56",
          5505 => x"05",
          5506 => x"e3",
          5507 => x"c8",
          5508 => x"76",
          5509 => x"0c",
          5510 => x"04",
          5511 => x"82",
          5512 => x"ff",
          5513 => x"9d",
          5514 => x"fa",
          5515 => x"c8",
          5516 => x"c8",
          5517 => x"81",
          5518 => x"83",
          5519 => x"53",
          5520 => x"3d",
          5521 => x"ff",
          5522 => x"73",
          5523 => x"70",
          5524 => x"52",
          5525 => x"9f",
          5526 => x"bc",
          5527 => x"74",
          5528 => x"6d",
          5529 => x"70",
          5530 => x"af",
          5531 => x"f8",
          5532 => x"2e",
          5533 => x"70",
          5534 => x"57",
          5535 => x"fd",
          5536 => x"c8",
          5537 => x"8d",
          5538 => x"2b",
          5539 => x"81",
          5540 => x"86",
          5541 => x"c8",
          5542 => x"9f",
          5543 => x"ff",
          5544 => x"54",
          5545 => x"8a",
          5546 => x"70",
          5547 => x"06",
          5548 => x"ff",
          5549 => x"38",
          5550 => x"15",
          5551 => x"80",
          5552 => x"74",
          5553 => x"d8",
          5554 => x"89",
          5555 => x"c8",
          5556 => x"81",
          5557 => x"88",
          5558 => x"26",
          5559 => x"39",
          5560 => x"86",
          5561 => x"81",
          5562 => x"ff",
          5563 => x"38",
          5564 => x"54",
          5565 => x"81",
          5566 => x"81",
          5567 => x"78",
          5568 => x"5a",
          5569 => x"6d",
          5570 => x"81",
          5571 => x"57",
          5572 => x"9f",
          5573 => x"38",
          5574 => x"54",
          5575 => x"81",
          5576 => x"b1",
          5577 => x"2e",
          5578 => x"a7",
          5579 => x"15",
          5580 => x"54",
          5581 => x"09",
          5582 => x"38",
          5583 => x"76",
          5584 => x"41",
          5585 => x"52",
          5586 => x"52",
          5587 => x"b3",
          5588 => x"c8",
          5589 => x"f8",
          5590 => x"f7",
          5591 => x"74",
          5592 => x"e5",
          5593 => x"c8",
          5594 => x"f8",
          5595 => x"38",
          5596 => x"38",
          5597 => x"74",
          5598 => x"39",
          5599 => x"08",
          5600 => x"81",
          5601 => x"38",
          5602 => x"74",
          5603 => x"38",
          5604 => x"51",
          5605 => x"3f",
          5606 => x"08",
          5607 => x"c8",
          5608 => x"a0",
          5609 => x"c8",
          5610 => x"51",
          5611 => x"3f",
          5612 => x"0b",
          5613 => x"8b",
          5614 => x"67",
          5615 => x"a7",
          5616 => x"81",
          5617 => x"34",
          5618 => x"ad",
          5619 => x"f8",
          5620 => x"73",
          5621 => x"f8",
          5622 => x"3d",
          5623 => x"3d",
          5624 => x"02",
          5625 => x"cb",
          5626 => x"3d",
          5627 => x"72",
          5628 => x"5a",
          5629 => x"81",
          5630 => x"58",
          5631 => x"08",
          5632 => x"91",
          5633 => x"77",
          5634 => x"7c",
          5635 => x"38",
          5636 => x"59",
          5637 => x"90",
          5638 => x"81",
          5639 => x"06",
          5640 => x"73",
          5641 => x"54",
          5642 => x"82",
          5643 => x"39",
          5644 => x"8b",
          5645 => x"11",
          5646 => x"2b",
          5647 => x"54",
          5648 => x"fe",
          5649 => x"ff",
          5650 => x"70",
          5651 => x"07",
          5652 => x"f8",
          5653 => x"8c",
          5654 => x"40",
          5655 => x"55",
          5656 => x"88",
          5657 => x"08",
          5658 => x"38",
          5659 => x"77",
          5660 => x"56",
          5661 => x"51",
          5662 => x"3f",
          5663 => x"55",
          5664 => x"08",
          5665 => x"38",
          5666 => x"f8",
          5667 => x"2e",
          5668 => x"81",
          5669 => x"ff",
          5670 => x"38",
          5671 => x"08",
          5672 => x"16",
          5673 => x"2e",
          5674 => x"87",
          5675 => x"74",
          5676 => x"74",
          5677 => x"81",
          5678 => x"38",
          5679 => x"ff",
          5680 => x"2e",
          5681 => x"7b",
          5682 => x"80",
          5683 => x"81",
          5684 => x"81",
          5685 => x"06",
          5686 => x"56",
          5687 => x"52",
          5688 => x"af",
          5689 => x"f8",
          5690 => x"81",
          5691 => x"80",
          5692 => x"81",
          5693 => x"56",
          5694 => x"d3",
          5695 => x"ff",
          5696 => x"7c",
          5697 => x"55",
          5698 => x"b3",
          5699 => x"1b",
          5700 => x"1b",
          5701 => x"33",
          5702 => x"54",
          5703 => x"34",
          5704 => x"fe",
          5705 => x"08",
          5706 => x"74",
          5707 => x"75",
          5708 => x"16",
          5709 => x"33",
          5710 => x"73",
          5711 => x"77",
          5712 => x"f8",
          5713 => x"3d",
          5714 => x"3d",
          5715 => x"02",
          5716 => x"eb",
          5717 => x"3d",
          5718 => x"59",
          5719 => x"8b",
          5720 => x"81",
          5721 => x"24",
          5722 => x"81",
          5723 => x"84",
          5724 => x"f8",
          5725 => x"51",
          5726 => x"2e",
          5727 => x"75",
          5728 => x"c8",
          5729 => x"06",
          5730 => x"7e",
          5731 => x"d0",
          5732 => x"c8",
          5733 => x"06",
          5734 => x"56",
          5735 => x"74",
          5736 => x"76",
          5737 => x"81",
          5738 => x"8a",
          5739 => x"b2",
          5740 => x"fc",
          5741 => x"52",
          5742 => x"a4",
          5743 => x"f8",
          5744 => x"38",
          5745 => x"80",
          5746 => x"74",
          5747 => x"26",
          5748 => x"15",
          5749 => x"74",
          5750 => x"38",
          5751 => x"80",
          5752 => x"84",
          5753 => x"92",
          5754 => x"80",
          5755 => x"38",
          5756 => x"06",
          5757 => x"2e",
          5758 => x"56",
          5759 => x"78",
          5760 => x"89",
          5761 => x"2b",
          5762 => x"43",
          5763 => x"38",
          5764 => x"30",
          5765 => x"77",
          5766 => x"91",
          5767 => x"c2",
          5768 => x"f8",
          5769 => x"52",
          5770 => x"a4",
          5771 => x"56",
          5772 => x"08",
          5773 => x"77",
          5774 => x"77",
          5775 => x"c8",
          5776 => x"45",
          5777 => x"bf",
          5778 => x"8e",
          5779 => x"26",
          5780 => x"74",
          5781 => x"48",
          5782 => x"75",
          5783 => x"38",
          5784 => x"81",
          5785 => x"fa",
          5786 => x"2a",
          5787 => x"56",
          5788 => x"2e",
          5789 => x"87",
          5790 => x"82",
          5791 => x"38",
          5792 => x"55",
          5793 => x"83",
          5794 => x"81",
          5795 => x"56",
          5796 => x"80",
          5797 => x"38",
          5798 => x"83",
          5799 => x"06",
          5800 => x"78",
          5801 => x"91",
          5802 => x"0b",
          5803 => x"22",
          5804 => x"80",
          5805 => x"74",
          5806 => x"38",
          5807 => x"56",
          5808 => x"17",
          5809 => x"57",
          5810 => x"2e",
          5811 => x"75",
          5812 => x"79",
          5813 => x"fe",
          5814 => x"81",
          5815 => x"84",
          5816 => x"05",
          5817 => x"5e",
          5818 => x"80",
          5819 => x"c8",
          5820 => x"8a",
          5821 => x"fd",
          5822 => x"75",
          5823 => x"38",
          5824 => x"78",
          5825 => x"8c",
          5826 => x"0b",
          5827 => x"22",
          5828 => x"80",
          5829 => x"74",
          5830 => x"38",
          5831 => x"56",
          5832 => x"17",
          5833 => x"57",
          5834 => x"2e",
          5835 => x"75",
          5836 => x"79",
          5837 => x"fe",
          5838 => x"81",
          5839 => x"10",
          5840 => x"81",
          5841 => x"9f",
          5842 => x"38",
          5843 => x"f8",
          5844 => x"81",
          5845 => x"05",
          5846 => x"2a",
          5847 => x"56",
          5848 => x"17",
          5849 => x"81",
          5850 => x"60",
          5851 => x"65",
          5852 => x"12",
          5853 => x"30",
          5854 => x"74",
          5855 => x"59",
          5856 => x"7d",
          5857 => x"81",
          5858 => x"76",
          5859 => x"41",
          5860 => x"76",
          5861 => x"90",
          5862 => x"62",
          5863 => x"51",
          5864 => x"26",
          5865 => x"75",
          5866 => x"31",
          5867 => x"65",
          5868 => x"fe",
          5869 => x"81",
          5870 => x"58",
          5871 => x"09",
          5872 => x"38",
          5873 => x"08",
          5874 => x"26",
          5875 => x"78",
          5876 => x"79",
          5877 => x"78",
          5878 => x"86",
          5879 => x"82",
          5880 => x"06",
          5881 => x"83",
          5882 => x"81",
          5883 => x"27",
          5884 => x"8f",
          5885 => x"55",
          5886 => x"26",
          5887 => x"59",
          5888 => x"62",
          5889 => x"74",
          5890 => x"38",
          5891 => x"88",
          5892 => x"c8",
          5893 => x"26",
          5894 => x"86",
          5895 => x"1a",
          5896 => x"79",
          5897 => x"38",
          5898 => x"80",
          5899 => x"2e",
          5900 => x"83",
          5901 => x"9f",
          5902 => x"8b",
          5903 => x"06",
          5904 => x"74",
          5905 => x"84",
          5906 => x"52",
          5907 => x"a2",
          5908 => x"53",
          5909 => x"52",
          5910 => x"a2",
          5911 => x"80",
          5912 => x"51",
          5913 => x"3f",
          5914 => x"34",
          5915 => x"ff",
          5916 => x"1b",
          5917 => x"a2",
          5918 => x"90",
          5919 => x"83",
          5920 => x"70",
          5921 => x"80",
          5922 => x"55",
          5923 => x"ff",
          5924 => x"66",
          5925 => x"ff",
          5926 => x"38",
          5927 => x"ff",
          5928 => x"1b",
          5929 => x"f2",
          5930 => x"74",
          5931 => x"51",
          5932 => x"3f",
          5933 => x"1c",
          5934 => x"98",
          5935 => x"a0",
          5936 => x"ff",
          5937 => x"51",
          5938 => x"3f",
          5939 => x"1b",
          5940 => x"e4",
          5941 => x"2e",
          5942 => x"80",
          5943 => x"88",
          5944 => x"80",
          5945 => x"ff",
          5946 => x"7c",
          5947 => x"51",
          5948 => x"3f",
          5949 => x"1b",
          5950 => x"bc",
          5951 => x"b0",
          5952 => x"a0",
          5953 => x"52",
          5954 => x"ff",
          5955 => x"ff",
          5956 => x"c0",
          5957 => x"0b",
          5958 => x"34",
          5959 => x"e6",
          5960 => x"c7",
          5961 => x"39",
          5962 => x"0a",
          5963 => x"51",
          5964 => x"3f",
          5965 => x"ff",
          5966 => x"1b",
          5967 => x"da",
          5968 => x"0b",
          5969 => x"a9",
          5970 => x"34",
          5971 => x"e6",
          5972 => x"1b",
          5973 => x"8f",
          5974 => x"d5",
          5975 => x"1b",
          5976 => x"ff",
          5977 => x"81",
          5978 => x"7a",
          5979 => x"ff",
          5980 => x"81",
          5981 => x"c8",
          5982 => x"38",
          5983 => x"09",
          5984 => x"ee",
          5985 => x"60",
          5986 => x"7a",
          5987 => x"ff",
          5988 => x"84",
          5989 => x"52",
          5990 => x"9f",
          5991 => x"8b",
          5992 => x"52",
          5993 => x"9f",
          5994 => x"8a",
          5995 => x"52",
          5996 => x"51",
          5997 => x"3f",
          5998 => x"83",
          5999 => x"ff",
          6000 => x"82",
          6001 => x"1b",
          6002 => x"ec",
          6003 => x"d5",
          6004 => x"ff",
          6005 => x"75",
          6006 => x"05",
          6007 => x"7e",
          6008 => x"e5",
          6009 => x"60",
          6010 => x"52",
          6011 => x"9a",
          6012 => x"53",
          6013 => x"51",
          6014 => x"3f",
          6015 => x"58",
          6016 => x"09",
          6017 => x"38",
          6018 => x"51",
          6019 => x"3f",
          6020 => x"1b",
          6021 => x"a0",
          6022 => x"52",
          6023 => x"91",
          6024 => x"ff",
          6025 => x"81",
          6026 => x"f8",
          6027 => x"7a",
          6028 => x"84",
          6029 => x"61",
          6030 => x"26",
          6031 => x"57",
          6032 => x"53",
          6033 => x"51",
          6034 => x"3f",
          6035 => x"08",
          6036 => x"84",
          6037 => x"f8",
          6038 => x"7a",
          6039 => x"aa",
          6040 => x"75",
          6041 => x"56",
          6042 => x"81",
          6043 => x"80",
          6044 => x"38",
          6045 => x"83",
          6046 => x"63",
          6047 => x"74",
          6048 => x"38",
          6049 => x"54",
          6050 => x"52",
          6051 => x"99",
          6052 => x"f8",
          6053 => x"c1",
          6054 => x"75",
          6055 => x"56",
          6056 => x"8c",
          6057 => x"2e",
          6058 => x"56",
          6059 => x"ff",
          6060 => x"84",
          6061 => x"2e",
          6062 => x"56",
          6063 => x"58",
          6064 => x"38",
          6065 => x"77",
          6066 => x"ff",
          6067 => x"82",
          6068 => x"78",
          6069 => x"c2",
          6070 => x"1b",
          6071 => x"34",
          6072 => x"16",
          6073 => x"82",
          6074 => x"83",
          6075 => x"84",
          6076 => x"67",
          6077 => x"fd",
          6078 => x"51",
          6079 => x"3f",
          6080 => x"16",
          6081 => x"c8",
          6082 => x"bf",
          6083 => x"86",
          6084 => x"f8",
          6085 => x"16",
          6086 => x"83",
          6087 => x"ff",
          6088 => x"66",
          6089 => x"1b",
          6090 => x"8c",
          6091 => x"77",
          6092 => x"7e",
          6093 => x"91",
          6094 => x"81",
          6095 => x"a2",
          6096 => x"80",
          6097 => x"ff",
          6098 => x"81",
          6099 => x"c8",
          6100 => x"89",
          6101 => x"8a",
          6102 => x"86",
          6103 => x"c8",
          6104 => x"81",
          6105 => x"99",
          6106 => x"f5",
          6107 => x"60",
          6108 => x"79",
          6109 => x"5a",
          6110 => x"78",
          6111 => x"8d",
          6112 => x"55",
          6113 => x"fc",
          6114 => x"51",
          6115 => x"7a",
          6116 => x"81",
          6117 => x"8c",
          6118 => x"74",
          6119 => x"38",
          6120 => x"81",
          6121 => x"81",
          6122 => x"8a",
          6123 => x"06",
          6124 => x"76",
          6125 => x"76",
          6126 => x"55",
          6127 => x"c8",
          6128 => x"0d",
          6129 => x"0d",
          6130 => x"05",
          6131 => x"59",
          6132 => x"2e",
          6133 => x"87",
          6134 => x"76",
          6135 => x"84",
          6136 => x"80",
          6137 => x"38",
          6138 => x"77",
          6139 => x"56",
          6140 => x"34",
          6141 => x"bb",
          6142 => x"38",
          6143 => x"05",
          6144 => x"8c",
          6145 => x"08",
          6146 => x"3f",
          6147 => x"70",
          6148 => x"07",
          6149 => x"30",
          6150 => x"56",
          6151 => x"0c",
          6152 => x"18",
          6153 => x"0d",
          6154 => x"0d",
          6155 => x"08",
          6156 => x"75",
          6157 => x"89",
          6158 => x"54",
          6159 => x"16",
          6160 => x"51",
          6161 => x"81",
          6162 => x"91",
          6163 => x"08",
          6164 => x"81",
          6165 => x"88",
          6166 => x"83",
          6167 => x"74",
          6168 => x"0c",
          6169 => x"04",
          6170 => x"75",
          6171 => x"53",
          6172 => x"51",
          6173 => x"3f",
          6174 => x"85",
          6175 => x"ea",
          6176 => x"80",
          6177 => x"6a",
          6178 => x"70",
          6179 => x"d8",
          6180 => x"72",
          6181 => x"3f",
          6182 => x"8d",
          6183 => x"0d",
          6184 => x"0d",
          6185 => x"70",
          6186 => x"74",
          6187 => x"e1",
          6188 => x"77",
          6189 => x"85",
          6190 => x"80",
          6191 => x"33",
          6192 => x"2e",
          6193 => x"86",
          6194 => x"55",
          6195 => x"57",
          6196 => x"81",
          6197 => x"70",
          6198 => x"fe",
          6199 => x"81",
          6200 => x"81",
          6201 => x"54",
          6202 => x"08",
          6203 => x"db",
          6204 => x"f8",
          6205 => x"38",
          6206 => x"54",
          6207 => x"ff",
          6208 => x"17",
          6209 => x"06",
          6210 => x"77",
          6211 => x"ff",
          6212 => x"f8",
          6213 => x"3d",
          6214 => x"3d",
          6215 => x"71",
          6216 => x"8e",
          6217 => x"29",
          6218 => x"05",
          6219 => x"04",
          6220 => x"51",
          6221 => x"81",
          6222 => x"80",
          6223 => x"e9",
          6224 => x"f2",
          6225 => x"e8",
          6226 => x"39",
          6227 => x"51",
          6228 => x"81",
          6229 => x"80",
          6230 => x"ea",
          6231 => x"d6",
          6232 => x"ac",
          6233 => x"39",
          6234 => x"51",
          6235 => x"81",
          6236 => x"80",
          6237 => x"ea",
          6238 => x"39",
          6239 => x"51",
          6240 => x"eb",
          6241 => x"39",
          6242 => x"51",
          6243 => x"eb",
          6244 => x"39",
          6245 => x"51",
          6246 => x"ec",
          6247 => x"39",
          6248 => x"51",
          6249 => x"ec",
          6250 => x"39",
          6251 => x"51",
          6252 => x"ec",
          6253 => x"f2",
          6254 => x"3d",
          6255 => x"3d",
          6256 => x"56",
          6257 => x"e7",
          6258 => x"74",
          6259 => x"e8",
          6260 => x"39",
          6261 => x"74",
          6262 => x"d2",
          6263 => x"c8",
          6264 => x"51",
          6265 => x"3f",
          6266 => x"08",
          6267 => x"75",
          6268 => x"fc",
          6269 => x"d3",
          6270 => x"0d",
          6271 => x"0d",
          6272 => x"05",
          6273 => x"33",
          6274 => x"68",
          6275 => x"7a",
          6276 => x"51",
          6277 => x"78",
          6278 => x"ff",
          6279 => x"81",
          6280 => x"07",
          6281 => x"06",
          6282 => x"56",
          6283 => x"38",
          6284 => x"52",
          6285 => x"52",
          6286 => x"c9",
          6287 => x"c8",
          6288 => x"f8",
          6289 => x"38",
          6290 => x"08",
          6291 => x"88",
          6292 => x"c8",
          6293 => x"3d",
          6294 => x"84",
          6295 => x"52",
          6296 => x"86",
          6297 => x"c8",
          6298 => x"f8",
          6299 => x"38",
          6300 => x"80",
          6301 => x"74",
          6302 => x"59",
          6303 => x"96",
          6304 => x"51",
          6305 => x"76",
          6306 => x"07",
          6307 => x"30",
          6308 => x"72",
          6309 => x"51",
          6310 => x"2e",
          6311 => x"ed",
          6312 => x"c0",
          6313 => x"52",
          6314 => x"92",
          6315 => x"75",
          6316 => x"0c",
          6317 => x"04",
          6318 => x"7b",
          6319 => x"b3",
          6320 => x"58",
          6321 => x"53",
          6322 => x"51",
          6323 => x"81",
          6324 => x"a4",
          6325 => x"2e",
          6326 => x"81",
          6327 => x"98",
          6328 => x"7f",
          6329 => x"c8",
          6330 => x"7d",
          6331 => x"81",
          6332 => x"57",
          6333 => x"04",
          6334 => x"c8",
          6335 => x"0d",
          6336 => x"0d",
          6337 => x"02",
          6338 => x"cf",
          6339 => x"73",
          6340 => x"5f",
          6341 => x"5e",
          6342 => x"81",
          6343 => x"fe",
          6344 => x"81",
          6345 => x"fe",
          6346 => x"80",
          6347 => x"27",
          6348 => x"7b",
          6349 => x"38",
          6350 => x"a7",
          6351 => x"39",
          6352 => x"72",
          6353 => x"38",
          6354 => x"81",
          6355 => x"fe",
          6356 => x"89",
          6357 => x"c0",
          6358 => x"8b",
          6359 => x"55",
          6360 => x"74",
          6361 => x"7a",
          6362 => x"72",
          6363 => x"ed",
          6364 => x"f4",
          6365 => x"39",
          6366 => x"51",
          6367 => x"3f",
          6368 => x"a1",
          6369 => x"53",
          6370 => x"8e",
          6371 => x"52",
          6372 => x"51",
          6373 => x"3f",
          6374 => x"ed",
          6375 => x"ee",
          6376 => x"15",
          6377 => x"fe",
          6378 => x"ff",
          6379 => x"ed",
          6380 => x"ee",
          6381 => x"55",
          6382 => x"bc",
          6383 => x"70",
          6384 => x"80",
          6385 => x"27",
          6386 => x"56",
          6387 => x"74",
          6388 => x"81",
          6389 => x"06",
          6390 => x"06",
          6391 => x"80",
          6392 => x"73",
          6393 => x"85",
          6394 => x"83",
          6395 => x"fe",
          6396 => x"81",
          6397 => x"39",
          6398 => x"51",
          6399 => x"3f",
          6400 => x"1c",
          6401 => x"de",
          6402 => x"f8",
          6403 => x"2b",
          6404 => x"51",
          6405 => x"2e",
          6406 => x"ab",
          6407 => x"c0",
          6408 => x"c8",
          6409 => x"70",
          6410 => x"a0",
          6411 => x"72",
          6412 => x"30",
          6413 => x"73",
          6414 => x"51",
          6415 => x"57",
          6416 => x"73",
          6417 => x"76",
          6418 => x"81",
          6419 => x"80",
          6420 => x"7c",
          6421 => x"78",
          6422 => x"38",
          6423 => x"81",
          6424 => x"8f",
          6425 => x"fc",
          6426 => x"9b",
          6427 => x"ed",
          6428 => x"ed",
          6429 => x"fe",
          6430 => x"81",
          6431 => x"51",
          6432 => x"3f",
          6433 => x"54",
          6434 => x"53",
          6435 => x"33",
          6436 => x"80",
          6437 => x"b3",
          6438 => x"2e",
          6439 => x"e2",
          6440 => x"3d",
          6441 => x"3d",
          6442 => x"96",
          6443 => x"fe",
          6444 => x"81",
          6445 => x"bc",
          6446 => x"9c",
          6447 => x"b4",
          6448 => x"fe",
          6449 => x"72",
          6450 => x"81",
          6451 => x"71",
          6452 => x"38",
          6453 => x"d9",
          6454 => x"ee",
          6455 => x"db",
          6456 => x"51",
          6457 => x"3f",
          6458 => x"70",
          6459 => x"52",
          6460 => x"95",
          6461 => x"fe",
          6462 => x"81",
          6463 => x"fe",
          6464 => x"80",
          6465 => x"ec",
          6466 => x"2a",
          6467 => x"51",
          6468 => x"2e",
          6469 => x"51",
          6470 => x"3f",
          6471 => x"51",
          6472 => x"3f",
          6473 => x"d8",
          6474 => x"84",
          6475 => x"06",
          6476 => x"80",
          6477 => x"81",
          6478 => x"b8",
          6479 => x"ec",
          6480 => x"b0",
          6481 => x"fe",
          6482 => x"72",
          6483 => x"81",
          6484 => x"71",
          6485 => x"38",
          6486 => x"d8",
          6487 => x"ef",
          6488 => x"da",
          6489 => x"51",
          6490 => x"3f",
          6491 => x"70",
          6492 => x"52",
          6493 => x"95",
          6494 => x"fe",
          6495 => x"81",
          6496 => x"fe",
          6497 => x"80",
          6498 => x"e8",
          6499 => x"2a",
          6500 => x"51",
          6501 => x"2e",
          6502 => x"51",
          6503 => x"3f",
          6504 => x"51",
          6505 => x"3f",
          6506 => x"d7",
          6507 => x"88",
          6508 => x"06",
          6509 => x"80",
          6510 => x"81",
          6511 => x"b4",
          6512 => x"bc",
          6513 => x"ac",
          6514 => x"fe",
          6515 => x"fe",
          6516 => x"84",
          6517 => x"fb",
          6518 => x"02",
          6519 => x"05",
          6520 => x"56",
          6521 => x"75",
          6522 => x"e4",
          6523 => x"b4",
          6524 => x"a7",
          6525 => x"81",
          6526 => x"82",
          6527 => x"ff",
          6528 => x"81",
          6529 => x"30",
          6530 => x"c8",
          6531 => x"25",
          6532 => x"51",
          6533 => x"81",
          6534 => x"81",
          6535 => x"54",
          6536 => x"09",
          6537 => x"38",
          6538 => x"53",
          6539 => x"51",
          6540 => x"81",
          6541 => x"80",
          6542 => x"81",
          6543 => x"51",
          6544 => x"3f",
          6545 => x"8f",
          6546 => x"aa",
          6547 => x"81",
          6548 => x"81",
          6549 => x"54",
          6550 => x"09",
          6551 => x"38",
          6552 => x"51",
          6553 => x"3f",
          6554 => x"f8",
          6555 => x"3d",
          6556 => x"3d",
          6557 => x"71",
          6558 => x"0c",
          6559 => x"52",
          6560 => x"86",
          6561 => x"f8",
          6562 => x"ff",
          6563 => x"7d",
          6564 => x"06",
          6565 => x"f0",
          6566 => x"3d",
          6567 => x"fe",
          6568 => x"7c",
          6569 => x"81",
          6570 => x"ff",
          6571 => x"81",
          6572 => x"7d",
          6573 => x"81",
          6574 => x"8d",
          6575 => x"70",
          6576 => x"f0",
          6577 => x"e8",
          6578 => x"3d",
          6579 => x"80",
          6580 => x"51",
          6581 => x"b4",
          6582 => x"05",
          6583 => x"3f",
          6584 => x"08",
          6585 => x"90",
          6586 => x"78",
          6587 => x"87",
          6588 => x"80",
          6589 => x"38",
          6590 => x"81",
          6591 => x"bd",
          6592 => x"78",
          6593 => x"ba",
          6594 => x"2e",
          6595 => x"8a",
          6596 => x"80",
          6597 => x"a1",
          6598 => x"c0",
          6599 => x"38",
          6600 => x"82",
          6601 => x"d2",
          6602 => x"f9",
          6603 => x"38",
          6604 => x"24",
          6605 => x"80",
          6606 => x"98",
          6607 => x"f8",
          6608 => x"38",
          6609 => x"78",
          6610 => x"8a",
          6611 => x"81",
          6612 => x"38",
          6613 => x"2e",
          6614 => x"8a",
          6615 => x"81",
          6616 => x"8f",
          6617 => x"39",
          6618 => x"80",
          6619 => x"84",
          6620 => x"ee",
          6621 => x"f8",
          6622 => x"2e",
          6623 => x"b4",
          6624 => x"11",
          6625 => x"05",
          6626 => x"b4",
          6627 => x"c8",
          6628 => x"fe",
          6629 => x"3d",
          6630 => x"53",
          6631 => x"51",
          6632 => x"3f",
          6633 => x"08",
          6634 => x"f8",
          6635 => x"81",
          6636 => x"fe",
          6637 => x"63",
          6638 => x"79",
          6639 => x"f2",
          6640 => x"78",
          6641 => x"05",
          6642 => x"7a",
          6643 => x"81",
          6644 => x"3d",
          6645 => x"53",
          6646 => x"51",
          6647 => x"3f",
          6648 => x"08",
          6649 => x"da",
          6650 => x"fe",
          6651 => x"ff",
          6652 => x"fe",
          6653 => x"81",
          6654 => x"80",
          6655 => x"38",
          6656 => x"f8",
          6657 => x"84",
          6658 => x"ed",
          6659 => x"f8",
          6660 => x"2e",
          6661 => x"81",
          6662 => x"fe",
          6663 => x"63",
          6664 => x"27",
          6665 => x"61",
          6666 => x"81",
          6667 => x"79",
          6668 => x"05",
          6669 => x"b4",
          6670 => x"11",
          6671 => x"05",
          6672 => x"fc",
          6673 => x"c8",
          6674 => x"fc",
          6675 => x"3d",
          6676 => x"53",
          6677 => x"51",
          6678 => x"3f",
          6679 => x"08",
          6680 => x"de",
          6681 => x"fe",
          6682 => x"ff",
          6683 => x"fe",
          6684 => x"81",
          6685 => x"80",
          6686 => x"38",
          6687 => x"51",
          6688 => x"3f",
          6689 => x"63",
          6690 => x"61",
          6691 => x"33",
          6692 => x"78",
          6693 => x"38",
          6694 => x"54",
          6695 => x"79",
          6696 => x"f8",
          6697 => x"a3",
          6698 => x"62",
          6699 => x"5a",
          6700 => x"f1",
          6701 => x"bd",
          6702 => x"ff",
          6703 => x"ff",
          6704 => x"fe",
          6705 => x"81",
          6706 => x"80",
          6707 => x"f4",
          6708 => x"78",
          6709 => x"38",
          6710 => x"08",
          6711 => x"39",
          6712 => x"33",
          6713 => x"2e",
          6714 => x"f3",
          6715 => x"bc",
          6716 => x"8e",
          6717 => x"80",
          6718 => x"81",
          6719 => x"44",
          6720 => x"f4",
          6721 => x"78",
          6722 => x"38",
          6723 => x"08",
          6724 => x"81",
          6725 => x"59",
          6726 => x"88",
          6727 => x"e4",
          6728 => x"39",
          6729 => x"08",
          6730 => x"44",
          6731 => x"fc",
          6732 => x"84",
          6733 => x"eb",
          6734 => x"f8",
          6735 => x"de",
          6736 => x"8c",
          6737 => x"80",
          6738 => x"81",
          6739 => x"43",
          6740 => x"81",
          6741 => x"59",
          6742 => x"88",
          6743 => x"d0",
          6744 => x"39",
          6745 => x"33",
          6746 => x"2e",
          6747 => x"f3",
          6748 => x"aa",
          6749 => x"8f",
          6750 => x"80",
          6751 => x"81",
          6752 => x"43",
          6753 => x"f4",
          6754 => x"78",
          6755 => x"38",
          6756 => x"08",
          6757 => x"81",
          6758 => x"88",
          6759 => x"3d",
          6760 => x"53",
          6761 => x"51",
          6762 => x"3f",
          6763 => x"08",
          6764 => x"38",
          6765 => x"5c",
          6766 => x"83",
          6767 => x"7a",
          6768 => x"30",
          6769 => x"9f",
          6770 => x"06",
          6771 => x"5a",
          6772 => x"88",
          6773 => x"2e",
          6774 => x"42",
          6775 => x"51",
          6776 => x"3f",
          6777 => x"54",
          6778 => x"52",
          6779 => x"91",
          6780 => x"a4",
          6781 => x"ef",
          6782 => x"39",
          6783 => x"80",
          6784 => x"84",
          6785 => x"e9",
          6786 => x"f8",
          6787 => x"2e",
          6788 => x"b4",
          6789 => x"11",
          6790 => x"05",
          6791 => x"a0",
          6792 => x"c8",
          6793 => x"a5",
          6794 => x"02",
          6795 => x"33",
          6796 => x"81",
          6797 => x"3d",
          6798 => x"53",
          6799 => x"51",
          6800 => x"3f",
          6801 => x"08",
          6802 => x"f6",
          6803 => x"33",
          6804 => x"f1",
          6805 => x"e6",
          6806 => x"f8",
          6807 => x"fe",
          6808 => x"79",
          6809 => x"59",
          6810 => x"f8",
          6811 => x"79",
          6812 => x"b4",
          6813 => x"11",
          6814 => x"05",
          6815 => x"c0",
          6816 => x"c8",
          6817 => x"91",
          6818 => x"02",
          6819 => x"33",
          6820 => x"81",
          6821 => x"b5",
          6822 => x"bc",
          6823 => x"c7",
          6824 => x"39",
          6825 => x"f4",
          6826 => x"84",
          6827 => x"ea",
          6828 => x"f8",
          6829 => x"2e",
          6830 => x"b4",
          6831 => x"11",
          6832 => x"05",
          6833 => x"ea",
          6834 => x"c8",
          6835 => x"a6",
          6836 => x"02",
          6837 => x"79",
          6838 => x"5b",
          6839 => x"b4",
          6840 => x"11",
          6841 => x"05",
          6842 => x"c6",
          6843 => x"c8",
          6844 => x"f7",
          6845 => x"70",
          6846 => x"81",
          6847 => x"fe",
          6848 => x"80",
          6849 => x"51",
          6850 => x"3f",
          6851 => x"33",
          6852 => x"2e",
          6853 => x"78",
          6854 => x"38",
          6855 => x"41",
          6856 => x"3d",
          6857 => x"53",
          6858 => x"51",
          6859 => x"3f",
          6860 => x"08",
          6861 => x"38",
          6862 => x"be",
          6863 => x"70",
          6864 => x"23",
          6865 => x"ae",
          6866 => x"bc",
          6867 => x"97",
          6868 => x"39",
          6869 => x"f4",
          6870 => x"84",
          6871 => x"e8",
          6872 => x"f8",
          6873 => x"2e",
          6874 => x"b4",
          6875 => x"11",
          6876 => x"05",
          6877 => x"ba",
          6878 => x"c8",
          6879 => x"a1",
          6880 => x"71",
          6881 => x"84",
          6882 => x"3d",
          6883 => x"53",
          6884 => x"51",
          6885 => x"3f",
          6886 => x"08",
          6887 => x"a2",
          6888 => x"08",
          6889 => x"f1",
          6890 => x"e4",
          6891 => x"f8",
          6892 => x"fe",
          6893 => x"79",
          6894 => x"59",
          6895 => x"f6",
          6896 => x"79",
          6897 => x"b4",
          6898 => x"11",
          6899 => x"05",
          6900 => x"de",
          6901 => x"c8",
          6902 => x"8d",
          6903 => x"71",
          6904 => x"84",
          6905 => x"b9",
          6906 => x"bc",
          6907 => x"f7",
          6908 => x"39",
          6909 => x"80",
          6910 => x"84",
          6911 => x"e5",
          6912 => x"f8",
          6913 => x"2e",
          6914 => x"63",
          6915 => x"dc",
          6916 => x"b7",
          6917 => x"78",
          6918 => x"ff",
          6919 => x"ff",
          6920 => x"fe",
          6921 => x"81",
          6922 => x"80",
          6923 => x"38",
          6924 => x"f1",
          6925 => x"e3",
          6926 => x"59",
          6927 => x"f8",
          6928 => x"2e",
          6929 => x"81",
          6930 => x"52",
          6931 => x"51",
          6932 => x"3f",
          6933 => x"81",
          6934 => x"fe",
          6935 => x"fe",
          6936 => x"f4",
          6937 => x"f2",
          6938 => x"dc",
          6939 => x"59",
          6940 => x"fe",
          6941 => x"f4",
          6942 => x"45",
          6943 => x"78",
          6944 => x"be",
          6945 => x"06",
          6946 => x"2e",
          6947 => x"b4",
          6948 => x"05",
          6949 => x"8d",
          6950 => x"c8",
          6951 => x"5b",
          6952 => x"b2",
          6953 => x"24",
          6954 => x"81",
          6955 => x"80",
          6956 => x"83",
          6957 => x"80",
          6958 => x"f2",
          6959 => x"55",
          6960 => x"54",
          6961 => x"f2",
          6962 => x"3d",
          6963 => x"51",
          6964 => x"3f",
          6965 => x"f3",
          6966 => x"3d",
          6967 => x"51",
          6968 => x"3f",
          6969 => x"55",
          6970 => x"54",
          6971 => x"f2",
          6972 => x"3d",
          6973 => x"51",
          6974 => x"3f",
          6975 => x"54",
          6976 => x"f3",
          6977 => x"3d",
          6978 => x"51",
          6979 => x"3f",
          6980 => x"58",
          6981 => x"57",
          6982 => x"55",
          6983 => x"80",
          6984 => x"80",
          6985 => x"3d",
          6986 => x"51",
          6987 => x"81",
          6988 => x"81",
          6989 => x"09",
          6990 => x"72",
          6991 => x"51",
          6992 => x"80",
          6993 => x"26",
          6994 => x"5a",
          6995 => x"59",
          6996 => x"8d",
          6997 => x"70",
          6998 => x"5c",
          6999 => x"c0",
          7000 => x"32",
          7001 => x"07",
          7002 => x"38",
          7003 => x"09",
          7004 => x"ce",
          7005 => x"8c",
          7006 => x"cf",
          7007 => x"39",
          7008 => x"80",
          7009 => x"90",
          7010 => x"94",
          7011 => x"54",
          7012 => x"80",
          7013 => x"fe",
          7014 => x"81",
          7015 => x"90",
          7016 => x"55",
          7017 => x"80",
          7018 => x"fe",
          7019 => x"72",
          7020 => x"08",
          7021 => x"87",
          7022 => x"70",
          7023 => x"87",
          7024 => x"72",
          7025 => x"e6",
          7026 => x"c8",
          7027 => x"75",
          7028 => x"87",
          7029 => x"73",
          7030 => x"d2",
          7031 => x"f8",
          7032 => x"75",
          7033 => x"83",
          7034 => x"94",
          7035 => x"80",
          7036 => x"c0",
          7037 => x"a3",
          7038 => x"f8",
          7039 => x"8c",
          7040 => x"e0",
          7041 => x"b0",
          7042 => x"d7",
          7043 => x"9c",
          7044 => x"d3",
          7045 => x"a8",
          7046 => x"cb",
          7047 => x"a3",
          7048 => x"ba",
          7049 => x"ec",
          7050 => x"c6",
          7051 => x"00",
          7052 => x"ff",
          7053 => x"ff",
          7054 => x"ff",
          7055 => x"00",
          7056 => x"00",
          7057 => x"00",
          7058 => x"00",
          7059 => x"00",
          7060 => x"00",
          7061 => x"00",
          7062 => x"00",
          7063 => x"00",
          7064 => x"00",
          7065 => x"00",
          7066 => x"00",
          7067 => x"00",
          7068 => x"00",
          7069 => x"00",
          7070 => x"00",
          7071 => x"00",
          7072 => x"00",
          7073 => x"00",
          7074 => x"00",
          7075 => x"00",
          7076 => x"00",
          7077 => x"00",
          7078 => x"00",
          7079 => x"00",
          7080 => x"00",
          7081 => x"00",
          7082 => x"00",
          7083 => x"00",
          7084 => x"00",
          7085 => x"00",
          7086 => x"00",
          7087 => x"00",
          7088 => x"00",
          7089 => x"00",
          7090 => x"00",
          7091 => x"00",
          7092 => x"25",
          7093 => x"64",
          7094 => x"20",
          7095 => x"25",
          7096 => x"64",
          7097 => x"25",
          7098 => x"53",
          7099 => x"43",
          7100 => x"69",
          7101 => x"61",
          7102 => x"6e",
          7103 => x"20",
          7104 => x"6f",
          7105 => x"6f",
          7106 => x"6f",
          7107 => x"67",
          7108 => x"3a",
          7109 => x"76",
          7110 => x"73",
          7111 => x"70",
          7112 => x"65",
          7113 => x"64",
          7114 => x"20",
          7115 => x"57",
          7116 => x"44",
          7117 => x"20",
          7118 => x"30",
          7119 => x"25",
          7120 => x"29",
          7121 => x"20",
          7122 => x"53",
          7123 => x"4d",
          7124 => x"20",
          7125 => x"30",
          7126 => x"25",
          7127 => x"29",
          7128 => x"20",
          7129 => x"49",
          7130 => x"20",
          7131 => x"4d",
          7132 => x"30",
          7133 => x"25",
          7134 => x"29",
          7135 => x"20",
          7136 => x"42",
          7137 => x"20",
          7138 => x"20",
          7139 => x"30",
          7140 => x"25",
          7141 => x"29",
          7142 => x"20",
          7143 => x"52",
          7144 => x"20",
          7145 => x"20",
          7146 => x"30",
          7147 => x"25",
          7148 => x"29",
          7149 => x"20",
          7150 => x"53",
          7151 => x"41",
          7152 => x"20",
          7153 => x"65",
          7154 => x"65",
          7155 => x"25",
          7156 => x"29",
          7157 => x"20",
          7158 => x"54",
          7159 => x"52",
          7160 => x"20",
          7161 => x"69",
          7162 => x"73",
          7163 => x"25",
          7164 => x"29",
          7165 => x"20",
          7166 => x"49",
          7167 => x"20",
          7168 => x"4c",
          7169 => x"68",
          7170 => x"65",
          7171 => x"25",
          7172 => x"29",
          7173 => x"20",
          7174 => x"57",
          7175 => x"42",
          7176 => x"20",
          7177 => x"0a",
          7178 => x"20",
          7179 => x"57",
          7180 => x"32",
          7181 => x"20",
          7182 => x"49",
          7183 => x"4c",
          7184 => x"20",
          7185 => x"50",
          7186 => x"00",
          7187 => x"20",
          7188 => x"53",
          7189 => x"00",
          7190 => x"41",
          7191 => x"65",
          7192 => x"73",
          7193 => x"20",
          7194 => x"43",
          7195 => x"52",
          7196 => x"74",
          7197 => x"63",
          7198 => x"20",
          7199 => x"72",
          7200 => x"20",
          7201 => x"30",
          7202 => x"00",
          7203 => x"20",
          7204 => x"43",
          7205 => x"4d",
          7206 => x"72",
          7207 => x"74",
          7208 => x"20",
          7209 => x"72",
          7210 => x"20",
          7211 => x"30",
          7212 => x"00",
          7213 => x"20",
          7214 => x"53",
          7215 => x"6b",
          7216 => x"61",
          7217 => x"41",
          7218 => x"65",
          7219 => x"20",
          7220 => x"20",
          7221 => x"30",
          7222 => x"00",
          7223 => x"4d",
          7224 => x"3a",
          7225 => x"20",
          7226 => x"5a",
          7227 => x"49",
          7228 => x"20",
          7229 => x"20",
          7230 => x"20",
          7231 => x"20",
          7232 => x"20",
          7233 => x"30",
          7234 => x"00",
          7235 => x"20",
          7236 => x"53",
          7237 => x"65",
          7238 => x"6c",
          7239 => x"20",
          7240 => x"71",
          7241 => x"20",
          7242 => x"20",
          7243 => x"64",
          7244 => x"34",
          7245 => x"7a",
          7246 => x"20",
          7247 => x"53",
          7248 => x"4d",
          7249 => x"6f",
          7250 => x"46",
          7251 => x"20",
          7252 => x"20",
          7253 => x"20",
          7254 => x"64",
          7255 => x"34",
          7256 => x"7a",
          7257 => x"20",
          7258 => x"57",
          7259 => x"62",
          7260 => x"20",
          7261 => x"41",
          7262 => x"6c",
          7263 => x"20",
          7264 => x"71",
          7265 => x"64",
          7266 => x"34",
          7267 => x"7a",
          7268 => x"53",
          7269 => x"6c",
          7270 => x"4d",
          7271 => x"75",
          7272 => x"46",
          7273 => x"00",
          7274 => x"45",
          7275 => x"45",
          7276 => x"69",
          7277 => x"55",
          7278 => x"6f",
          7279 => x"68",
          7280 => x"6f",
          7281 => x"74",
          7282 => x"68",
          7283 => x"6f",
          7284 => x"68",
          7285 => x"00",
          7286 => x"21",
          7287 => x"25",
          7288 => x"20",
          7289 => x"0a",
          7290 => x"46",
          7291 => x"65",
          7292 => x"6f",
          7293 => x"73",
          7294 => x"74",
          7295 => x"68",
          7296 => x"6f",
          7297 => x"66",
          7298 => x"20",
          7299 => x"45",
          7300 => x"0a",
          7301 => x"43",
          7302 => x"6f",
          7303 => x"70",
          7304 => x"63",
          7305 => x"74",
          7306 => x"69",
          7307 => x"72",
          7308 => x"69",
          7309 => x"20",
          7310 => x"61",
          7311 => x"6e",
          7312 => x"00",
          7313 => x"00",
          7314 => x"01",
          7315 => x"00",
          7316 => x"00",
          7317 => x"01",
          7318 => x"00",
          7319 => x"00",
          7320 => x"04",
          7321 => x"00",
          7322 => x"00",
          7323 => x"04",
          7324 => x"00",
          7325 => x"00",
          7326 => x"04",
          7327 => x"00",
          7328 => x"00",
          7329 => x"04",
          7330 => x"00",
          7331 => x"00",
          7332 => x"04",
          7333 => x"00",
          7334 => x"00",
          7335 => x"03",
          7336 => x"00",
          7337 => x"00",
          7338 => x"03",
          7339 => x"00",
          7340 => x"00",
          7341 => x"03",
          7342 => x"00",
          7343 => x"00",
          7344 => x"03",
          7345 => x"00",
          7346 => x"1b",
          7347 => x"1b",
          7348 => x"1b",
          7349 => x"1b",
          7350 => x"1b",
          7351 => x"1b",
          7352 => x"1b",
          7353 => x"1b",
          7354 => x"1b",
          7355 => x"0d",
          7356 => x"08",
          7357 => x"53",
          7358 => x"22",
          7359 => x"3a",
          7360 => x"3e",
          7361 => x"7c",
          7362 => x"46",
          7363 => x"46",
          7364 => x"32",
          7365 => x"eb",
          7366 => x"53",
          7367 => x"35",
          7368 => x"4e",
          7369 => x"41",
          7370 => x"20",
          7371 => x"41",
          7372 => x"20",
          7373 => x"4e",
          7374 => x"41",
          7375 => x"20",
          7376 => x"41",
          7377 => x"20",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"80",
          7383 => x"8e",
          7384 => x"45",
          7385 => x"49",
          7386 => x"90",
          7387 => x"99",
          7388 => x"59",
          7389 => x"9c",
          7390 => x"41",
          7391 => x"a5",
          7392 => x"a8",
          7393 => x"ac",
          7394 => x"b0",
          7395 => x"b4",
          7396 => x"b8",
          7397 => x"bc",
          7398 => x"c0",
          7399 => x"c4",
          7400 => x"c8",
          7401 => x"cc",
          7402 => x"d0",
          7403 => x"d4",
          7404 => x"d8",
          7405 => x"dc",
          7406 => x"e0",
          7407 => x"e4",
          7408 => x"e8",
          7409 => x"ec",
          7410 => x"f0",
          7411 => x"f4",
          7412 => x"f8",
          7413 => x"fc",
          7414 => x"2b",
          7415 => x"3d",
          7416 => x"5c",
          7417 => x"3c",
          7418 => x"7f",
          7419 => x"00",
          7420 => x"00",
          7421 => x"01",
          7422 => x"00",
          7423 => x"00",
          7424 => x"00",
          7425 => x"00",
          7426 => x"00",
          7427 => x"64",
          7428 => x"74",
          7429 => x"64",
          7430 => x"74",
          7431 => x"66",
          7432 => x"74",
          7433 => x"66",
          7434 => x"64",
          7435 => x"66",
          7436 => x"63",
          7437 => x"6d",
          7438 => x"61",
          7439 => x"6d",
          7440 => x"79",
          7441 => x"6d",
          7442 => x"66",
          7443 => x"6d",
          7444 => x"70",
          7445 => x"6d",
          7446 => x"6d",
          7447 => x"6d",
          7448 => x"68",
          7449 => x"68",
          7450 => x"68",
          7451 => x"68",
          7452 => x"63",
          7453 => x"00",
          7454 => x"6a",
          7455 => x"72",
          7456 => x"61",
          7457 => x"72",
          7458 => x"74",
          7459 => x"69",
          7460 => x"00",
          7461 => x"74",
          7462 => x"00",
          7463 => x"74",
          7464 => x"69",
          7465 => x"6d",
          7466 => x"69",
          7467 => x"6b",
          7468 => x"00",
          7469 => x"44",
          7470 => x"20",
          7471 => x"6f",
          7472 => x"49",
          7473 => x"72",
          7474 => x"20",
          7475 => x"6f",
          7476 => x"00",
          7477 => x"44",
          7478 => x"20",
          7479 => x"20",
          7480 => x"64",
          7481 => x"00",
          7482 => x"4e",
          7483 => x"69",
          7484 => x"66",
          7485 => x"64",
          7486 => x"4e",
          7487 => x"61",
          7488 => x"66",
          7489 => x"64",
          7490 => x"49",
          7491 => x"6c",
          7492 => x"66",
          7493 => x"6e",
          7494 => x"2e",
          7495 => x"41",
          7496 => x"73",
          7497 => x"65",
          7498 => x"64",
          7499 => x"46",
          7500 => x"20",
          7501 => x"65",
          7502 => x"20",
          7503 => x"73",
          7504 => x"0a",
          7505 => x"46",
          7506 => x"20",
          7507 => x"64",
          7508 => x"69",
          7509 => x"6c",
          7510 => x"0a",
          7511 => x"53",
          7512 => x"73",
          7513 => x"69",
          7514 => x"70",
          7515 => x"65",
          7516 => x"64",
          7517 => x"44",
          7518 => x"65",
          7519 => x"6d",
          7520 => x"20",
          7521 => x"69",
          7522 => x"6c",
          7523 => x"0a",
          7524 => x"44",
          7525 => x"20",
          7526 => x"20",
          7527 => x"62",
          7528 => x"2e",
          7529 => x"4e",
          7530 => x"6f",
          7531 => x"74",
          7532 => x"65",
          7533 => x"6c",
          7534 => x"73",
          7535 => x"20",
          7536 => x"6e",
          7537 => x"6e",
          7538 => x"73",
          7539 => x"00",
          7540 => x"46",
          7541 => x"61",
          7542 => x"62",
          7543 => x"65",
          7544 => x"00",
          7545 => x"54",
          7546 => x"6f",
          7547 => x"20",
          7548 => x"72",
          7549 => x"6f",
          7550 => x"61",
          7551 => x"6c",
          7552 => x"2e",
          7553 => x"46",
          7554 => x"20",
          7555 => x"6c",
          7556 => x"65",
          7557 => x"00",
          7558 => x"49",
          7559 => x"66",
          7560 => x"69",
          7561 => x"20",
          7562 => x"6f",
          7563 => x"0a",
          7564 => x"54",
          7565 => x"6d",
          7566 => x"20",
          7567 => x"6e",
          7568 => x"6c",
          7569 => x"0a",
          7570 => x"50",
          7571 => x"6d",
          7572 => x"72",
          7573 => x"6e",
          7574 => x"72",
          7575 => x"2e",
          7576 => x"53",
          7577 => x"65",
          7578 => x"0a",
          7579 => x"55",
          7580 => x"6f",
          7581 => x"65",
          7582 => x"72",
          7583 => x"0a",
          7584 => x"20",
          7585 => x"65",
          7586 => x"73",
          7587 => x"20",
          7588 => x"20",
          7589 => x"65",
          7590 => x"65",
          7591 => x"00",
          7592 => x"72",
          7593 => x"00",
          7594 => x"25",
          7595 => x"00",
          7596 => x"3a",
          7597 => x"25",
          7598 => x"00",
          7599 => x"20",
          7600 => x"20",
          7601 => x"00",
          7602 => x"25",
          7603 => x"00",
          7604 => x"20",
          7605 => x"20",
          7606 => x"7c",
          7607 => x"7a",
          7608 => x"0a",
          7609 => x"25",
          7610 => x"00",
          7611 => x"31",
          7612 => x"34",
          7613 => x"32",
          7614 => x"76",
          7615 => x"31",
          7616 => x"20",
          7617 => x"2c",
          7618 => x"76",
          7619 => x"32",
          7620 => x"25",
          7621 => x"73",
          7622 => x"0a",
          7623 => x"5a",
          7624 => x"49",
          7625 => x"72",
          7626 => x"74",
          7627 => x"6e",
          7628 => x"72",
          7629 => x"54",
          7630 => x"72",
          7631 => x"74",
          7632 => x"75",
          7633 => x"00",
          7634 => x"50",
          7635 => x"69",
          7636 => x"72",
          7637 => x"74",
          7638 => x"49",
          7639 => x"4c",
          7640 => x"20",
          7641 => x"65",
          7642 => x"70",
          7643 => x"49",
          7644 => x"4c",
          7645 => x"20",
          7646 => x"65",
          7647 => x"70",
          7648 => x"55",
          7649 => x"30",
          7650 => x"20",
          7651 => x"65",
          7652 => x"70",
          7653 => x"55",
          7654 => x"30",
          7655 => x"20",
          7656 => x"65",
          7657 => x"70",
          7658 => x"55",
          7659 => x"31",
          7660 => x"20",
          7661 => x"65",
          7662 => x"70",
          7663 => x"55",
          7664 => x"31",
          7665 => x"20",
          7666 => x"65",
          7667 => x"70",
          7668 => x"53",
          7669 => x"69",
          7670 => x"75",
          7671 => x"69",
          7672 => x"2e",
          7673 => x"00",
          7674 => x"45",
          7675 => x"6c",
          7676 => x"20",
          7677 => x"65",
          7678 => x"2e",
          7679 => x"61",
          7680 => x"65",
          7681 => x"2e",
          7682 => x"00",
          7683 => x"30",
          7684 => x"46",
          7685 => x"65",
          7686 => x"6f",
          7687 => x"69",
          7688 => x"6c",
          7689 => x"20",
          7690 => x"63",
          7691 => x"20",
          7692 => x"70",
          7693 => x"73",
          7694 => x"6e",
          7695 => x"6d",
          7696 => x"61",
          7697 => x"2e",
          7698 => x"2a",
          7699 => x"43",
          7700 => x"72",
          7701 => x"2e",
          7702 => x"00",
          7703 => x"43",
          7704 => x"69",
          7705 => x"2e",
          7706 => x"43",
          7707 => x"61",
          7708 => x"67",
          7709 => x"00",
          7710 => x"25",
          7711 => x"78",
          7712 => x"38",
          7713 => x"3e",
          7714 => x"6c",
          7715 => x"30",
          7716 => x"0a",
          7717 => x"44",
          7718 => x"20",
          7719 => x"6f",
          7720 => x"00",
          7721 => x"0a",
          7722 => x"70",
          7723 => x"65",
          7724 => x"25",
          7725 => x"20",
          7726 => x"58",
          7727 => x"3f",
          7728 => x"00",
          7729 => x"25",
          7730 => x"20",
          7731 => x"58",
          7732 => x"25",
          7733 => x"20",
          7734 => x"58",
          7735 => x"45",
          7736 => x"75",
          7737 => x"67",
          7738 => x"64",
          7739 => x"20",
          7740 => x"78",
          7741 => x"2e",
          7742 => x"43",
          7743 => x"69",
          7744 => x"63",
          7745 => x"20",
          7746 => x"30",
          7747 => x"2e",
          7748 => x"00",
          7749 => x"43",
          7750 => x"20",
          7751 => x"75",
          7752 => x"64",
          7753 => x"64",
          7754 => x"25",
          7755 => x"0a",
          7756 => x"52",
          7757 => x"61",
          7758 => x"6e",
          7759 => x"70",
          7760 => x"63",
          7761 => x"6f",
          7762 => x"2e",
          7763 => x"43",
          7764 => x"20",
          7765 => x"6f",
          7766 => x"6e",
          7767 => x"2e",
          7768 => x"5a",
          7769 => x"62",
          7770 => x"25",
          7771 => x"25",
          7772 => x"73",
          7773 => x"00",
          7774 => x"25",
          7775 => x"25",
          7776 => x"73",
          7777 => x"25",
          7778 => x"25",
          7779 => x"42",
          7780 => x"63",
          7781 => x"61",
          7782 => x"0a",
          7783 => x"52",
          7784 => x"69",
          7785 => x"2e",
          7786 => x"45",
          7787 => x"6c",
          7788 => x"20",
          7789 => x"65",
          7790 => x"70",
          7791 => x"2e",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"01",
          7802 => x"01",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"05",
          7808 => x"05",
          7809 => x"05",
          7810 => x"00",
          7811 => x"01",
          7812 => x"01",
          7813 => x"01",
          7814 => x"01",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"01",
          7848 => x"00",
          7849 => x"01",
          7850 => x"00",
          7851 => x"02",
          7852 => x"01",
          7853 => x"00",
          7854 => x"00",
          7855 => x"01",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"01",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"01",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"01",
          7868 => x"00",
          7869 => x"00",
          7870 => x"00",
          7871 => x"01",
          7872 => x"00",
          7873 => x"00",
          7874 => x"00",
          7875 => x"01",
          7876 => x"00",
          7877 => x"00",
          7878 => x"00",
          7879 => x"01",
          7880 => x"00",
          7881 => x"00",
          7882 => x"00",
          7883 => x"01",
          7884 => x"00",
          7885 => x"00",
          7886 => x"00",
          7887 => x"01",
          7888 => x"00",
          7889 => x"00",
          7890 => x"00",
          7891 => x"01",
          7892 => x"00",
          7893 => x"00",
          7894 => x"00",
          7895 => x"01",
          7896 => x"00",
          7897 => x"00",
          7898 => x"00",
          7899 => x"01",
          7900 => x"00",
          7901 => x"00",
          7902 => x"00",
          7903 => x"01",
          7904 => x"00",
          7905 => x"00",
          7906 => x"00",
          7907 => x"01",
          7908 => x"00",
          7909 => x"00",
          7910 => x"00",
          7911 => x"01",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"01",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"01",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"01",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"01",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"01",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"01",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"01",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"01",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"01",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"01",
          7952 => x"00",
          7953 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
