-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b704",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9b040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92fe",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b8299",
          2210 => x"a0738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93830400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80cf",
          2219 => x"942d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80d1",
          2227 => x"802d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"ef040b0b",
          2326 => x"0b8cfe04",
          2327 => x"0b0b0b8d",
          2328 => x"8d040b0b",
          2329 => x"0b8d9c04",
          2330 => x"0b0b0b8d",
          2331 => x"ab040b0b",
          2332 => x"0b8dbb04",
          2333 => x"0b0b0b8d",
          2334 => x"cb040b0b",
          2335 => x"0b8ddb04",
          2336 => x"0b0b0b8d",
          2337 => x"eb040b0b",
          2338 => x"0b8dfb04",
          2339 => x"0b0b0b8e",
          2340 => x"8b040b0b",
          2341 => x"0b8e9b04",
          2342 => x"0b0b0b8e",
          2343 => x"ab040b0b",
          2344 => x"0b8ebb04",
          2345 => x"0b0b0b8e",
          2346 => x"cb040b0b",
          2347 => x"0b8edb04",
          2348 => x"0b0b0b8e",
          2349 => x"eb040b0b",
          2350 => x"0b8efb04",
          2351 => x"0b0b0b8f",
          2352 => x"8b040b0b",
          2353 => x"0b8f9b04",
          2354 => x"0b0b0b8f",
          2355 => x"ab040b0b",
          2356 => x"0b8fbb04",
          2357 => x"0b0b0b8f",
          2358 => x"cb040b0b",
          2359 => x"0b8fdb04",
          2360 => x"0b0b0b8f",
          2361 => x"eb040b0b",
          2362 => x"0b8ffb04",
          2363 => x"0b0b0b90",
          2364 => x"8b040b0b",
          2365 => x"0b909b04",
          2366 => x"0b0b0b90",
          2367 => x"ab040b0b",
          2368 => x"0b90bb04",
          2369 => x"0b0b0b90",
          2370 => x"cb040b0b",
          2371 => x"0b90db04",
          2372 => x"0b0b0b90",
          2373 => x"eb040b0b",
          2374 => x"0b90fb04",
          2375 => x"0b0b0b91",
          2376 => x"8b040b0b",
          2377 => x"0b919b04",
          2378 => x"0b0b0b91",
          2379 => x"ab040b0b",
          2380 => x"0b91bb04",
          2381 => x"0b0b0b91",
          2382 => x"cb040b0b",
          2383 => x"0b91db04",
          2384 => x"0b0b0b91",
          2385 => x"eb040b0b",
          2386 => x"0b91fb04",
          2387 => x"0b0b0b92",
          2388 => x"8b040b0b",
          2389 => x"0b929b04",
          2390 => x"0b0b0b92",
          2391 => x"ab040b0b",
          2392 => x"0b92bb04",
          2393 => x"0b0b0b92",
          2394 => x"cb04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482bba4",
          2434 => x"0c80f8f5",
          2435 => x"2d82bba4",
          2436 => x"0882e090",
          2437 => x"0482bba4",
          2438 => x"0cbed22d",
          2439 => x"82bba408",
          2440 => x"82e09004",
          2441 => x"82bba40c",
          2442 => x"bb832d82",
          2443 => x"bba40882",
          2444 => x"e0900482",
          2445 => x"bba40cb4",
          2446 => x"fc2d82bb",
          2447 => x"a40882e0",
          2448 => x"900482bb",
          2449 => x"a40c94ab",
          2450 => x"2d82bba4",
          2451 => x"0882e090",
          2452 => x"0482bba4",
          2453 => x"0cbce22d",
          2454 => x"82bba408",
          2455 => x"82e09004",
          2456 => x"82bba40c",
          2457 => x"b5b22d82",
          2458 => x"bba40882",
          2459 => x"e0900482",
          2460 => x"bba40caf",
          2461 => x"ab2d82bb",
          2462 => x"a40882e0",
          2463 => x"900482bb",
          2464 => x"a40c93d6",
          2465 => x"2d82bba4",
          2466 => x"0882e090",
          2467 => x"0482bba4",
          2468 => x"0c96be2d",
          2469 => x"82bba408",
          2470 => x"82e09004",
          2471 => x"82bba40c",
          2472 => x"97cb2d82",
          2473 => x"bba40882",
          2474 => x"e0900482",
          2475 => x"bba40c80",
          2476 => x"fc9f2d82",
          2477 => x"bba40882",
          2478 => x"e0900482",
          2479 => x"bba40c80",
          2480 => x"fcfd2d82",
          2481 => x"bba40882",
          2482 => x"e0900482",
          2483 => x"bba40c80",
          2484 => x"f4b92d82",
          2485 => x"bba40882",
          2486 => x"e0900482",
          2487 => x"bba40c80",
          2488 => x"f6b12d82",
          2489 => x"bba40882",
          2490 => x"e0900482",
          2491 => x"bba40c80",
          2492 => x"f7e42d82",
          2493 => x"bba40882",
          2494 => x"e0900482",
          2495 => x"bba40c81",
          2496 => x"dc842d82",
          2497 => x"bba40882",
          2498 => x"e0900482",
          2499 => x"bba40c81",
          2500 => x"e8f52d82",
          2501 => x"bba40882",
          2502 => x"e0900482",
          2503 => x"bba40c81",
          2504 => x"e0e92d82",
          2505 => x"bba40882",
          2506 => x"e0900482",
          2507 => x"bba40c81",
          2508 => x"e3e62d82",
          2509 => x"bba40882",
          2510 => x"e0900482",
          2511 => x"bba40c81",
          2512 => x"ee842d82",
          2513 => x"bba40882",
          2514 => x"e0900482",
          2515 => x"bba40c81",
          2516 => x"f6e42d82",
          2517 => x"bba40882",
          2518 => x"e0900482",
          2519 => x"bba40c81",
          2520 => x"e7d72d82",
          2521 => x"bba40882",
          2522 => x"e0900482",
          2523 => x"bba40c81",
          2524 => x"f1a32d82",
          2525 => x"bba40882",
          2526 => x"e0900482",
          2527 => x"bba40c81",
          2528 => x"f2c22d82",
          2529 => x"bba40882",
          2530 => x"e0900482",
          2531 => x"bba40c81",
          2532 => x"f2e12d82",
          2533 => x"bba40882",
          2534 => x"e0900482",
          2535 => x"bba40c81",
          2536 => x"facb2d82",
          2537 => x"bba40882",
          2538 => x"e0900482",
          2539 => x"bba40c81",
          2540 => x"f8b12d82",
          2541 => x"bba40882",
          2542 => x"e0900482",
          2543 => x"bba40c81",
          2544 => x"fd9f2d82",
          2545 => x"bba40882",
          2546 => x"e0900482",
          2547 => x"bba40c81",
          2548 => x"f3e52d82",
          2549 => x"bba40882",
          2550 => x"e0900482",
          2551 => x"bba40c82",
          2552 => x"809f2d82",
          2553 => x"bba40882",
          2554 => x"e0900482",
          2555 => x"bba40c82",
          2556 => x"81a02d82",
          2557 => x"bba40882",
          2558 => x"e0900482",
          2559 => x"bba40c81",
          2560 => x"e9d52d82",
          2561 => x"bba40882",
          2562 => x"e0900482",
          2563 => x"bba40c81",
          2564 => x"e9ae2d82",
          2565 => x"bba40882",
          2566 => x"e0900482",
          2567 => x"bba40c81",
          2568 => x"ead92d82",
          2569 => x"bba40882",
          2570 => x"e0900482",
          2571 => x"bba40c81",
          2572 => x"f4bc2d82",
          2573 => x"bba40882",
          2574 => x"e0900482",
          2575 => x"bba40c82",
          2576 => x"82912d82",
          2577 => x"bba40882",
          2578 => x"e0900482",
          2579 => x"bba40c82",
          2580 => x"849b2d82",
          2581 => x"bba40882",
          2582 => x"e0900482",
          2583 => x"bba40c82",
          2584 => x"87dd2d82",
          2585 => x"bba40882",
          2586 => x"e0900482",
          2587 => x"bba40c81",
          2588 => x"dba32d82",
          2589 => x"bba40882",
          2590 => x"e0900482",
          2591 => x"bba40c82",
          2592 => x"8ac92d82",
          2593 => x"bba40882",
          2594 => x"e0900482",
          2595 => x"bba40c82",
          2596 => x"98fe2d82",
          2597 => x"bba40882",
          2598 => x"e0900482",
          2599 => x"bba40c82",
          2600 => x"96ea2d82",
          2601 => x"bba40882",
          2602 => x"e0900482",
          2603 => x"bba40c81",
          2604 => x"acde2d82",
          2605 => x"bba40882",
          2606 => x"e0900482",
          2607 => x"bba40c81",
          2608 => x"aec82d82",
          2609 => x"bba40882",
          2610 => x"e0900482",
          2611 => x"bba40c81",
          2612 => x"b0ac2d82",
          2613 => x"bba40882",
          2614 => x"e0900482",
          2615 => x"bba40c80",
          2616 => x"f4e22d82",
          2617 => x"bba40882",
          2618 => x"e0900482",
          2619 => x"bba40c80",
          2620 => x"f6862d82",
          2621 => x"bba40882",
          2622 => x"e0900482",
          2623 => x"bba40c80",
          2624 => x"f9ea2d82",
          2625 => x"bba40882",
          2626 => x"e0900482",
          2627 => x"bba40c80",
          2628 => x"d6962d82",
          2629 => x"bba40882",
          2630 => x"e0900482",
          2631 => x"bba40c81",
          2632 => x"a6f22d82",
          2633 => x"bba40882",
          2634 => x"e0900482",
          2635 => x"bba40c81",
          2636 => x"a79a2d82",
          2637 => x"bba40882",
          2638 => x"e0900482",
          2639 => x"bba40c81",
          2640 => x"ab922d82",
          2641 => x"bba40882",
          2642 => x"e0900482",
          2643 => x"bba40c81",
          2644 => x"a3dc2d82",
          2645 => x"bba40882",
          2646 => x"e090043c",
          2647 => x"04000010",
          2648 => x"10101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10105351",
          2656 => x"04000073",
          2657 => x"81ff0673",
          2658 => x"83060981",
          2659 => x"05830510",
          2660 => x"10102b07",
          2661 => x"72fc060c",
          2662 => x"51510472",
          2663 => x"72807281",
          2664 => x"06ff0509",
          2665 => x"72060571",
          2666 => x"1052720a",
          2667 => x"100a5372",
          2668 => x"ed385151",
          2669 => x"53510482",
          2670 => x"bb987082",
          2671 => x"d2f4278e",
          2672 => x"38807170",
          2673 => x"8405530c",
          2674 => x"0b0b0b93",
          2675 => x"ba048c81",
          2676 => x"5180f2fe",
          2677 => x"040082bb",
          2678 => x"a4080282",
          2679 => x"bba40cfb",
          2680 => x"3d0d82bb",
          2681 => x"a4088c05",
          2682 => x"7082bba4",
          2683 => x"08fc050c",
          2684 => x"82bba408",
          2685 => x"fc050854",
          2686 => x"82bba408",
          2687 => x"88050853",
          2688 => x"82d2ec08",
          2689 => x"5254849a",
          2690 => x"3f82bb98",
          2691 => x"087082bb",
          2692 => x"a408f805",
          2693 => x"0c82bba4",
          2694 => x"08f80508",
          2695 => x"7082bb98",
          2696 => x"0c515487",
          2697 => x"3d0d82bb",
          2698 => x"a40c0482",
          2699 => x"bba40802",
          2700 => x"82bba40c",
          2701 => x"fb3d0d82",
          2702 => x"bba40890",
          2703 => x"05088511",
          2704 => x"33708132",
          2705 => x"70810651",
          2706 => x"51515271",
          2707 => x"8f38800b",
          2708 => x"82bba408",
          2709 => x"8c050825",
          2710 => x"83388d39",
          2711 => x"800b82bb",
          2712 => x"a408f405",
          2713 => x"0c81c439",
          2714 => x"82bba408",
          2715 => x"8c0508ff",
          2716 => x"0582bba4",
          2717 => x"088c050c",
          2718 => x"800b82bb",
          2719 => x"a408f805",
          2720 => x"0c82bba4",
          2721 => x"08880508",
          2722 => x"82bba408",
          2723 => x"fc050c82",
          2724 => x"bba408f8",
          2725 => x"05088a2e",
          2726 => x"80f63880",
          2727 => x"0b82bba4",
          2728 => x"088c0508",
          2729 => x"2580e938",
          2730 => x"82bba408",
          2731 => x"90050851",
          2732 => x"abb23f82",
          2733 => x"bb980870",
          2734 => x"82bba408",
          2735 => x"f8050c52",
          2736 => x"82bba408",
          2737 => x"f80508ff",
          2738 => x"2e098106",
          2739 => x"8d38800b",
          2740 => x"82bba408",
          2741 => x"f4050c80",
          2742 => x"d23982bb",
          2743 => x"a408fc05",
          2744 => x"0882bba4",
          2745 => x"08f80508",
          2746 => x"53537173",
          2747 => x"3482bba4",
          2748 => x"088c0508",
          2749 => x"ff0582bb",
          2750 => x"a4088c05",
          2751 => x"0c82bba4",
          2752 => x"08fc0508",
          2753 => x"810582bb",
          2754 => x"a408fc05",
          2755 => x"0cff8039",
          2756 => x"82bba408",
          2757 => x"fc050852",
          2758 => x"80723482",
          2759 => x"bba40888",
          2760 => x"05087082",
          2761 => x"bba408f4",
          2762 => x"050c5282",
          2763 => x"bba408f4",
          2764 => x"050882bb",
          2765 => x"980c873d",
          2766 => x"0d82bba4",
          2767 => x"0c0482bb",
          2768 => x"a4080282",
          2769 => x"bba40cf4",
          2770 => x"3d0d860b",
          2771 => x"82bba408",
          2772 => x"e5053482",
          2773 => x"bba40888",
          2774 => x"050882bb",
          2775 => x"a408e005",
          2776 => x"0cfe0a0b",
          2777 => x"82bba408",
          2778 => x"e8050c82",
          2779 => x"bba40890",
          2780 => x"057082bb",
          2781 => x"a408fc05",
          2782 => x"0c82bba4",
          2783 => x"08fc0508",
          2784 => x"5482bba4",
          2785 => x"088c0508",
          2786 => x"5382bba4",
          2787 => x"08e00570",
          2788 => x"53515481",
          2789 => x"8d3f82bb",
          2790 => x"98087082",
          2791 => x"bba408dc",
          2792 => x"050c82bb",
          2793 => x"a408ec05",
          2794 => x"0882bba4",
          2795 => x"08880508",
          2796 => x"05515480",
          2797 => x"743482bb",
          2798 => x"a408dc05",
          2799 => x"087082bb",
          2800 => x"980c548e",
          2801 => x"3d0d82bb",
          2802 => x"a40c0482",
          2803 => x"bba40802",
          2804 => x"82bba40c",
          2805 => x"fb3d0d82",
          2806 => x"bba40890",
          2807 => x"057082bb",
          2808 => x"a408fc05",
          2809 => x"0c82bba4",
          2810 => x"08fc0508",
          2811 => x"5482bba4",
          2812 => x"088c0508",
          2813 => x"5382bba4",
          2814 => x"08880508",
          2815 => x"5254a33f",
          2816 => x"82bb9808",
          2817 => x"7082bba4",
          2818 => x"08f8050c",
          2819 => x"82bba408",
          2820 => x"f8050870",
          2821 => x"82bb980c",
          2822 => x"5154873d",
          2823 => x"0d82bba4",
          2824 => x"0c0482bb",
          2825 => x"a4080282",
          2826 => x"bba40ced",
          2827 => x"3d0d800b",
          2828 => x"82bba408",
          2829 => x"e4052382",
          2830 => x"bba40888",
          2831 => x"05085380",
          2832 => x"0b8c140c",
          2833 => x"82bba408",
          2834 => x"88050885",
          2835 => x"11337081",
          2836 => x"2a708132",
          2837 => x"70810651",
          2838 => x"51515153",
          2839 => x"72802e8d",
          2840 => x"38ff0b82",
          2841 => x"bba408e0",
          2842 => x"050c96ac",
          2843 => x"3982bba4",
          2844 => x"088c0508",
          2845 => x"53723353",
          2846 => x"7282bba4",
          2847 => x"08f80534",
          2848 => x"7281ff06",
          2849 => x"5372802e",
          2850 => x"95fa3882",
          2851 => x"bba4088c",
          2852 => x"05088105",
          2853 => x"82bba408",
          2854 => x"8c050c82",
          2855 => x"bba408e4",
          2856 => x"05227081",
          2857 => x"06515372",
          2858 => x"802e958b",
          2859 => x"3882bba4",
          2860 => x"08f80533",
          2861 => x"53af7327",
          2862 => x"81fc3882",
          2863 => x"bba408f8",
          2864 => x"05335372",
          2865 => x"b92681ee",
          2866 => x"3882bba4",
          2867 => x"08f80533",
          2868 => x"5372b02e",
          2869 => x"09810680",
          2870 => x"c53882bb",
          2871 => x"a408e805",
          2872 => x"3370982b",
          2873 => x"70982c51",
          2874 => x"515372b2",
          2875 => x"3882bba4",
          2876 => x"08e40522",
          2877 => x"70832a70",
          2878 => x"81327081",
          2879 => x"06515151",
          2880 => x"5372802e",
          2881 => x"993882bb",
          2882 => x"a408e405",
          2883 => x"22708280",
          2884 => x"07515372",
          2885 => x"82bba408",
          2886 => x"e40523fe",
          2887 => x"d03982bb",
          2888 => x"a408e805",
          2889 => x"3370982b",
          2890 => x"70982c70",
          2891 => x"70832b72",
          2892 => x"11731151",
          2893 => x"51515351",
          2894 => x"55537282",
          2895 => x"bba408e8",
          2896 => x"053482bb",
          2897 => x"a408e805",
          2898 => x"335482bb",
          2899 => x"a408f805",
          2900 => x"337015d0",
          2901 => x"11515153",
          2902 => x"7282bba4",
          2903 => x"08e80534",
          2904 => x"82bba408",
          2905 => x"e8053370",
          2906 => x"982b7098",
          2907 => x"2c515153",
          2908 => x"7280258b",
          2909 => x"3880ff0b",
          2910 => x"82bba408",
          2911 => x"e8053482",
          2912 => x"bba408e4",
          2913 => x"05227083",
          2914 => x"2a708106",
          2915 => x"51515372",
          2916 => x"fddb3882",
          2917 => x"bba408e8",
          2918 => x"05337088",
          2919 => x"2b70902b",
          2920 => x"70902c70",
          2921 => x"882c5151",
          2922 => x"51515372",
          2923 => x"82bba408",
          2924 => x"ec0523fd",
          2925 => x"b83982bb",
          2926 => x"a408e405",
          2927 => x"2270832a",
          2928 => x"70810651",
          2929 => x"51537280",
          2930 => x"2e9d3882",
          2931 => x"bba408e8",
          2932 => x"05337098",
          2933 => x"2b70982c",
          2934 => x"51515372",
          2935 => x"8a38810b",
          2936 => x"82bba408",
          2937 => x"e8053482",
          2938 => x"bba408f8",
          2939 => x"0533e011",
          2940 => x"82bba408",
          2941 => x"c4050c53",
          2942 => x"82bba408",
          2943 => x"c4050880",
          2944 => x"d8269294",
          2945 => x"3882bba4",
          2946 => x"08c40508",
          2947 => x"70822b82",
          2948 => x"9aec1170",
          2949 => x"08515151",
          2950 => x"53720482",
          2951 => x"bba408e4",
          2952 => x"05227090",
          2953 => x"07515372",
          2954 => x"82bba408",
          2955 => x"e4052382",
          2956 => x"bba408e4",
          2957 => x"052270a0",
          2958 => x"07515372",
          2959 => x"82bba408",
          2960 => x"e40523fc",
          2961 => x"a83982bb",
          2962 => x"a408e405",
          2963 => x"22708180",
          2964 => x"07515372",
          2965 => x"82bba408",
          2966 => x"e40523fc",
          2967 => x"903982bb",
          2968 => x"a408e405",
          2969 => x"227080c0",
          2970 => x"07515372",
          2971 => x"82bba408",
          2972 => x"e40523fb",
          2973 => x"f83982bb",
          2974 => x"a408e405",
          2975 => x"22708807",
          2976 => x"51537282",
          2977 => x"bba408e4",
          2978 => x"0523800b",
          2979 => x"82bba408",
          2980 => x"e80534fb",
          2981 => x"d83982bb",
          2982 => x"a408e405",
          2983 => x"22708407",
          2984 => x"51537282",
          2985 => x"bba408e4",
          2986 => x"0523fbc1",
          2987 => x"39bf0b82",
          2988 => x"bba408fc",
          2989 => x"053482bb",
          2990 => x"a408ec05",
          2991 => x"22ff1151",
          2992 => x"537282bb",
          2993 => x"a408ec05",
          2994 => x"2380e30b",
          2995 => x"82bba408",
          2996 => x"f805348d",
          2997 => x"a83982bb",
          2998 => x"a4089005",
          2999 => x"0882bba4",
          3000 => x"08900508",
          3001 => x"840582bb",
          3002 => x"a4089005",
          3003 => x"0c700851",
          3004 => x"537282bb",
          3005 => x"a408fc05",
          3006 => x"3482bba4",
          3007 => x"08ec0522",
          3008 => x"ff115153",
          3009 => x"7282bba4",
          3010 => x"08ec0523",
          3011 => x"8cef3982",
          3012 => x"bba40890",
          3013 => x"050882bb",
          3014 => x"a4089005",
          3015 => x"08840582",
          3016 => x"bba40890",
          3017 => x"050c7008",
          3018 => x"82bba408",
          3019 => x"fc050c82",
          3020 => x"bba408e4",
          3021 => x"05227083",
          3022 => x"2a708106",
          3023 => x"51515153",
          3024 => x"72802eab",
          3025 => x"3882bba4",
          3026 => x"08e80533",
          3027 => x"70982b53",
          3028 => x"72982c53",
          3029 => x"82bba408",
          3030 => x"fc050852",
          3031 => x"53adfa3f",
          3032 => x"82bb9808",
          3033 => x"537282bb",
          3034 => x"a408f405",
          3035 => x"23993982",
          3036 => x"bba408fc",
          3037 => x"050851a8",
          3038 => x"ac3f82bb",
          3039 => x"98085372",
          3040 => x"82bba408",
          3041 => x"f4052382",
          3042 => x"bba408ec",
          3043 => x"05225382",
          3044 => x"bba408f4",
          3045 => x"05227371",
          3046 => x"31545472",
          3047 => x"82bba408",
          3048 => x"ec05238b",
          3049 => x"d83982bb",
          3050 => x"a4089005",
          3051 => x"0882bba4",
          3052 => x"08900508",
          3053 => x"840582bb",
          3054 => x"a4089005",
          3055 => x"0c700882",
          3056 => x"bba408fc",
          3057 => x"050c82bb",
          3058 => x"a408e405",
          3059 => x"2270832a",
          3060 => x"70810651",
          3061 => x"51515372",
          3062 => x"802eab38",
          3063 => x"82bba408",
          3064 => x"e8053370",
          3065 => x"982b5372",
          3066 => x"982c5382",
          3067 => x"bba408fc",
          3068 => x"05085253",
          3069 => x"ace33f82",
          3070 => x"bb980853",
          3071 => x"7282bba4",
          3072 => x"08f40523",
          3073 => x"993982bb",
          3074 => x"a408fc05",
          3075 => x"0851a795",
          3076 => x"3f82bb98",
          3077 => x"08537282",
          3078 => x"bba408f4",
          3079 => x"052382bb",
          3080 => x"a408ec05",
          3081 => x"225382bb",
          3082 => x"a408f405",
          3083 => x"22737131",
          3084 => x"54547282",
          3085 => x"bba408ec",
          3086 => x"05238ac1",
          3087 => x"3982bba4",
          3088 => x"08e40522",
          3089 => x"70822a70",
          3090 => x"81065151",
          3091 => x"5372802e",
          3092 => x"a43882bb",
          3093 => x"a4089005",
          3094 => x"0882bba4",
          3095 => x"08900508",
          3096 => x"840582bb",
          3097 => x"a4089005",
          3098 => x"0c700882",
          3099 => x"bba408dc",
          3100 => x"050c53a2",
          3101 => x"3982bba4",
          3102 => x"08900508",
          3103 => x"82bba408",
          3104 => x"90050884",
          3105 => x"0582bba4",
          3106 => x"0890050c",
          3107 => x"700882bb",
          3108 => x"a408dc05",
          3109 => x"0c5382bb",
          3110 => x"a408dc05",
          3111 => x"0882bba4",
          3112 => x"08fc050c",
          3113 => x"82bba408",
          3114 => x"fc050880",
          3115 => x"25a43882",
          3116 => x"bba408e4",
          3117 => x"05227082",
          3118 => x"07515372",
          3119 => x"82bba408",
          3120 => x"e4052382",
          3121 => x"bba408fc",
          3122 => x"05083082",
          3123 => x"bba408fc",
          3124 => x"050c82bb",
          3125 => x"a408e405",
          3126 => x"2270ffbf",
          3127 => x"06515372",
          3128 => x"82bba408",
          3129 => x"e4052381",
          3130 => x"af39880b",
          3131 => x"82bba408",
          3132 => x"f40523a9",
          3133 => x"3982bba4",
          3134 => x"08e40522",
          3135 => x"7080c007",
          3136 => x"51537282",
          3137 => x"bba408e4",
          3138 => x"052380f8",
          3139 => x"0b82bba4",
          3140 => x"08f80534",
          3141 => x"900b82bb",
          3142 => x"a408f405",
          3143 => x"2382bba4",
          3144 => x"08e40522",
          3145 => x"70822a70",
          3146 => x"81065151",
          3147 => x"5372802e",
          3148 => x"a43882bb",
          3149 => x"a4089005",
          3150 => x"0882bba4",
          3151 => x"08900508",
          3152 => x"840582bb",
          3153 => x"a4089005",
          3154 => x"0c700882",
          3155 => x"bba408d8",
          3156 => x"050c53a2",
          3157 => x"3982bba4",
          3158 => x"08900508",
          3159 => x"82bba408",
          3160 => x"90050884",
          3161 => x"0582bba4",
          3162 => x"0890050c",
          3163 => x"700882bb",
          3164 => x"a408d805",
          3165 => x"0c5382bb",
          3166 => x"a408d805",
          3167 => x"0882bba4",
          3168 => x"08fc050c",
          3169 => x"82bba408",
          3170 => x"e4052270",
          3171 => x"cf065153",
          3172 => x"7282bba4",
          3173 => x"08e40523",
          3174 => x"82bba80b",
          3175 => x"82bba408",
          3176 => x"f0050c82",
          3177 => x"bba408f0",
          3178 => x"050882bb",
          3179 => x"a408f405",
          3180 => x"2282bba4",
          3181 => x"08fc0508",
          3182 => x"71557054",
          3183 => x"565455af",
          3184 => x"953f82bb",
          3185 => x"98085372",
          3186 => x"753482bb",
          3187 => x"a408f005",
          3188 => x"0882bba4",
          3189 => x"08d4050c",
          3190 => x"82bba408",
          3191 => x"f0050870",
          3192 => x"33515389",
          3193 => x"7327a438",
          3194 => x"82bba408",
          3195 => x"f0050853",
          3196 => x"72335482",
          3197 => x"bba408f8",
          3198 => x"05337015",
          3199 => x"df115151",
          3200 => x"537282bb",
          3201 => x"a408d005",
          3202 => x"34973982",
          3203 => x"bba408f0",
          3204 => x"05085372",
          3205 => x"33b01151",
          3206 => x"537282bb",
          3207 => x"a408d005",
          3208 => x"3482bba4",
          3209 => x"08d40508",
          3210 => x"5382bba4",
          3211 => x"08d00533",
          3212 => x"733482bb",
          3213 => x"a408f005",
          3214 => x"08810582",
          3215 => x"bba408f0",
          3216 => x"050c82bb",
          3217 => x"a408f405",
          3218 => x"22705382",
          3219 => x"bba408fc",
          3220 => x"05085253",
          3221 => x"adcd3f82",
          3222 => x"bb980870",
          3223 => x"82bba408",
          3224 => x"fc050c53",
          3225 => x"82bba408",
          3226 => x"fc050880",
          3227 => x"2e8438fe",
          3228 => x"b23982bb",
          3229 => x"a408f005",
          3230 => x"0882bba8",
          3231 => x"54557254",
          3232 => x"74707531",
          3233 => x"51537282",
          3234 => x"bba408fc",
          3235 => x"053482bb",
          3236 => x"a408e405",
          3237 => x"2270b206",
          3238 => x"51537280",
          3239 => x"2e943882",
          3240 => x"bba408ec",
          3241 => x"0522ff11",
          3242 => x"51537282",
          3243 => x"bba408ec",
          3244 => x"052382bb",
          3245 => x"a408e405",
          3246 => x"2270862a",
          3247 => x"70810651",
          3248 => x"51537280",
          3249 => x"2e80e738",
          3250 => x"82bba408",
          3251 => x"ec052270",
          3252 => x"902b82bb",
          3253 => x"a408cc05",
          3254 => x"0c82bba4",
          3255 => x"08cc0508",
          3256 => x"902c82bb",
          3257 => x"a408cc05",
          3258 => x"0c82bba4",
          3259 => x"08f40522",
          3260 => x"51537290",
          3261 => x"2e098106",
          3262 => x"953882bb",
          3263 => x"a408cc05",
          3264 => x"08fe0553",
          3265 => x"7282bba4",
          3266 => x"08c80523",
          3267 => x"933982bb",
          3268 => x"a408cc05",
          3269 => x"08ff0553",
          3270 => x"7282bba4",
          3271 => x"08c80523",
          3272 => x"82bba408",
          3273 => x"c8052282",
          3274 => x"bba408ec",
          3275 => x"052382bb",
          3276 => x"a408e405",
          3277 => x"2270832a",
          3278 => x"70810651",
          3279 => x"51537280",
          3280 => x"2e80d038",
          3281 => x"82bba408",
          3282 => x"e8053370",
          3283 => x"982b7098",
          3284 => x"2c82bba4",
          3285 => x"08fc0533",
          3286 => x"57515153",
          3287 => x"72742497",
          3288 => x"3882bba4",
          3289 => x"08e40522",
          3290 => x"70f70651",
          3291 => x"537282bb",
          3292 => x"a408e405",
          3293 => x"239d3982",
          3294 => x"bba408e8",
          3295 => x"05335382",
          3296 => x"bba408fc",
          3297 => x"05337371",
          3298 => x"31545472",
          3299 => x"82bba408",
          3300 => x"e8053482",
          3301 => x"bba408e4",
          3302 => x"05227083",
          3303 => x"2a708106",
          3304 => x"51515372",
          3305 => x"802eb138",
          3306 => x"82bba408",
          3307 => x"e8053370",
          3308 => x"882b7090",
          3309 => x"2b70902c",
          3310 => x"70882c51",
          3311 => x"51515153",
          3312 => x"725482bb",
          3313 => x"a408ec05",
          3314 => x"22707531",
          3315 => x"51537282",
          3316 => x"bba408ec",
          3317 => x"0523af39",
          3318 => x"82bba408",
          3319 => x"fc053370",
          3320 => x"882b7090",
          3321 => x"2b70902c",
          3322 => x"70882c51",
          3323 => x"51515153",
          3324 => x"725482bb",
          3325 => x"a408ec05",
          3326 => x"22707531",
          3327 => x"51537282",
          3328 => x"bba408ec",
          3329 => x"052382bb",
          3330 => x"a408e405",
          3331 => x"22708380",
          3332 => x"06515372",
          3333 => x"b03882bb",
          3334 => x"a408ec05",
          3335 => x"22ff1154",
          3336 => x"547282bb",
          3337 => x"a408ec05",
          3338 => x"2373902b",
          3339 => x"70902c51",
          3340 => x"53807325",
          3341 => x"903882bb",
          3342 => x"a4088805",
          3343 => x"0852a051",
          3344 => x"96903fd2",
          3345 => x"3982bba4",
          3346 => x"08e40522",
          3347 => x"70812a70",
          3348 => x"81065151",
          3349 => x"5372802e",
          3350 => x"913882bb",
          3351 => x"a4088805",
          3352 => x"0852ad51",
          3353 => x"95ec3f80",
          3354 => x"c73982bb",
          3355 => x"a408e405",
          3356 => x"2270842a",
          3357 => x"70810651",
          3358 => x"51537280",
          3359 => x"2e903882",
          3360 => x"bba40888",
          3361 => x"050852ab",
          3362 => x"5195c73f",
          3363 => x"a33982bb",
          3364 => x"a408e405",
          3365 => x"2270852a",
          3366 => x"70810651",
          3367 => x"51537280",
          3368 => x"2e8e3882",
          3369 => x"bba40888",
          3370 => x"050852a0",
          3371 => x"5195a33f",
          3372 => x"82bba408",
          3373 => x"e4052270",
          3374 => x"862a7081",
          3375 => x"06515153",
          3376 => x"72802eb1",
          3377 => x"3882bba4",
          3378 => x"08880508",
          3379 => x"52b05195",
          3380 => x"813f82bb",
          3381 => x"a408f405",
          3382 => x"22537290",
          3383 => x"2e098106",
          3384 => x"943882bb",
          3385 => x"a4088805",
          3386 => x"085282bb",
          3387 => x"a408f805",
          3388 => x"335194de",
          3389 => x"3f82bba4",
          3390 => x"08e40522",
          3391 => x"70882a70",
          3392 => x"81065151",
          3393 => x"5372802e",
          3394 => x"b03882bb",
          3395 => x"a408ec05",
          3396 => x"22ff1154",
          3397 => x"547282bb",
          3398 => x"a408ec05",
          3399 => x"2373902b",
          3400 => x"70902c51",
          3401 => x"53807325",
          3402 => x"903882bb",
          3403 => x"a4088805",
          3404 => x"0852b051",
          3405 => x"949c3fd2",
          3406 => x"3982bba4",
          3407 => x"08e40522",
          3408 => x"70832a70",
          3409 => x"81065151",
          3410 => x"5372802e",
          3411 => x"b03882bb",
          3412 => x"a408e805",
          3413 => x"33ff1154",
          3414 => x"547282bb",
          3415 => x"a408e805",
          3416 => x"3473982b",
          3417 => x"70982c51",
          3418 => x"53807325",
          3419 => x"903882bb",
          3420 => x"a4088805",
          3421 => x"0852b051",
          3422 => x"93d83fd2",
          3423 => x"3982bba4",
          3424 => x"08e40522",
          3425 => x"70872a70",
          3426 => x"81065151",
          3427 => x"5372b038",
          3428 => x"82bba408",
          3429 => x"ec0522ff",
          3430 => x"11545472",
          3431 => x"82bba408",
          3432 => x"ec052373",
          3433 => x"902b7090",
          3434 => x"2c515380",
          3435 => x"73259038",
          3436 => x"82bba408",
          3437 => x"88050852",
          3438 => x"a0519396",
          3439 => x"3fd23982",
          3440 => x"bba408f8",
          3441 => x"05335372",
          3442 => x"80e32e09",
          3443 => x"81069738",
          3444 => x"82bba408",
          3445 => x"88050852",
          3446 => x"82bba408",
          3447 => x"fc053351",
          3448 => x"92f03f81",
          3449 => x"ee3982bb",
          3450 => x"a408f805",
          3451 => x"33537280",
          3452 => x"f32e0981",
          3453 => x"0680cb38",
          3454 => x"82bba408",
          3455 => x"f40522ff",
          3456 => x"11515372",
          3457 => x"82bba408",
          3458 => x"f4052372",
          3459 => x"83ffff06",
          3460 => x"537283ff",
          3461 => x"ff2e81bb",
          3462 => x"3882bba4",
          3463 => x"08880508",
          3464 => x"5282bba4",
          3465 => x"08fc0508",
          3466 => x"70335282",
          3467 => x"bba408fc",
          3468 => x"05088105",
          3469 => x"82bba408",
          3470 => x"fc050c53",
          3471 => x"92943fff",
          3472 => x"b73982bb",
          3473 => x"a408f805",
          3474 => x"33537280",
          3475 => x"d32e0981",
          3476 => x"0680cb38",
          3477 => x"82bba408",
          3478 => x"f40522ff",
          3479 => x"11515372",
          3480 => x"82bba408",
          3481 => x"f4052372",
          3482 => x"83ffff06",
          3483 => x"537283ff",
          3484 => x"ff2e80df",
          3485 => x"3882bba4",
          3486 => x"08880508",
          3487 => x"5282bba4",
          3488 => x"08fc0508",
          3489 => x"70335253",
          3490 => x"91c83f82",
          3491 => x"bba408fc",
          3492 => x"05088105",
          3493 => x"82bba408",
          3494 => x"fc050cff",
          3495 => x"b73982bb",
          3496 => x"a408f005",
          3497 => x"0882bba8",
          3498 => x"2ea93882",
          3499 => x"bba40888",
          3500 => x"05085282",
          3501 => x"bba408f0",
          3502 => x"0508ff05",
          3503 => x"82bba408",
          3504 => x"f0050c82",
          3505 => x"bba408f0",
          3506 => x"05087033",
          3507 => x"52539182",
          3508 => x"3fcc3982",
          3509 => x"bba408e4",
          3510 => x"05227087",
          3511 => x"2a708106",
          3512 => x"51515372",
          3513 => x"802e80c3",
          3514 => x"3882bba4",
          3515 => x"08ec0522",
          3516 => x"ff115454",
          3517 => x"7282bba4",
          3518 => x"08ec0523",
          3519 => x"73902b70",
          3520 => x"902c5153",
          3521 => x"807325a3",
          3522 => x"3882bba4",
          3523 => x"08880508",
          3524 => x"52a05190",
          3525 => x"bd3fd239",
          3526 => x"82bba408",
          3527 => x"88050852",
          3528 => x"82bba408",
          3529 => x"f8053351",
          3530 => x"90a83f80",
          3531 => x"0b82bba4",
          3532 => x"08e40523",
          3533 => x"eab73982",
          3534 => x"bba408f8",
          3535 => x"05335372",
          3536 => x"a52e0981",
          3537 => x"06a83881",
          3538 => x"0b82bba4",
          3539 => x"08e40523",
          3540 => x"800b82bb",
          3541 => x"a408ec05",
          3542 => x"23800b82",
          3543 => x"bba408e8",
          3544 => x"05348a0b",
          3545 => x"82bba408",
          3546 => x"f40523ea",
          3547 => x"803982bb",
          3548 => x"a4088805",
          3549 => x"085282bb",
          3550 => x"a408f805",
          3551 => x"33518fd2",
          3552 => x"3fe9ea39",
          3553 => x"82bba408",
          3554 => x"8805088c",
          3555 => x"11087082",
          3556 => x"bba408e0",
          3557 => x"050c5153",
          3558 => x"82bba408",
          3559 => x"e0050882",
          3560 => x"bb980c95",
          3561 => x"3d0d82bb",
          3562 => x"a40c0482",
          3563 => x"bba40802",
          3564 => x"82bba40c",
          3565 => x"f73d0d80",
          3566 => x"0b82bba4",
          3567 => x"08f00534",
          3568 => x"82bba408",
          3569 => x"8c050853",
          3570 => x"80730c82",
          3571 => x"bba40888",
          3572 => x"05087008",
          3573 => x"51537233",
          3574 => x"537282bb",
          3575 => x"a408f805",
          3576 => x"347281ff",
          3577 => x"065372a0",
          3578 => x"2e098106",
          3579 => x"913882bb",
          3580 => x"a4088805",
          3581 => x"08700881",
          3582 => x"05710c53",
          3583 => x"ce3982bb",
          3584 => x"a408f805",
          3585 => x"335372ad",
          3586 => x"2e098106",
          3587 => x"a438810b",
          3588 => x"82bba408",
          3589 => x"f0053482",
          3590 => x"bba40888",
          3591 => x"05087008",
          3592 => x"8105710c",
          3593 => x"70085153",
          3594 => x"723382bb",
          3595 => x"a408f805",
          3596 => x"3482bba4",
          3597 => x"08f80533",
          3598 => x"5372b02e",
          3599 => x"09810681",
          3600 => x"dc3882bb",
          3601 => x"a4088805",
          3602 => x"08700881",
          3603 => x"05710c70",
          3604 => x"08515372",
          3605 => x"3382bba4",
          3606 => x"08f80534",
          3607 => x"82bba408",
          3608 => x"f8053382",
          3609 => x"bba408e8",
          3610 => x"050c82bb",
          3611 => x"a408e805",
          3612 => x"0880e22e",
          3613 => x"b63882bb",
          3614 => x"a408e805",
          3615 => x"0880f82e",
          3616 => x"843880cd",
          3617 => x"39900b82",
          3618 => x"bba408f4",
          3619 => x"053482bb",
          3620 => x"a4088805",
          3621 => x"08700881",
          3622 => x"05710c70",
          3623 => x"08515372",
          3624 => x"3382bba4",
          3625 => x"08f80534",
          3626 => x"81a43982",
          3627 => x"0b82bba4",
          3628 => x"08f40534",
          3629 => x"82bba408",
          3630 => x"88050870",
          3631 => x"08810571",
          3632 => x"0c700851",
          3633 => x"53723382",
          3634 => x"bba408f8",
          3635 => x"053480fe",
          3636 => x"3982bba4",
          3637 => x"08f80533",
          3638 => x"5372a026",
          3639 => x"8d38810b",
          3640 => x"82bba408",
          3641 => x"ec050c83",
          3642 => x"803982bb",
          3643 => x"a408f805",
          3644 => x"3353af73",
          3645 => x"27903882",
          3646 => x"bba408f8",
          3647 => x"05335372",
          3648 => x"b9268338",
          3649 => x"8d39800b",
          3650 => x"82bba408",
          3651 => x"ec050c82",
          3652 => x"d839880b",
          3653 => x"82bba408",
          3654 => x"f40534b2",
          3655 => x"3982bba4",
          3656 => x"08f80533",
          3657 => x"53af7327",
          3658 => x"903882bb",
          3659 => x"a408f805",
          3660 => x"335372b9",
          3661 => x"2683388d",
          3662 => x"39800b82",
          3663 => x"bba408ec",
          3664 => x"050c82a5",
          3665 => x"398a0b82",
          3666 => x"bba408f4",
          3667 => x"0534800b",
          3668 => x"82bba408",
          3669 => x"fc050c82",
          3670 => x"bba408f8",
          3671 => x"053353a0",
          3672 => x"732781cf",
          3673 => x"3882bba4",
          3674 => x"08f80533",
          3675 => x"5380e073",
          3676 => x"27943882",
          3677 => x"bba408f8",
          3678 => x"0533e011",
          3679 => x"51537282",
          3680 => x"bba408f8",
          3681 => x"053482bb",
          3682 => x"a408f805",
          3683 => x"33d01151",
          3684 => x"537282bb",
          3685 => x"a408f805",
          3686 => x"3482bba4",
          3687 => x"08f80533",
          3688 => x"53907327",
          3689 => x"ad3882bb",
          3690 => x"a408f805",
          3691 => x"33f91151",
          3692 => x"537282bb",
          3693 => x"a408f805",
          3694 => x"3482bba4",
          3695 => x"08f80533",
          3696 => x"53728926",
          3697 => x"8d38800b",
          3698 => x"82bba408",
          3699 => x"ec050c81",
          3700 => x"983982bb",
          3701 => x"a408f805",
          3702 => x"3382bba4",
          3703 => x"08f40533",
          3704 => x"54547274",
          3705 => x"268d3880",
          3706 => x"0b82bba4",
          3707 => x"08ec050c",
          3708 => x"80f73982",
          3709 => x"bba408f4",
          3710 => x"05337082",
          3711 => x"bba408fc",
          3712 => x"05082982",
          3713 => x"bba408f8",
          3714 => x"05337012",
          3715 => x"82bba408",
          3716 => x"fc050c82",
          3717 => x"bba40888",
          3718 => x"05087008",
          3719 => x"8105710c",
          3720 => x"70085151",
          3721 => x"52555372",
          3722 => x"3382bba4",
          3723 => x"08f80534",
          3724 => x"fea53982",
          3725 => x"bba408f0",
          3726 => x"05335372",
          3727 => x"802e9038",
          3728 => x"82bba408",
          3729 => x"fc050830",
          3730 => x"82bba408",
          3731 => x"fc050c82",
          3732 => x"bba4088c",
          3733 => x"050882bb",
          3734 => x"a408fc05",
          3735 => x"08710c53",
          3736 => x"810b82bb",
          3737 => x"a408ec05",
          3738 => x"0c82bba4",
          3739 => x"08ec0508",
          3740 => x"82bb980c",
          3741 => x"8b3d0d82",
          3742 => x"bba40c04",
          3743 => x"82bba408",
          3744 => x"0282bba4",
          3745 => x"0cfd3d0d",
          3746 => x"82d2e808",
          3747 => x"5382bba4",
          3748 => x"088c0508",
          3749 => x"5282bba4",
          3750 => x"08880508",
          3751 => x"51df8c3f",
          3752 => x"82bb9808",
          3753 => x"7082bb98",
          3754 => x"0c54853d",
          3755 => x"0d82bba4",
          3756 => x"0c0482bb",
          3757 => x"a4080282",
          3758 => x"bba40cf7",
          3759 => x"3d0d800b",
          3760 => x"82bba408",
          3761 => x"f0053482",
          3762 => x"bba4088c",
          3763 => x"05085380",
          3764 => x"730c82bb",
          3765 => x"a4088805",
          3766 => x"08700851",
          3767 => x"53723353",
          3768 => x"7282bba4",
          3769 => x"08f80534",
          3770 => x"7281ff06",
          3771 => x"5372a02e",
          3772 => x"09810691",
          3773 => x"3882bba4",
          3774 => x"08880508",
          3775 => x"70088105",
          3776 => x"710c53ce",
          3777 => x"3982bba4",
          3778 => x"08f80533",
          3779 => x"5372ad2e",
          3780 => x"098106a4",
          3781 => x"38810b82",
          3782 => x"bba408f0",
          3783 => x"053482bb",
          3784 => x"a4088805",
          3785 => x"08700881",
          3786 => x"05710c70",
          3787 => x"08515372",
          3788 => x"3382bba4",
          3789 => x"08f80534",
          3790 => x"82bba408",
          3791 => x"f8053353",
          3792 => x"72b02e09",
          3793 => x"810681dc",
          3794 => x"3882bba4",
          3795 => x"08880508",
          3796 => x"70088105",
          3797 => x"710c7008",
          3798 => x"51537233",
          3799 => x"82bba408",
          3800 => x"f8053482",
          3801 => x"bba408f8",
          3802 => x"053382bb",
          3803 => x"a408e805",
          3804 => x"0c82bba4",
          3805 => x"08e80508",
          3806 => x"80e22eb6",
          3807 => x"3882bba4",
          3808 => x"08e80508",
          3809 => x"80f82e84",
          3810 => x"3880cd39",
          3811 => x"900b82bb",
          3812 => x"a408f405",
          3813 => x"3482bba4",
          3814 => x"08880508",
          3815 => x"70088105",
          3816 => x"710c7008",
          3817 => x"51537233",
          3818 => x"82bba408",
          3819 => x"f8053481",
          3820 => x"a439820b",
          3821 => x"82bba408",
          3822 => x"f4053482",
          3823 => x"bba40888",
          3824 => x"05087008",
          3825 => x"8105710c",
          3826 => x"70085153",
          3827 => x"723382bb",
          3828 => x"a408f805",
          3829 => x"3480fe39",
          3830 => x"82bba408",
          3831 => x"f8053353",
          3832 => x"72a0268d",
          3833 => x"38810b82",
          3834 => x"bba408ec",
          3835 => x"050c8380",
          3836 => x"3982bba4",
          3837 => x"08f80533",
          3838 => x"53af7327",
          3839 => x"903882bb",
          3840 => x"a408f805",
          3841 => x"335372b9",
          3842 => x"2683388d",
          3843 => x"39800b82",
          3844 => x"bba408ec",
          3845 => x"050c82d8",
          3846 => x"39880b82",
          3847 => x"bba408f4",
          3848 => x"0534b239",
          3849 => x"82bba408",
          3850 => x"f8053353",
          3851 => x"af732790",
          3852 => x"3882bba4",
          3853 => x"08f80533",
          3854 => x"5372b926",
          3855 => x"83388d39",
          3856 => x"800b82bb",
          3857 => x"a408ec05",
          3858 => x"0c82a539",
          3859 => x"8a0b82bb",
          3860 => x"a408f405",
          3861 => x"34800b82",
          3862 => x"bba408fc",
          3863 => x"050c82bb",
          3864 => x"a408f805",
          3865 => x"3353a073",
          3866 => x"2781cf38",
          3867 => x"82bba408",
          3868 => x"f8053353",
          3869 => x"80e07327",
          3870 => x"943882bb",
          3871 => x"a408f805",
          3872 => x"33e01151",
          3873 => x"537282bb",
          3874 => x"a408f805",
          3875 => x"3482bba4",
          3876 => x"08f80533",
          3877 => x"d0115153",
          3878 => x"7282bba4",
          3879 => x"08f80534",
          3880 => x"82bba408",
          3881 => x"f8053353",
          3882 => x"907327ad",
          3883 => x"3882bba4",
          3884 => x"08f80533",
          3885 => x"f9115153",
          3886 => x"7282bba4",
          3887 => x"08f80534",
          3888 => x"82bba408",
          3889 => x"f8053353",
          3890 => x"7289268d",
          3891 => x"38800b82",
          3892 => x"bba408ec",
          3893 => x"050c8198",
          3894 => x"3982bba4",
          3895 => x"08f80533",
          3896 => x"82bba408",
          3897 => x"f4053354",
          3898 => x"54727426",
          3899 => x"8d38800b",
          3900 => x"82bba408",
          3901 => x"ec050c80",
          3902 => x"f73982bb",
          3903 => x"a408f405",
          3904 => x"337082bb",
          3905 => x"a408fc05",
          3906 => x"082982bb",
          3907 => x"a408f805",
          3908 => x"33701282",
          3909 => x"bba408fc",
          3910 => x"050c82bb",
          3911 => x"a4088805",
          3912 => x"08700881",
          3913 => x"05710c70",
          3914 => x"08515152",
          3915 => x"55537233",
          3916 => x"82bba408",
          3917 => x"f80534fe",
          3918 => x"a53982bb",
          3919 => x"a408f005",
          3920 => x"33537280",
          3921 => x"2e903882",
          3922 => x"bba408fc",
          3923 => x"05083082",
          3924 => x"bba408fc",
          3925 => x"050c82bb",
          3926 => x"a4088c05",
          3927 => x"0882bba4",
          3928 => x"08fc0508",
          3929 => x"710c5381",
          3930 => x"0b82bba4",
          3931 => x"08ec050c",
          3932 => x"82bba408",
          3933 => x"ec050882",
          3934 => x"bb980c8b",
          3935 => x"3d0d82bb",
          3936 => x"a40c0482",
          3937 => x"bba40802",
          3938 => x"82bba40c",
          3939 => x"fb3d0d80",
          3940 => x"0b82bba4",
          3941 => x"08f8050c",
          3942 => x"82d2ec08",
          3943 => x"85113370",
          3944 => x"812a7081",
          3945 => x"32708106",
          3946 => x"51515151",
          3947 => x"5372802e",
          3948 => x"8d38ff0b",
          3949 => x"82bba408",
          3950 => x"f4050c81",
          3951 => x"923982bb",
          3952 => x"a4088805",
          3953 => x"08537233",
          3954 => x"82bba408",
          3955 => x"88050881",
          3956 => x"0582bba4",
          3957 => x"0888050c",
          3958 => x"537282bb",
          3959 => x"a408fc05",
          3960 => x"347281ff",
          3961 => x"06537280",
          3962 => x"2eb03882",
          3963 => x"d2ec0882",
          3964 => x"d2ec0853",
          3965 => x"82bba408",
          3966 => x"fc053352",
          3967 => x"90110851",
          3968 => x"53722d82",
          3969 => x"bb980853",
          3970 => x"72802eff",
          3971 => x"b138ff0b",
          3972 => x"82bba408",
          3973 => x"f8050cff",
          3974 => x"a53982d2",
          3975 => x"ec0882d2",
          3976 => x"ec085353",
          3977 => x"8a519013",
          3978 => x"0853722d",
          3979 => x"82bb9808",
          3980 => x"5372802e",
          3981 => x"8a38ff0b",
          3982 => x"82bba408",
          3983 => x"f8050c82",
          3984 => x"bba408f8",
          3985 => x"05087082",
          3986 => x"bba408f4",
          3987 => x"050c5382",
          3988 => x"bba408f4",
          3989 => x"050882bb",
          3990 => x"980c873d",
          3991 => x"0d82bba4",
          3992 => x"0c0482bb",
          3993 => x"a4080282",
          3994 => x"bba40cfb",
          3995 => x"3d0d800b",
          3996 => x"82bba408",
          3997 => x"f8050c82",
          3998 => x"bba4088c",
          3999 => x"05088511",
          4000 => x"3370812a",
          4001 => x"70813270",
          4002 => x"81065151",
          4003 => x"51515372",
          4004 => x"802e8d38",
          4005 => x"ff0b82bb",
          4006 => x"a408f405",
          4007 => x"0c80f339",
          4008 => x"82bba408",
          4009 => x"88050853",
          4010 => x"723382bb",
          4011 => x"a4088805",
          4012 => x"08810582",
          4013 => x"bba40888",
          4014 => x"050c5372",
          4015 => x"82bba408",
          4016 => x"fc053472",
          4017 => x"81ff0653",
          4018 => x"72802eb6",
          4019 => x"3882bba4",
          4020 => x"088c0508",
          4021 => x"82bba408",
          4022 => x"8c050853",
          4023 => x"82bba408",
          4024 => x"fc053352",
          4025 => x"90110851",
          4026 => x"53722d82",
          4027 => x"bb980853",
          4028 => x"72802eff",
          4029 => x"ab38ff0b",
          4030 => x"82bba408",
          4031 => x"f8050cff",
          4032 => x"9f3982bb",
          4033 => x"a408f805",
          4034 => x"087082bb",
          4035 => x"a408f405",
          4036 => x"0c5382bb",
          4037 => x"a408f405",
          4038 => x"0882bb98",
          4039 => x"0c873d0d",
          4040 => x"82bba40c",
          4041 => x"0482bba4",
          4042 => x"080282bb",
          4043 => x"a40cfe3d",
          4044 => x"0d82d2ec",
          4045 => x"085282bb",
          4046 => x"a4088805",
          4047 => x"0851933f",
          4048 => x"82bb9808",
          4049 => x"7082bb98",
          4050 => x"0c53843d",
          4051 => x"0d82bba4",
          4052 => x"0c0482bb",
          4053 => x"a4080282",
          4054 => x"bba40cfb",
          4055 => x"3d0d82bb",
          4056 => x"a4088c05",
          4057 => x"08851133",
          4058 => x"70812a70",
          4059 => x"81327081",
          4060 => x"06515151",
          4061 => x"51537280",
          4062 => x"2e8d38ff",
          4063 => x"0b82bba4",
          4064 => x"08fc050c",
          4065 => x"81cb3982",
          4066 => x"bba4088c",
          4067 => x"05088511",
          4068 => x"3370822a",
          4069 => x"70810651",
          4070 => x"51515372",
          4071 => x"802e80db",
          4072 => x"3882bba4",
          4073 => x"088c0508",
          4074 => x"82bba408",
          4075 => x"8c050854",
          4076 => x"548c1408",
          4077 => x"88140825",
          4078 => x"9f3882bb",
          4079 => x"a4088c05",
          4080 => x"08700870",
          4081 => x"82bba408",
          4082 => x"88050852",
          4083 => x"57545472",
          4084 => x"75347308",
          4085 => x"8105740c",
          4086 => x"82bba408",
          4087 => x"8c05088c",
          4088 => x"11088105",
          4089 => x"8c120c82",
          4090 => x"bba40888",
          4091 => x"05087082",
          4092 => x"bba408fc",
          4093 => x"050c5153",
          4094 => x"80d73982",
          4095 => x"bba4088c",
          4096 => x"050882bb",
          4097 => x"a4088c05",
          4098 => x"085382bb",
          4099 => x"a4088805",
          4100 => x"087081ff",
          4101 => x"06539012",
          4102 => x"08515454",
          4103 => x"722d82bb",
          4104 => x"98085372",
          4105 => x"a33882bb",
          4106 => x"a4088c05",
          4107 => x"088c1108",
          4108 => x"81058c12",
          4109 => x"0c82bba4",
          4110 => x"08880508",
          4111 => x"7082bba4",
          4112 => x"08fc050c",
          4113 => x"51538a39",
          4114 => x"ff0b82bb",
          4115 => x"a408fc05",
          4116 => x"0c82bba4",
          4117 => x"08fc0508",
          4118 => x"82bb980c",
          4119 => x"873d0d82",
          4120 => x"bba40c04",
          4121 => x"82bba408",
          4122 => x"0282bba4",
          4123 => x"0cf93d0d",
          4124 => x"82bba408",
          4125 => x"88050885",
          4126 => x"11337081",
          4127 => x"32708106",
          4128 => x"51515152",
          4129 => x"71802e8d",
          4130 => x"38ff0b82",
          4131 => x"bba408f8",
          4132 => x"050c8394",
          4133 => x"3982bba4",
          4134 => x"08880508",
          4135 => x"85113370",
          4136 => x"862a7081",
          4137 => x"06515151",
          4138 => x"5271802e",
          4139 => x"80c53882",
          4140 => x"bba40888",
          4141 => x"050882bb",
          4142 => x"a4088805",
          4143 => x"08535385",
          4144 => x"123370ff",
          4145 => x"bf065152",
          4146 => x"71851434",
          4147 => x"82bba408",
          4148 => x"8805088c",
          4149 => x"11088105",
          4150 => x"8c120c82",
          4151 => x"bba40888",
          4152 => x"05088411",
          4153 => x"337082bb",
          4154 => x"a408f805",
          4155 => x"0c515152",
          4156 => x"82b63982",
          4157 => x"bba40888",
          4158 => x"05088511",
          4159 => x"3370822a",
          4160 => x"70810651",
          4161 => x"51515271",
          4162 => x"802e80d7",
          4163 => x"3882bba4",
          4164 => x"08880508",
          4165 => x"70087033",
          4166 => x"82bba408",
          4167 => x"fc050c51",
          4168 => x"5282bba4",
          4169 => x"08fc0508",
          4170 => x"a93882bb",
          4171 => x"a4088805",
          4172 => x"0882bba4",
          4173 => x"08880508",
          4174 => x"53538512",
          4175 => x"3370a007",
          4176 => x"51527185",
          4177 => x"1434ff0b",
          4178 => x"82bba408",
          4179 => x"f8050c81",
          4180 => x"d73982bb",
          4181 => x"a4088805",
          4182 => x"08700881",
          4183 => x"05710c52",
          4184 => x"81a13982",
          4185 => x"bba40888",
          4186 => x"050882bb",
          4187 => x"a4088805",
          4188 => x"08529411",
          4189 => x"08515271",
          4190 => x"2d82bb98",
          4191 => x"087082bb",
          4192 => x"a408fc05",
          4193 => x"0c5282bb",
          4194 => x"a408fc05",
          4195 => x"08802580",
          4196 => x"f23882bb",
          4197 => x"a4088805",
          4198 => x"0882bba4",
          4199 => x"08f4050c",
          4200 => x"82bba408",
          4201 => x"88050885",
          4202 => x"113382bb",
          4203 => x"a408f005",
          4204 => x"0c5282bb",
          4205 => x"a408fc05",
          4206 => x"08ff2e09",
          4207 => x"81069538",
          4208 => x"82bba408",
          4209 => x"f0050890",
          4210 => x"07527182",
          4211 => x"bba408ec",
          4212 => x"05349339",
          4213 => x"82bba408",
          4214 => x"f00508a0",
          4215 => x"07527182",
          4216 => x"bba408ec",
          4217 => x"053482bb",
          4218 => x"a408f405",
          4219 => x"085282bb",
          4220 => x"a408ec05",
          4221 => x"33851334",
          4222 => x"ff0b82bb",
          4223 => x"a408f805",
          4224 => x"0ca63982",
          4225 => x"bba40888",
          4226 => x"05088c11",
          4227 => x"0881058c",
          4228 => x"120c82bb",
          4229 => x"a408fc05",
          4230 => x"087081ff",
          4231 => x"067082bb",
          4232 => x"a408f805",
          4233 => x"0c515152",
          4234 => x"82bba408",
          4235 => x"f8050882",
          4236 => x"bb980c89",
          4237 => x"3d0d82bb",
          4238 => x"a40c0482",
          4239 => x"bba40802",
          4240 => x"82bba40c",
          4241 => x"fd3d0d82",
          4242 => x"bba40888",
          4243 => x"050882bb",
          4244 => x"a408fc05",
          4245 => x"0c82bba4",
          4246 => x"088c0508",
          4247 => x"82bba408",
          4248 => x"f8050c82",
          4249 => x"bba40890",
          4250 => x"0508802e",
          4251 => x"82a23882",
          4252 => x"bba408f8",
          4253 => x"050882bb",
          4254 => x"a408fc05",
          4255 => x"082681ac",
          4256 => x"3882bba4",
          4257 => x"08f80508",
          4258 => x"82bba408",
          4259 => x"90050805",
          4260 => x"5182bba4",
          4261 => x"08fc0508",
          4262 => x"71278190",
          4263 => x"3882bba4",
          4264 => x"08fc0508",
          4265 => x"82bba408",
          4266 => x"90050805",
          4267 => x"82bba408",
          4268 => x"fc050c82",
          4269 => x"bba408f8",
          4270 => x"050882bb",
          4271 => x"a4089005",
          4272 => x"080582bb",
          4273 => x"a408f805",
          4274 => x"0c82bba4",
          4275 => x"08900508",
          4276 => x"810582bb",
          4277 => x"a4089005",
          4278 => x"0c82bba4",
          4279 => x"08900508",
          4280 => x"ff0582bb",
          4281 => x"a4089005",
          4282 => x"0c82bba4",
          4283 => x"08900508",
          4284 => x"802e819c",
          4285 => x"3882bba4",
          4286 => x"08fc0508",
          4287 => x"ff0582bb",
          4288 => x"a408fc05",
          4289 => x"0c82bba4",
          4290 => x"08f80508",
          4291 => x"ff0582bb",
          4292 => x"a408f805",
          4293 => x"0c82bba4",
          4294 => x"08fc0508",
          4295 => x"82bba408",
          4296 => x"f8050853",
          4297 => x"51713371",
          4298 => x"34ffae39",
          4299 => x"82bba408",
          4300 => x"90050881",
          4301 => x"0582bba4",
          4302 => x"0890050c",
          4303 => x"82bba408",
          4304 => x"900508ff",
          4305 => x"0582bba4",
          4306 => x"0890050c",
          4307 => x"82bba408",
          4308 => x"90050880",
          4309 => x"2eba3882",
          4310 => x"bba408f8",
          4311 => x"05085170",
          4312 => x"3382bba4",
          4313 => x"08f80508",
          4314 => x"810582bb",
          4315 => x"a408f805",
          4316 => x"0c82bba4",
          4317 => x"08fc0508",
          4318 => x"52527171",
          4319 => x"3482bba4",
          4320 => x"08fc0508",
          4321 => x"810582bb",
          4322 => x"a408fc05",
          4323 => x"0cffad39",
          4324 => x"82bba408",
          4325 => x"88050870",
          4326 => x"82bb980c",
          4327 => x"51853d0d",
          4328 => x"82bba40c",
          4329 => x"0482bba4",
          4330 => x"080282bb",
          4331 => x"a40cfe3d",
          4332 => x"0d82bba4",
          4333 => x"08880508",
          4334 => x"82bba408",
          4335 => x"fc050c82",
          4336 => x"bba408fc",
          4337 => x"05085271",
          4338 => x"3382bba4",
          4339 => x"08fc0508",
          4340 => x"810582bb",
          4341 => x"a408fc05",
          4342 => x"0c7081ff",
          4343 => x"06515170",
          4344 => x"802e8338",
          4345 => x"da3982bb",
          4346 => x"a408fc05",
          4347 => x"08ff0582",
          4348 => x"bba408fc",
          4349 => x"050c82bb",
          4350 => x"a408fc05",
          4351 => x"0882bba4",
          4352 => x"08880508",
          4353 => x"317082bb",
          4354 => x"980c5184",
          4355 => x"3d0d82bb",
          4356 => x"a40c0482",
          4357 => x"bba40802",
          4358 => x"82bba40c",
          4359 => x"fe3d0d82",
          4360 => x"bba40888",
          4361 => x"050882bb",
          4362 => x"a408fc05",
          4363 => x"0c82bba4",
          4364 => x"088c0508",
          4365 => x"52713382",
          4366 => x"bba4088c",
          4367 => x"05088105",
          4368 => x"82bba408",
          4369 => x"8c050c82",
          4370 => x"bba408fc",
          4371 => x"05085351",
          4372 => x"70723482",
          4373 => x"bba408fc",
          4374 => x"05088105",
          4375 => x"82bba408",
          4376 => x"fc050c70",
          4377 => x"81ff0651",
          4378 => x"70802e84",
          4379 => x"38ffbe39",
          4380 => x"82bba408",
          4381 => x"88050870",
          4382 => x"82bb980c",
          4383 => x"51843d0d",
          4384 => x"82bba40c",
          4385 => x"0482bba4",
          4386 => x"080282bb",
          4387 => x"a40cfd3d",
          4388 => x"0d82bba4",
          4389 => x"08880508",
          4390 => x"82bba408",
          4391 => x"fc050c82",
          4392 => x"bba4088c",
          4393 => x"050882bb",
          4394 => x"a408f805",
          4395 => x"0c82bba4",
          4396 => x"08900508",
          4397 => x"802e80e5",
          4398 => x"3882bba4",
          4399 => x"08900508",
          4400 => x"810582bb",
          4401 => x"a4089005",
          4402 => x"0c82bba4",
          4403 => x"08900508",
          4404 => x"ff0582bb",
          4405 => x"a4089005",
          4406 => x"0c82bba4",
          4407 => x"08900508",
          4408 => x"802eba38",
          4409 => x"82bba408",
          4410 => x"f8050851",
          4411 => x"703382bb",
          4412 => x"a408f805",
          4413 => x"08810582",
          4414 => x"bba408f8",
          4415 => x"050c82bb",
          4416 => x"a408fc05",
          4417 => x"08525271",
          4418 => x"713482bb",
          4419 => x"a408fc05",
          4420 => x"08810582",
          4421 => x"bba408fc",
          4422 => x"050cffad",
          4423 => x"3982bba4",
          4424 => x"08880508",
          4425 => x"7082bb98",
          4426 => x"0c51853d",
          4427 => x"0d82bba4",
          4428 => x"0c0482bb",
          4429 => x"a4080282",
          4430 => x"bba40cfd",
          4431 => x"3d0d82bb",
          4432 => x"a4089005",
          4433 => x"08802e81",
          4434 => x"f43882bb",
          4435 => x"a4088c05",
          4436 => x"08527133",
          4437 => x"82bba408",
          4438 => x"8c050881",
          4439 => x"0582bba4",
          4440 => x"088c050c",
          4441 => x"82bba408",
          4442 => x"88050870",
          4443 => x"337281ff",
          4444 => x"06535454",
          4445 => x"5171712e",
          4446 => x"843880ce",
          4447 => x"3982bba4",
          4448 => x"08880508",
          4449 => x"52713382",
          4450 => x"bba40888",
          4451 => x"05088105",
          4452 => x"82bba408",
          4453 => x"88050c70",
          4454 => x"81ff0651",
          4455 => x"51708d38",
          4456 => x"800b82bb",
          4457 => x"a408fc05",
          4458 => x"0c819b39",
          4459 => x"82bba408",
          4460 => x"900508ff",
          4461 => x"0582bba4",
          4462 => x"0890050c",
          4463 => x"82bba408",
          4464 => x"90050880",
          4465 => x"2e8438ff",
          4466 => x"813982bb",
          4467 => x"a4089005",
          4468 => x"08802e80",
          4469 => x"e83882bb",
          4470 => x"a4088805",
          4471 => x"08703352",
          4472 => x"53708d38",
          4473 => x"ff0b82bb",
          4474 => x"a408fc05",
          4475 => x"0c80d739",
          4476 => x"82bba408",
          4477 => x"8c0508ff",
          4478 => x"0582bba4",
          4479 => x"088c050c",
          4480 => x"82bba408",
          4481 => x"8c050870",
          4482 => x"33525270",
          4483 => x"8c38810b",
          4484 => x"82bba408",
          4485 => x"fc050cae",
          4486 => x"3982bba4",
          4487 => x"08880508",
          4488 => x"703382bb",
          4489 => x"a4088c05",
          4490 => x"08703372",
          4491 => x"71317082",
          4492 => x"bba408fc",
          4493 => x"050c5355",
          4494 => x"5252538a",
          4495 => x"39800b82",
          4496 => x"bba408fc",
          4497 => x"050c82bb",
          4498 => x"a408fc05",
          4499 => x"0882bb98",
          4500 => x"0c853d0d",
          4501 => x"82bba40c",
          4502 => x"0482bba4",
          4503 => x"080282bb",
          4504 => x"a40cfd3d",
          4505 => x"0d82bba4",
          4506 => x"08880508",
          4507 => x"82bba408",
          4508 => x"f8050c82",
          4509 => x"bba4088c",
          4510 => x"05088d38",
          4511 => x"800b82bb",
          4512 => x"a408fc05",
          4513 => x"0c80ec39",
          4514 => x"82bba408",
          4515 => x"f8050852",
          4516 => x"713382bb",
          4517 => x"a408f805",
          4518 => x"08810582",
          4519 => x"bba408f8",
          4520 => x"050c7081",
          4521 => x"ff065151",
          4522 => x"70802e9f",
          4523 => x"3882bba4",
          4524 => x"088c0508",
          4525 => x"ff0582bb",
          4526 => x"a4088c05",
          4527 => x"0c82bba4",
          4528 => x"088c0508",
          4529 => x"ff2e8438",
          4530 => x"ffbe3982",
          4531 => x"bba408f8",
          4532 => x"0508ff05",
          4533 => x"82bba408",
          4534 => x"f8050c82",
          4535 => x"bba408f8",
          4536 => x"050882bb",
          4537 => x"a4088805",
          4538 => x"08317082",
          4539 => x"bba408fc",
          4540 => x"050c5182",
          4541 => x"bba408fc",
          4542 => x"050882bb",
          4543 => x"980c853d",
          4544 => x"0d82bba4",
          4545 => x"0c0482bb",
          4546 => x"a4080282",
          4547 => x"bba40cfe",
          4548 => x"3d0d82bb",
          4549 => x"a4088805",
          4550 => x"0882bba4",
          4551 => x"08fc050c",
          4552 => x"82bba408",
          4553 => x"90050880",
          4554 => x"2e80d438",
          4555 => x"82bba408",
          4556 => x"90050881",
          4557 => x"0582bba4",
          4558 => x"0890050c",
          4559 => x"82bba408",
          4560 => x"900508ff",
          4561 => x"0582bba4",
          4562 => x"0890050c",
          4563 => x"82bba408",
          4564 => x"90050880",
          4565 => x"2ea93882",
          4566 => x"bba4088c",
          4567 => x"05085170",
          4568 => x"82bba408",
          4569 => x"fc050852",
          4570 => x"52717134",
          4571 => x"82bba408",
          4572 => x"fc050881",
          4573 => x"0582bba4",
          4574 => x"08fc050c",
          4575 => x"ffbe3982",
          4576 => x"bba40888",
          4577 => x"05087082",
          4578 => x"bb980c51",
          4579 => x"843d0d82",
          4580 => x"bba40c04",
          4581 => x"82bba408",
          4582 => x"0282bba4",
          4583 => x"0cf93d0d",
          4584 => x"800b82bb",
          4585 => x"a408fc05",
          4586 => x"0c82bba4",
          4587 => x"08880508",
          4588 => x"8025b938",
          4589 => x"82bba408",
          4590 => x"88050830",
          4591 => x"82bba408",
          4592 => x"88050c80",
          4593 => x"0b82bba4",
          4594 => x"08f4050c",
          4595 => x"82bba408",
          4596 => x"fc05088a",
          4597 => x"38810b82",
          4598 => x"bba408f4",
          4599 => x"050c82bb",
          4600 => x"a408f405",
          4601 => x"0882bba4",
          4602 => x"08fc050c",
          4603 => x"82bba408",
          4604 => x"8c050880",
          4605 => x"25b93882",
          4606 => x"bba4088c",
          4607 => x"05083082",
          4608 => x"bba4088c",
          4609 => x"050c800b",
          4610 => x"82bba408",
          4611 => x"f0050c82",
          4612 => x"bba408fc",
          4613 => x"05088a38",
          4614 => x"810b82bb",
          4615 => x"a408f005",
          4616 => x"0c82bba4",
          4617 => x"08f00508",
          4618 => x"82bba408",
          4619 => x"fc050c80",
          4620 => x"5382bba4",
          4621 => x"088c0508",
          4622 => x"5282bba4",
          4623 => x"08880508",
          4624 => x"5182c53f",
          4625 => x"82bb9808",
          4626 => x"7082bba4",
          4627 => x"08f8050c",
          4628 => x"5482bba4",
          4629 => x"08fc0508",
          4630 => x"802e9038",
          4631 => x"82bba408",
          4632 => x"f8050830",
          4633 => x"82bba408",
          4634 => x"f8050c82",
          4635 => x"bba408f8",
          4636 => x"05087082",
          4637 => x"bb980c54",
          4638 => x"893d0d82",
          4639 => x"bba40c04",
          4640 => x"82bba408",
          4641 => x"0282bba4",
          4642 => x"0cfb3d0d",
          4643 => x"800b82bb",
          4644 => x"a408fc05",
          4645 => x"0c82bba4",
          4646 => x"08880508",
          4647 => x"80259938",
          4648 => x"82bba408",
          4649 => x"88050830",
          4650 => x"82bba408",
          4651 => x"88050c81",
          4652 => x"0b82bba4",
          4653 => x"08fc050c",
          4654 => x"82bba408",
          4655 => x"8c050880",
          4656 => x"25903882",
          4657 => x"bba4088c",
          4658 => x"05083082",
          4659 => x"bba4088c",
          4660 => x"050c8153",
          4661 => x"82bba408",
          4662 => x"8c050852",
          4663 => x"82bba408",
          4664 => x"88050851",
          4665 => x"81a23f82",
          4666 => x"bb980870",
          4667 => x"82bba408",
          4668 => x"f8050c54",
          4669 => x"82bba408",
          4670 => x"fc050880",
          4671 => x"2e903882",
          4672 => x"bba408f8",
          4673 => x"05083082",
          4674 => x"bba408f8",
          4675 => x"050c82bb",
          4676 => x"a408f805",
          4677 => x"087082bb",
          4678 => x"980c5487",
          4679 => x"3d0d82bb",
          4680 => x"a40c0482",
          4681 => x"bba40802",
          4682 => x"82bba40c",
          4683 => x"fd3d0d80",
          4684 => x"5382bba4",
          4685 => x"088c0508",
          4686 => x"5282bba4",
          4687 => x"08880508",
          4688 => x"5180c53f",
          4689 => x"82bb9808",
          4690 => x"7082bb98",
          4691 => x"0c54853d",
          4692 => x"0d82bba4",
          4693 => x"0c0482bb",
          4694 => x"a4080282",
          4695 => x"bba40cfd",
          4696 => x"3d0d8153",
          4697 => x"82bba408",
          4698 => x"8c050852",
          4699 => x"82bba408",
          4700 => x"88050851",
          4701 => x"933f82bb",
          4702 => x"98087082",
          4703 => x"bb980c54",
          4704 => x"853d0d82",
          4705 => x"bba40c04",
          4706 => x"82bba408",
          4707 => x"0282bba4",
          4708 => x"0cfd3d0d",
          4709 => x"810b82bb",
          4710 => x"a408fc05",
          4711 => x"0c800b82",
          4712 => x"bba408f8",
          4713 => x"050c82bb",
          4714 => x"a4088c05",
          4715 => x"0882bba4",
          4716 => x"08880508",
          4717 => x"27b93882",
          4718 => x"bba408fc",
          4719 => x"0508802e",
          4720 => x"ae38800b",
          4721 => x"82bba408",
          4722 => x"8c050824",
          4723 => x"a23882bb",
          4724 => x"a4088c05",
          4725 => x"081082bb",
          4726 => x"a4088c05",
          4727 => x"0c82bba4",
          4728 => x"08fc0508",
          4729 => x"1082bba4",
          4730 => x"08fc050c",
          4731 => x"ffb83982",
          4732 => x"bba408fc",
          4733 => x"0508802e",
          4734 => x"80e13882",
          4735 => x"bba4088c",
          4736 => x"050882bb",
          4737 => x"a4088805",
          4738 => x"0826ad38",
          4739 => x"82bba408",
          4740 => x"88050882",
          4741 => x"bba4088c",
          4742 => x"05083182",
          4743 => x"bba40888",
          4744 => x"050c82bb",
          4745 => x"a408f805",
          4746 => x"0882bba4",
          4747 => x"08fc0508",
          4748 => x"0782bba4",
          4749 => x"08f8050c",
          4750 => x"82bba408",
          4751 => x"fc050881",
          4752 => x"2a82bba4",
          4753 => x"08fc050c",
          4754 => x"82bba408",
          4755 => x"8c050881",
          4756 => x"2a82bba4",
          4757 => x"088c050c",
          4758 => x"ff953982",
          4759 => x"bba40890",
          4760 => x"0508802e",
          4761 => x"933882bb",
          4762 => x"a4088805",
          4763 => x"087082bb",
          4764 => x"a408f405",
          4765 => x"0c519139",
          4766 => x"82bba408",
          4767 => x"f8050870",
          4768 => x"82bba408",
          4769 => x"f4050c51",
          4770 => x"82bba408",
          4771 => x"f4050882",
          4772 => x"bb980c85",
          4773 => x"3d0d82bb",
          4774 => x"a40c04f9",
          4775 => x"3d0d7970",
          4776 => x"08705656",
          4777 => x"5874802e",
          4778 => x"80e33895",
          4779 => x"39750851",
          4780 => x"f1f33f82",
          4781 => x"bb980815",
          4782 => x"780c8516",
          4783 => x"335480cd",
          4784 => x"39743354",
          4785 => x"73a02e09",
          4786 => x"81068638",
          4787 => x"811555f1",
          4788 => x"39805776",
          4789 => x"902982b6",
          4790 => x"98057008",
          4791 => x"5256f1c5",
          4792 => x"3f82bb98",
          4793 => x"08537452",
          4794 => x"750851f4",
          4795 => x"c53f82bb",
          4796 => x"98088b38",
          4797 => x"84163354",
          4798 => x"73812eff",
          4799 => x"b0388117",
          4800 => x"7081ff06",
          4801 => x"58549977",
          4802 => x"27c938ff",
          4803 => x"547382bb",
          4804 => x"980c893d",
          4805 => x"0d04ff3d",
          4806 => x"0d735271",
          4807 => x"9326818e",
          4808 => x"38718429",
          4809 => x"8299b005",
          4810 => x"52710804",
          4811 => x"829efc51",
          4812 => x"81803982",
          4813 => x"9f885180",
          4814 => x"f939829f",
          4815 => x"9c5180f2",
          4816 => x"39829fb0",
          4817 => x"5180eb39",
          4818 => x"829fc051",
          4819 => x"80e43982",
          4820 => x"9fd05180",
          4821 => x"dd39829f",
          4822 => x"e45180d6",
          4823 => x"39829ff4",
          4824 => x"5180cf39",
          4825 => x"82a08c51",
          4826 => x"80c83982",
          4827 => x"a0a45180",
          4828 => x"c13982a0",
          4829 => x"bc51bb39",
          4830 => x"82a0d851",
          4831 => x"b53982a0",
          4832 => x"ec51af39",
          4833 => x"82a19851",
          4834 => x"a93982a1",
          4835 => x"ac51a339",
          4836 => x"82a1cc51",
          4837 => x"9d3982a1",
          4838 => x"e0519739",
          4839 => x"82a1f851",
          4840 => x"913982a2",
          4841 => x"90518b39",
          4842 => x"82a2a851",
          4843 => x"853982a2",
          4844 => x"b451e3cf",
          4845 => x"3f833d0d",
          4846 => x"04fb3d0d",
          4847 => x"77795656",
          4848 => x"7487e726",
          4849 => x"8a387452",
          4850 => x"7587e829",
          4851 => x"51903987",
          4852 => x"e8527451",
          4853 => x"facd3f82",
          4854 => x"bb980852",
          4855 => x"7551fac3",
          4856 => x"3f82bb98",
          4857 => x"08547953",
          4858 => x"755282a2",
          4859 => x"c451ffbb",
          4860 => x"e53f873d",
          4861 => x"0d04ec3d",
          4862 => x"0d660284",
          4863 => x"0580e305",
          4864 => x"335b5780",
          4865 => x"68783070",
          4866 => x"7a077325",
          4867 => x"51575959",
          4868 => x"78567787",
          4869 => x"ff268338",
          4870 => x"81567476",
          4871 => x"077081ff",
          4872 => x"06515593",
          4873 => x"56748182",
          4874 => x"38815376",
          4875 => x"528c3d70",
          4876 => x"52568183",
          4877 => x"cf3f82bb",
          4878 => x"98085782",
          4879 => x"bb9808b9",
          4880 => x"3882bb98",
          4881 => x"0887c098",
          4882 => x"880c82bb",
          4883 => x"98085996",
          4884 => x"3dd40554",
          4885 => x"84805377",
          4886 => x"52755181",
          4887 => x"888b3f82",
          4888 => x"bb980857",
          4889 => x"82bb9808",
          4890 => x"90387a55",
          4891 => x"74802e89",
          4892 => x"38741975",
          4893 => x"195959d7",
          4894 => x"39963dd8",
          4895 => x"0551818f",
          4896 => x"f43f7630",
          4897 => x"70780780",
          4898 => x"257b3070",
          4899 => x"9f2a7206",
          4900 => x"51575156",
          4901 => x"74802e90",
          4902 => x"3882a2e8",
          4903 => x"5387c098",
          4904 => x"88085278",
          4905 => x"51fe923f",
          4906 => x"76567582",
          4907 => x"bb980c96",
          4908 => x"3d0d04f8",
          4909 => x"3d0d7c02",
          4910 => x"8405b705",
          4911 => x"335859ff",
          4912 => x"5880537b",
          4913 => x"527a51fe",
          4914 => x"ad3f82bb",
          4915 => x"9808a638",
          4916 => x"76802e88",
          4917 => x"3876812e",
          4918 => x"9a389a39",
          4919 => x"62566155",
          4920 => x"605482bb",
          4921 => x"98537f52",
          4922 => x"7e51782d",
          4923 => x"82bb9808",
          4924 => x"58833978",
          4925 => x"047782bb",
          4926 => x"980c8a3d",
          4927 => x"0d04f33d",
          4928 => x"0d7f6163",
          4929 => x"028c0580",
          4930 => x"cf053373",
          4931 => x"73156841",
          4932 => x"5f5c5c5e",
          4933 => x"5e5e7a52",
          4934 => x"82a2f051",
          4935 => x"ffb9b73f",
          4936 => x"82a2f851",
          4937 => x"e0dd3f80",
          4938 => x"55747927",
          4939 => x"80fd387b",
          4940 => x"902e8938",
          4941 => x"7ba02ea6",
          4942 => x"3880c439",
          4943 => x"74185372",
          4944 => x"7a278e38",
          4945 => x"72225282",
          4946 => x"a2fc51ff",
          4947 => x"b9883f88",
          4948 => x"3982a388",
          4949 => x"51e0ac3f",
          4950 => x"82155580",
          4951 => x"c1397418",
          4952 => x"53727a27",
          4953 => x"8e387208",
          4954 => x"5282a2f0",
          4955 => x"51ffb8e6",
          4956 => x"3f883982",
          4957 => x"a38451e0",
          4958 => x"8a3f8415",
          4959 => x"55a03974",
          4960 => x"1853727a",
          4961 => x"278e3872",
          4962 => x"335282a3",
          4963 => x"9051ffb8",
          4964 => x"c53f8839",
          4965 => x"82a39851",
          4966 => x"dfe93f81",
          4967 => x"155582d2",
          4968 => x"ec0852a0",
          4969 => x"51e3ab3f",
          4970 => x"feff3982",
          4971 => x"a39c51df",
          4972 => x"d23f8055",
          4973 => x"74792780",
          4974 => x"c6387418",
          4975 => x"70335553",
          4976 => x"8056727a",
          4977 => x"27833881",
          4978 => x"5680539f",
          4979 => x"74278338",
          4980 => x"81537573",
          4981 => x"067081ff",
          4982 => x"06515372",
          4983 => x"802e9038",
          4984 => x"7380fe26",
          4985 => x"8a3882d2",
          4986 => x"ec085273",
          4987 => x"51883982",
          4988 => x"d2ec0852",
          4989 => x"a051e2da",
          4990 => x"3f811555",
          4991 => x"ffb63982",
          4992 => x"a3a051de",
          4993 => x"fe3f7818",
          4994 => x"791c5c58",
          4995 => x"a0ef3f82",
          4996 => x"bb980898",
          4997 => x"2b70982c",
          4998 => x"515776a0",
          4999 => x"2e098106",
          5000 => x"aa38a0d9",
          5001 => x"3f82bb98",
          5002 => x"08982b70",
          5003 => x"982c70a0",
          5004 => x"32703072",
          5005 => x"9b327030",
          5006 => x"70720773",
          5007 => x"75070651",
          5008 => x"58585957",
          5009 => x"51578073",
          5010 => x"24d83876",
          5011 => x"9b2e0981",
          5012 => x"06853880",
          5013 => x"538c397c",
          5014 => x"1e537278",
          5015 => x"26fdb738",
          5016 => x"ff537282",
          5017 => x"bb980c8f",
          5018 => x"3d0d04fc",
          5019 => x"3d0d029b",
          5020 => x"053382a3",
          5021 => x"a45382a3",
          5022 => x"ac5255ff",
          5023 => x"b6d83f82",
          5024 => x"b9f02251",
          5025 => x"a9ca3f82",
          5026 => x"a3b85482",
          5027 => x"a3c45382",
          5028 => x"b9f13352",
          5029 => x"82a3cc51",
          5030 => x"ffb6bb3f",
          5031 => x"74802e84",
          5032 => x"38a4fc3f",
          5033 => x"863d0d04",
          5034 => x"fe3d0d87",
          5035 => x"c0968008",
          5036 => x"53aaa73f",
          5037 => x"81519cb2",
          5038 => x"3f82a3e8",
          5039 => x"519dc73f",
          5040 => x"80519ca6",
          5041 => x"3f72812a",
          5042 => x"70810651",
          5043 => x"5271802e",
          5044 => x"92388151",
          5045 => x"9c943f82",
          5046 => x"a484519d",
          5047 => x"a93f8051",
          5048 => x"9c883f72",
          5049 => x"822a7081",
          5050 => x"06515271",
          5051 => x"802e9238",
          5052 => x"81519bf6",
          5053 => x"3f82a498",
          5054 => x"519d8b3f",
          5055 => x"80519bea",
          5056 => x"3f72832a",
          5057 => x"70810651",
          5058 => x"5271802e",
          5059 => x"92388151",
          5060 => x"9bd83f82",
          5061 => x"a4a8519c",
          5062 => x"ed3f8051",
          5063 => x"9bcc3f72",
          5064 => x"842a7081",
          5065 => x"06515271",
          5066 => x"802e9238",
          5067 => x"81519bba",
          5068 => x"3f82a4bc",
          5069 => x"519ccf3f",
          5070 => x"80519bae",
          5071 => x"3f72852a",
          5072 => x"70810651",
          5073 => x"5271802e",
          5074 => x"92388151",
          5075 => x"9b9c3f82",
          5076 => x"a4d0519c",
          5077 => x"b13f8051",
          5078 => x"9b903f72",
          5079 => x"862a7081",
          5080 => x"06515271",
          5081 => x"802e9238",
          5082 => x"81519afe",
          5083 => x"3f82a4e4",
          5084 => x"519c933f",
          5085 => x"80519af2",
          5086 => x"3f72872a",
          5087 => x"70810651",
          5088 => x"5271802e",
          5089 => x"92388151",
          5090 => x"9ae03f82",
          5091 => x"a4f8519b",
          5092 => x"f53f8051",
          5093 => x"9ad43f72",
          5094 => x"882a7081",
          5095 => x"06515271",
          5096 => x"802e9238",
          5097 => x"81519ac2",
          5098 => x"3f82a58c",
          5099 => x"519bd73f",
          5100 => x"80519ab6",
          5101 => x"3fa8ab3f",
          5102 => x"843d0d04",
          5103 => x"fb3d0d77",
          5104 => x"028405a3",
          5105 => x"05337055",
          5106 => x"56568052",
          5107 => x"7551eeb6",
          5108 => x"3f0b0b82",
          5109 => x"b6943354",
          5110 => x"73a93881",
          5111 => x"5382a5cc",
          5112 => x"5282d298",
          5113 => x"5180fc9c",
          5114 => x"3f82bb98",
          5115 => x"08307082",
          5116 => x"bb980807",
          5117 => x"80258271",
          5118 => x"31515154",
          5119 => x"730b0b82",
          5120 => x"b694340b",
          5121 => x"0b82b694",
          5122 => x"33547381",
          5123 => x"2e098106",
          5124 => x"af3882d2",
          5125 => x"98537452",
          5126 => x"755181b6",
          5127 => x"cd3f82bb",
          5128 => x"9808802e",
          5129 => x"8b3882bb",
          5130 => x"980851da",
          5131 => x"d63f9139",
          5132 => x"82d29851",
          5133 => x"8188be3f",
          5134 => x"820b0b0b",
          5135 => x"82b69434",
          5136 => x"0b0b82b6",
          5137 => x"94335473",
          5138 => x"822e0981",
          5139 => x"068c3882",
          5140 => x"a5dc5374",
          5141 => x"527551ae",
          5142 => x"953f800b",
          5143 => x"82bb980c",
          5144 => x"873d0d04",
          5145 => x"cd3d0d80",
          5146 => x"707182d2",
          5147 => x"940c405e",
          5148 => x"81527d51",
          5149 => x"80cae83f",
          5150 => x"82bb9808",
          5151 => x"81ff065a",
          5152 => x"797e2e09",
          5153 => x"8106a338",
          5154 => x"973d5a83",
          5155 => x"5382a5e8",
          5156 => x"527951e7",
          5157 => x"f03f7d53",
          5158 => x"795282bc",
          5159 => x"c45180fa",
          5160 => x"823f82bb",
          5161 => x"98087e2e",
          5162 => x"883882a5",
          5163 => x"ec5191c8",
          5164 => x"39817040",
          5165 => x"5e82a6a4",
          5166 => x"51d9c83f",
          5167 => x"973d7047",
          5168 => x"5b80f852",
          5169 => x"7a51fdf4",
          5170 => x"3fb53dff",
          5171 => x"840551f3",
          5172 => x"ca3f82bb",
          5173 => x"9808902b",
          5174 => x"70902c51",
          5175 => x"5a7980c1",
          5176 => x"2e89d438",
          5177 => x"7980c124",
          5178 => x"80d93879",
          5179 => x"ab2e83b9",
          5180 => x"3879ab24",
          5181 => x"a4387982",
          5182 => x"2e81b338",
          5183 => x"7982248a",
          5184 => x"3879802e",
          5185 => x"ffaf388e",
          5186 => x"ed397984",
          5187 => x"2e828338",
          5188 => x"79942e82",
          5189 => x"ad388ede",
          5190 => x"3979bd2e",
          5191 => x"84ff3879",
          5192 => x"bd249038",
          5193 => x"79b02e83",
          5194 => x"a63879bc",
          5195 => x"2e848838",
          5196 => x"8ec43979",
          5197 => x"bf2e85c6",
          5198 => x"387980c0",
          5199 => x"2e86bd38",
          5200 => x"8eb43979",
          5201 => x"80d52e8d",
          5202 => x"90387980",
          5203 => x"d524b038",
          5204 => x"7980d02e",
          5205 => x"8cc93879",
          5206 => x"80d02492",
          5207 => x"387980c2",
          5208 => x"2e89f638",
          5209 => x"7980c32e",
          5210 => x"8b9b388e",
          5211 => x"89397980",
          5212 => x"d12e8cba",
          5213 => x"387980d4",
          5214 => x"2e8cc238",
          5215 => x"8df83979",
          5216 => x"81822e8d",
          5217 => x"d1387981",
          5218 => x"82249238",
          5219 => x"7980f82e",
          5220 => x"8ce33879",
          5221 => x"80f92e8d",
          5222 => x"80388dda",
          5223 => x"39798183",
          5224 => x"2e8dc138",
          5225 => x"7981852e",
          5226 => x"8dc6388d",
          5227 => x"c939b53d",
          5228 => x"ff801153",
          5229 => x"ff840551",
          5230 => x"d1f83f82",
          5231 => x"bb980888",
          5232 => x"3882a6a8",
          5233 => x"518fb139",
          5234 => x"b53dfefc",
          5235 => x"1153ff84",
          5236 => x"0551d1de",
          5237 => x"3f82bb98",
          5238 => x"08802e88",
          5239 => x"38816425",
          5240 => x"83388044",
          5241 => x"0280cf05",
          5242 => x"33520280",
          5243 => x"d3053351",
          5244 => x"80c7ec3f",
          5245 => x"82bb9808",
          5246 => x"81ff065a",
          5247 => x"798d3882",
          5248 => x"a6b851d6",
          5249 => x"fe3f815f",
          5250 => x"fdab3982",
          5251 => x"a6c8518e",
          5252 => x"e739b53d",
          5253 => x"ff801153",
          5254 => x"ff840551",
          5255 => x"d1943f82",
          5256 => x"bb980880",
          5257 => x"2efd8e38",
          5258 => x"80538052",
          5259 => x"0280d305",
          5260 => x"335180cb",
          5261 => x"f73f82bb",
          5262 => x"98085282",
          5263 => x"a6e0518c",
          5264 => x"8e39b53d",
          5265 => x"ff801153",
          5266 => x"ff840551",
          5267 => x"d0e43f82",
          5268 => x"bb980880",
          5269 => x"2e873864",
          5270 => x"8926fcd9",
          5271 => x"38b53dfe",
          5272 => x"fc1153ff",
          5273 => x"840551d0",
          5274 => x"c93f82bb",
          5275 => x"98088638",
          5276 => x"82bb9808",
          5277 => x"44645382",
          5278 => x"a6e8527a",
          5279 => x"51ffb1be",
          5280 => x"3f0280cf",
          5281 => x"0533537a",
          5282 => x"526484b4",
          5283 => x"2982bcc4",
          5284 => x"055180f6",
          5285 => x"8e3f82bb",
          5286 => x"98088190",
          5287 => x"3882a6b8",
          5288 => x"51d5e03f",
          5289 => x"815efc8d",
          5290 => x"39b53dff",
          5291 => x"8405518f",
          5292 => x"b13f82bb",
          5293 => x"9808b63d",
          5294 => x"ff840552",
          5295 => x"5c90c73f",
          5296 => x"815382bb",
          5297 => x"9808527b",
          5298 => x"51f2ab3f",
          5299 => x"80d539b5",
          5300 => x"3dff8405",
          5301 => x"518f8b3f",
          5302 => x"82bb9808",
          5303 => x"b63dff84",
          5304 => x"05525c90",
          5305 => x"a13f82bb",
          5306 => x"9808b63d",
          5307 => x"ff840552",
          5308 => x"5b90933f",
          5309 => x"82bb9808",
          5310 => x"b63dff84",
          5311 => x"05525a90",
          5312 => x"853f82d2",
          5313 => x"e85982b9",
          5314 => x"bc5882bb",
          5315 => x"c8578056",
          5316 => x"805582bb",
          5317 => x"980881ff",
          5318 => x"06547953",
          5319 => x"7a527b51",
          5320 => x"f3913f82",
          5321 => x"bb980880",
          5322 => x"2efb8a38",
          5323 => x"82bb9808",
          5324 => x"51efe33f",
          5325 => x"faff39b5",
          5326 => x"3dff8011",
          5327 => x"53ff8405",
          5328 => x"51ceef3f",
          5329 => x"82bb9808",
          5330 => x"802efae9",
          5331 => x"38b53dfe",
          5332 => x"fc1153ff",
          5333 => x"840551ce",
          5334 => x"d93f82bb",
          5335 => x"9808802e",
          5336 => x"fad338b5",
          5337 => x"3dfef811",
          5338 => x"53ff8405",
          5339 => x"51cec33f",
          5340 => x"82bb9808",
          5341 => x"863882bb",
          5342 => x"98084382",
          5343 => x"a6ec51d4",
          5344 => x"823f6464",
          5345 => x"5d5b7a7c",
          5346 => x"2781ea38",
          5347 => x"625a797b",
          5348 => x"7084055d",
          5349 => x"0c7b7b26",
          5350 => x"f53881d9",
          5351 => x"39b53dff",
          5352 => x"801153ff",
          5353 => x"840551ce",
          5354 => x"893f82bb",
          5355 => x"9808802e",
          5356 => x"fa8338b5",
          5357 => x"3dfefc11",
          5358 => x"53ff8405",
          5359 => x"51cdf33f",
          5360 => x"82bb9808",
          5361 => x"802ef9ed",
          5362 => x"38b53dfe",
          5363 => x"f81153ff",
          5364 => x"840551cd",
          5365 => x"dd3f82bb",
          5366 => x"9808802e",
          5367 => x"f9d73882",
          5368 => x"a6fc51d3",
          5369 => x"9e3f645b",
          5370 => x"7a642781",
          5371 => x"8838625a",
          5372 => x"7a708105",
          5373 => x"5c337a34",
          5374 => x"62810543",
          5375 => x"eb39b53d",
          5376 => x"ff801153",
          5377 => x"ff840551",
          5378 => x"cda83f82",
          5379 => x"bb980880",
          5380 => x"2ef9a238",
          5381 => x"b53dfefc",
          5382 => x"1153ff84",
          5383 => x"0551cd92",
          5384 => x"3f82bb98",
          5385 => x"08802ef9",
          5386 => x"8c38b53d",
          5387 => x"fef81153",
          5388 => x"ff840551",
          5389 => x"ccfc3f82",
          5390 => x"bb980880",
          5391 => x"2ef8f638",
          5392 => x"82a78851",
          5393 => x"d2bd3f64",
          5394 => x"5b7a6427",
          5395 => x"a8386270",
          5396 => x"337c335f",
          5397 => x"5b5c797d",
          5398 => x"2e923879",
          5399 => x"557b547a",
          5400 => x"33537a52",
          5401 => x"82a79851",
          5402 => x"ffaaeb3f",
          5403 => x"811b6381",
          5404 => x"05445bd5",
          5405 => x"3982a7b0",
          5406 => x"5189fd39",
          5407 => x"b53dff80",
          5408 => x"1153ff84",
          5409 => x"0551ccaa",
          5410 => x"3f82bb98",
          5411 => x"0880df38",
          5412 => x"82ba8433",
          5413 => x"5a79802e",
          5414 => x"893882b9",
          5415 => x"bc084580",
          5416 => x"cd3982ba",
          5417 => x"85335a79",
          5418 => x"802e8838",
          5419 => x"82b9c408",
          5420 => x"45bc3982",
          5421 => x"ba86335a",
          5422 => x"79802e88",
          5423 => x"3882b9cc",
          5424 => x"0845ab39",
          5425 => x"82ba8733",
          5426 => x"5a79802e",
          5427 => x"883882b9",
          5428 => x"d408459a",
          5429 => x"3982ba82",
          5430 => x"335a7980",
          5431 => x"2e883882",
          5432 => x"b9dc0845",
          5433 => x"893982b9",
          5434 => x"ec08fc80",
          5435 => x"0545b53d",
          5436 => x"fefc1153",
          5437 => x"ff840551",
          5438 => x"cbb83f82",
          5439 => x"bb980880",
          5440 => x"de3882ba",
          5441 => x"84335a79",
          5442 => x"802e8938",
          5443 => x"82b9c008",
          5444 => x"4480cc39",
          5445 => x"82ba8533",
          5446 => x"5a79802e",
          5447 => x"883882b9",
          5448 => x"c80844bb",
          5449 => x"3982ba86",
          5450 => x"335a7980",
          5451 => x"2e883882",
          5452 => x"b9d00844",
          5453 => x"aa3982ba",
          5454 => x"87335a79",
          5455 => x"802e8838",
          5456 => x"82b9d808",
          5457 => x"44993982",
          5458 => x"ba82335a",
          5459 => x"79802e88",
          5460 => x"3882b9e0",
          5461 => x"08448839",
          5462 => x"82b9ec08",
          5463 => x"880544b5",
          5464 => x"3dfef811",
          5465 => x"53ff8405",
          5466 => x"51cac73f",
          5467 => x"82bb9808",
          5468 => x"802ea738",
          5469 => x"80635d5d",
          5470 => x"7b882e83",
          5471 => x"38815d7b",
          5472 => x"90327030",
          5473 => x"7072079f",
          5474 => x"2a706006",
          5475 => x"51515b5b",
          5476 => x"79802e88",
          5477 => x"387ba02e",
          5478 => x"83388843",
          5479 => x"82a7b451",
          5480 => x"cfe13fa0",
          5481 => x"55645462",
          5482 => x"53635264",
          5483 => x"51eecf3f",
          5484 => x"82a7c451",
          5485 => x"87c239b5",
          5486 => x"3dff8011",
          5487 => x"53ff8405",
          5488 => x"51c9ef3f",
          5489 => x"82bb9808",
          5490 => x"802ef5e9",
          5491 => x"38b53dfe",
          5492 => x"fc1153ff",
          5493 => x"840551c9",
          5494 => x"d93f82bb",
          5495 => x"9808802e",
          5496 => x"a438645a",
          5497 => x"0280cf05",
          5498 => x"337a3464",
          5499 => x"810545b5",
          5500 => x"3dfefc11",
          5501 => x"53ff8405",
          5502 => x"51c9b73f",
          5503 => x"82bb9808",
          5504 => x"e138f5b1",
          5505 => x"39647033",
          5506 => x"545282a7",
          5507 => x"d051ffa7",
          5508 => x"c53f80f8",
          5509 => x"527a51c8",
          5510 => x"e33f7a46",
          5511 => x"7a335a79",
          5512 => x"ae2ef591",
          5513 => x"389f7a27",
          5514 => x"9f38b53d",
          5515 => x"fefc1153",
          5516 => x"ff840551",
          5517 => x"c8fc3f82",
          5518 => x"bb980880",
          5519 => x"2e913864",
          5520 => x"5a0280cf",
          5521 => x"05337a34",
          5522 => x"64810545",
          5523 => x"ffb73982",
          5524 => x"a7dc51ce",
          5525 => x"ae3fffad",
          5526 => x"39b53dfe",
          5527 => x"f41153ff",
          5528 => x"840551c2",
          5529 => x"c63f82bb",
          5530 => x"9808802e",
          5531 => x"f4c738b5",
          5532 => x"3dfef011",
          5533 => x"53ff8405",
          5534 => x"51c2b03f",
          5535 => x"82bb9808",
          5536 => x"802ea638",
          5537 => x"615a0280",
          5538 => x"c205227a",
          5539 => x"7082055c",
          5540 => x"237942b5",
          5541 => x"3dfef011",
          5542 => x"53ff8405",
          5543 => x"51c28c3f",
          5544 => x"82bb9808",
          5545 => x"df38f48d",
          5546 => x"39617022",
          5547 => x"545282a7",
          5548 => x"e451ffa6",
          5549 => x"a13f80f8",
          5550 => x"527a51c7",
          5551 => x"bf3f7a46",
          5552 => x"7a335a79",
          5553 => x"ae2ef3ed",
          5554 => x"38799f26",
          5555 => x"87386182",
          5556 => x"0542d639",
          5557 => x"b53dfef0",
          5558 => x"1153ff84",
          5559 => x"0551c1cb",
          5560 => x"3f82bb98",
          5561 => x"08802e93",
          5562 => x"38615a02",
          5563 => x"80c20522",
          5564 => x"7a708205",
          5565 => x"5c237942",
          5566 => x"ffaf3982",
          5567 => x"a7dc51cd",
          5568 => x"823fffa5",
          5569 => x"39b53dfe",
          5570 => x"f41153ff",
          5571 => x"840551c1",
          5572 => x"9a3f82bb",
          5573 => x"9808802e",
          5574 => x"f39b38b5",
          5575 => x"3dfef011",
          5576 => x"53ff8405",
          5577 => x"51c1843f",
          5578 => x"82bb9808",
          5579 => x"802ea038",
          5580 => x"6161710c",
          5581 => x"5a618405",
          5582 => x"42b53dfe",
          5583 => x"f01153ff",
          5584 => x"840551c0",
          5585 => x"e63f82bb",
          5586 => x"9808e538",
          5587 => x"f2e73961",
          5588 => x"70085452",
          5589 => x"82a7f051",
          5590 => x"ffa4fb3f",
          5591 => x"80f8527a",
          5592 => x"51c6993f",
          5593 => x"7a467a33",
          5594 => x"5a79ae2e",
          5595 => x"f2c7389f",
          5596 => x"7a279b38",
          5597 => x"b53dfef0",
          5598 => x"1153ff84",
          5599 => x"0551c0ab",
          5600 => x"3f82bb98",
          5601 => x"08802e8d",
          5602 => x"38616171",
          5603 => x"0c5a6184",
          5604 => x"0542ffbb",
          5605 => x"3982a7dc",
          5606 => x"51cbe83f",
          5607 => x"ffb13982",
          5608 => x"a7fc51cb",
          5609 => x"de3f8251",
          5610 => x"988b3ff2",
          5611 => x"883982a8",
          5612 => x"9451cbcf",
          5613 => x"3fa25197",
          5614 => x"e03ff1f9",
          5615 => x"3982a8ac",
          5616 => x"51cbc03f",
          5617 => x"8480810b",
          5618 => x"87c09484",
          5619 => x"0c848081",
          5620 => x"0b87c094",
          5621 => x"940cf1dd",
          5622 => x"3982a8c0",
          5623 => x"51cba43f",
          5624 => x"8c80830b",
          5625 => x"87c09484",
          5626 => x"0c8c8083",
          5627 => x"0b87c094",
          5628 => x"940cf1c1",
          5629 => x"39b53dff",
          5630 => x"801153ff",
          5631 => x"840551c5",
          5632 => x"b13f82bb",
          5633 => x"9808802e",
          5634 => x"f1ab3864",
          5635 => x"5282a8d4",
          5636 => x"51ffa3c2",
          5637 => x"3f645a79",
          5638 => x"04b53dff",
          5639 => x"801153ff",
          5640 => x"840551c5",
          5641 => x"8d3f82bb",
          5642 => x"9808802e",
          5643 => x"f1873864",
          5644 => x"5282a8f0",
          5645 => x"51ffa39e",
          5646 => x"3f645a79",
          5647 => x"2d82bb98",
          5648 => x"08802ef0",
          5649 => x"f03882bb",
          5650 => x"98085282",
          5651 => x"a98c51ff",
          5652 => x"a3843ff0",
          5653 => x"e03982a9",
          5654 => x"a851caa7",
          5655 => x"3fffa2d7",
          5656 => x"3ff0d239",
          5657 => x"82a9c451",
          5658 => x"ca993f80",
          5659 => x"5affa839",
          5660 => x"91ad3ff0",
          5661 => x"c0397a46",
          5662 => x"7a335a79",
          5663 => x"802ef0b5",
          5664 => x"387e7e06",
          5665 => x"5a79802e",
          5666 => x"81d638b5",
          5667 => x"3dff8405",
          5668 => x"5183cf3f",
          5669 => x"82bb9808",
          5670 => x"5c815d7c",
          5671 => x"822eb238",
          5672 => x"7c822489",
          5673 => x"387c812e",
          5674 => x"8c3880cd",
          5675 => x"397c832e",
          5676 => x"b03880c5",
          5677 => x"3982a9d8",
          5678 => x"567b5582",
          5679 => x"a9dc5480",
          5680 => x"5382a9e0",
          5681 => x"52b53dff",
          5682 => x"b00551ff",
          5683 => x"a4f03fbb",
          5684 => x"3982aa80",
          5685 => x"52b53dff",
          5686 => x"b00551ff",
          5687 => x"a4e03fab",
          5688 => x"397b5582",
          5689 => x"a9dc5480",
          5690 => x"5382a9f0",
          5691 => x"52b53dff",
          5692 => x"b00551ff",
          5693 => x"a4c83f93",
          5694 => x"397b5480",
          5695 => x"5382a9fc",
          5696 => x"52b53dff",
          5697 => x"b00551ff",
          5698 => x"a4b43f82",
          5699 => x"d2e85982",
          5700 => x"b9bc5882",
          5701 => x"bbc85780",
          5702 => x"56655580",
          5703 => x"5482e080",
          5704 => x"5382e080",
          5705 => x"52b53dff",
          5706 => x"b00551e7",
          5707 => x"863f82bb",
          5708 => x"980882bb",
          5709 => x"98080970",
          5710 => x"30707207",
          5711 => x"8025515c",
          5712 => x"5c40805b",
          5713 => x"7c832683",
          5714 => x"38815b79",
          5715 => x"7b065a79",
          5716 => x"802e8d38",
          5717 => x"811d7081",
          5718 => x"ff065e5a",
          5719 => x"7cfebc38",
          5720 => x"7e81327e",
          5721 => x"8132075a",
          5722 => x"798a387f",
          5723 => x"ff2e0981",
          5724 => x"06eec238",
          5725 => x"82aa8451",
          5726 => x"c8893fee",
          5727 => x"b839f53d",
          5728 => x"0d800b82",
          5729 => x"bbc83487",
          5730 => x"c0948c70",
          5731 => x"08545587",
          5732 => x"84805272",
          5733 => x"51df8c3f",
          5734 => x"82bb9808",
          5735 => x"902b7508",
          5736 => x"55538784",
          5737 => x"80527351",
          5738 => x"def93f72",
          5739 => x"82bb9808",
          5740 => x"07750c87",
          5741 => x"c0949c70",
          5742 => x"08545587",
          5743 => x"84805272",
          5744 => x"51dee03f",
          5745 => x"82bb9808",
          5746 => x"902b7508",
          5747 => x"55538784",
          5748 => x"80527351",
          5749 => x"decd3f72",
          5750 => x"82bb9808",
          5751 => x"07750c8c",
          5752 => x"80830b87",
          5753 => x"c094840c",
          5754 => x"8c80830b",
          5755 => x"87c09494",
          5756 => x"0c80fa82",
          5757 => x"5a80fcee",
          5758 => x"5b830284",
          5759 => x"05990534",
          5760 => x"805c82d2",
          5761 => x"e80b873d",
          5762 => x"7088130c",
          5763 => x"70720c82",
          5764 => x"d2ec0c54",
          5765 => x"89bd3f93",
          5766 => x"c13f82aa",
          5767 => x"9451c6e3",
          5768 => x"3f82aaa0",
          5769 => x"51c6dc3f",
          5770 => x"80dda851",
          5771 => x"92e63f81",
          5772 => x"51e8b83f",
          5773 => x"ecae3f80",
          5774 => x"04fe3d0d",
          5775 => x"80528353",
          5776 => x"71882b52",
          5777 => x"87d93f82",
          5778 => x"bb980881",
          5779 => x"ff067207",
          5780 => x"ff145452",
          5781 => x"728025e8",
          5782 => x"387182bb",
          5783 => x"980c843d",
          5784 => x"0d04fc3d",
          5785 => x"0d767008",
          5786 => x"54558073",
          5787 => x"52547274",
          5788 => x"2e818a38",
          5789 => x"72335170",
          5790 => x"a02e0981",
          5791 => x"06863881",
          5792 => x"1353f139",
          5793 => x"72335170",
          5794 => x"a22e0981",
          5795 => x"06863881",
          5796 => x"13538154",
          5797 => x"72527381",
          5798 => x"2e098106",
          5799 => x"9f388439",
          5800 => x"81125280",
          5801 => x"72335254",
          5802 => x"70a22e83",
          5803 => x"38815470",
          5804 => x"802e9d38",
          5805 => x"73ea3898",
          5806 => x"39811252",
          5807 => x"80723352",
          5808 => x"5470a02e",
          5809 => x"83388154",
          5810 => x"70802e84",
          5811 => x"3873ea38",
          5812 => x"80723352",
          5813 => x"5470a02e",
          5814 => x"09810683",
          5815 => x"38815470",
          5816 => x"a2327030",
          5817 => x"70802576",
          5818 => x"07515151",
          5819 => x"70802e88",
          5820 => x"38807270",
          5821 => x"81055434",
          5822 => x"71750c72",
          5823 => x"517082bb",
          5824 => x"980c863d",
          5825 => x"0d04fc3d",
          5826 => x"0d765372",
          5827 => x"08802e92",
          5828 => x"38863dfc",
          5829 => x"05527251",
          5830 => x"ffb9903f",
          5831 => x"82bb9808",
          5832 => x"85388053",
          5833 => x"83397453",
          5834 => x"7282bb98",
          5835 => x"0c863d0d",
          5836 => x"04fc3d0d",
          5837 => x"76821133",
          5838 => x"ff055253",
          5839 => x"8152708b",
          5840 => x"26819838",
          5841 => x"831333ff",
          5842 => x"05518252",
          5843 => x"709e2681",
          5844 => x"8a388413",
          5845 => x"33518352",
          5846 => x"70972680",
          5847 => x"fe388513",
          5848 => x"33518452",
          5849 => x"70bb2680",
          5850 => x"f2388613",
          5851 => x"33518552",
          5852 => x"70bb2680",
          5853 => x"e6388813",
          5854 => x"22558652",
          5855 => x"7487e726",
          5856 => x"80d9388a",
          5857 => x"13225487",
          5858 => x"527387e7",
          5859 => x"2680cc38",
          5860 => x"810b87c0",
          5861 => x"989c0c72",
          5862 => x"2287c098",
          5863 => x"bc0c8213",
          5864 => x"3387c098",
          5865 => x"b80c8313",
          5866 => x"3387c098",
          5867 => x"b40c8413",
          5868 => x"3387c098",
          5869 => x"b00c8513",
          5870 => x"3387c098",
          5871 => x"ac0c8613",
          5872 => x"3387c098",
          5873 => x"a80c7487",
          5874 => x"c098a40c",
          5875 => x"7387c098",
          5876 => x"a00c800b",
          5877 => x"87c0989c",
          5878 => x"0c805271",
          5879 => x"82bb980c",
          5880 => x"863d0d04",
          5881 => x"f33d0d7f",
          5882 => x"5b87c098",
          5883 => x"9c5d817d",
          5884 => x"0c87c098",
          5885 => x"bc085e7d",
          5886 => x"7b2387c0",
          5887 => x"98b8085a",
          5888 => x"79821c34",
          5889 => x"87c098b4",
          5890 => x"085a7983",
          5891 => x"1c3487c0",
          5892 => x"98b0085a",
          5893 => x"79841c34",
          5894 => x"87c098ac",
          5895 => x"085a7985",
          5896 => x"1c3487c0",
          5897 => x"98a8085a",
          5898 => x"79861c34",
          5899 => x"87c098a4",
          5900 => x"085c7b88",
          5901 => x"1c2387c0",
          5902 => x"98a0085a",
          5903 => x"798a1c23",
          5904 => x"807d0c79",
          5905 => x"83ffff06",
          5906 => x"597b83ff",
          5907 => x"ff065886",
          5908 => x"1b335785",
          5909 => x"1b335684",
          5910 => x"1b335583",
          5911 => x"1b335482",
          5912 => x"1b33537d",
          5913 => x"83ffff06",
          5914 => x"5282aab8",
          5915 => x"51ff9ae6",
          5916 => x"3f8f3d0d",
          5917 => x"04fb3d0d",
          5918 => x"029f0533",
          5919 => x"82b9b833",
          5920 => x"7081ff06",
          5921 => x"58555587",
          5922 => x"c0948451",
          5923 => x"75802e86",
          5924 => x"3887c094",
          5925 => x"94517008",
          5926 => x"70962a70",
          5927 => x"81065354",
          5928 => x"5270802e",
          5929 => x"8c387191",
          5930 => x"2a708106",
          5931 => x"515170d7",
          5932 => x"38728132",
          5933 => x"70810651",
          5934 => x"5170802e",
          5935 => x"8d387193",
          5936 => x"2a708106",
          5937 => x"515170ff",
          5938 => x"be387381",
          5939 => x"ff065187",
          5940 => x"c0948052",
          5941 => x"70802e86",
          5942 => x"3887c094",
          5943 => x"90527472",
          5944 => x"0c7482bb",
          5945 => x"980c873d",
          5946 => x"0d04ff3d",
          5947 => x"0d028f05",
          5948 => x"33703070",
          5949 => x"9f2a5152",
          5950 => x"527082b9",
          5951 => x"b834833d",
          5952 => x"0d04f93d",
          5953 => x"0d02a705",
          5954 => x"3358778a",
          5955 => x"2e098106",
          5956 => x"87387a52",
          5957 => x"8d51eb3f",
          5958 => x"82b9b833",
          5959 => x"7081ff06",
          5960 => x"585687c0",
          5961 => x"94845376",
          5962 => x"802e8638",
          5963 => x"87c09494",
          5964 => x"53720870",
          5965 => x"962a7081",
          5966 => x"06555654",
          5967 => x"72802e8c",
          5968 => x"3873912a",
          5969 => x"70810651",
          5970 => x"5372d738",
          5971 => x"74813270",
          5972 => x"81065153",
          5973 => x"72802e8d",
          5974 => x"3873932a",
          5975 => x"70810651",
          5976 => x"5372ffbe",
          5977 => x"387581ff",
          5978 => x"065387c0",
          5979 => x"94805472",
          5980 => x"802e8638",
          5981 => x"87c09490",
          5982 => x"5477740c",
          5983 => x"800b82bb",
          5984 => x"980c893d",
          5985 => x"0d04f93d",
          5986 => x"0d795480",
          5987 => x"74337081",
          5988 => x"ff065353",
          5989 => x"5770772e",
          5990 => x"80fc3871",
          5991 => x"81ff0681",
          5992 => x"1582b9b8",
          5993 => x"337081ff",
          5994 => x"06595755",
          5995 => x"5887c094",
          5996 => x"84517580",
          5997 => x"2e863887",
          5998 => x"c0949451",
          5999 => x"70087096",
          6000 => x"2a708106",
          6001 => x"53545270",
          6002 => x"802e8c38",
          6003 => x"71912a70",
          6004 => x"81065151",
          6005 => x"70d73872",
          6006 => x"81327081",
          6007 => x"06515170",
          6008 => x"802e8d38",
          6009 => x"71932a70",
          6010 => x"81065151",
          6011 => x"70ffbe38",
          6012 => x"7481ff06",
          6013 => x"5187c094",
          6014 => x"80527080",
          6015 => x"2e863887",
          6016 => x"c0949052",
          6017 => x"77720c81",
          6018 => x"17743370",
          6019 => x"81ff0653",
          6020 => x"535770ff",
          6021 => x"86387682",
          6022 => x"bb980c89",
          6023 => x"3d0d04fe",
          6024 => x"3d0d82b9",
          6025 => x"b8337081",
          6026 => x"ff065452",
          6027 => x"87c09484",
          6028 => x"5172802e",
          6029 => x"863887c0",
          6030 => x"94945170",
          6031 => x"0870822a",
          6032 => x"70810651",
          6033 => x"51517080",
          6034 => x"2ee23871",
          6035 => x"81ff0651",
          6036 => x"87c09480",
          6037 => x"5270802e",
          6038 => x"863887c0",
          6039 => x"94905271",
          6040 => x"087081ff",
          6041 => x"0682bb98",
          6042 => x"0c51843d",
          6043 => x"0d04ffaf",
          6044 => x"3f82bb98",
          6045 => x"0881ff06",
          6046 => x"82bb980c",
          6047 => x"04fe3d0d",
          6048 => x"82b9b833",
          6049 => x"7081ff06",
          6050 => x"525387c0",
          6051 => x"94845270",
          6052 => x"802e8638",
          6053 => x"87c09494",
          6054 => x"52710870",
          6055 => x"822a7081",
          6056 => x"06515151",
          6057 => x"ff527080",
          6058 => x"2ea03872",
          6059 => x"81ff0651",
          6060 => x"87c09480",
          6061 => x"5270802e",
          6062 => x"863887c0",
          6063 => x"94905271",
          6064 => x"0870982b",
          6065 => x"70982c51",
          6066 => x"53517182",
          6067 => x"bb980c84",
          6068 => x"3d0d04ff",
          6069 => x"3d0d87c0",
          6070 => x"9e800870",
          6071 => x"9c2a8a06",
          6072 => x"51517080",
          6073 => x"2e84b438",
          6074 => x"87c09ea4",
          6075 => x"0882b9bc",
          6076 => x"0c87c09e",
          6077 => x"a80882b9",
          6078 => x"c00c87c0",
          6079 => x"9e940882",
          6080 => x"b9c40c87",
          6081 => x"c09e9808",
          6082 => x"82b9c80c",
          6083 => x"87c09e9c",
          6084 => x"0882b9cc",
          6085 => x"0c87c09e",
          6086 => x"a00882b9",
          6087 => x"d00c87c0",
          6088 => x"9eac0882",
          6089 => x"b9d40c87",
          6090 => x"c09eb008",
          6091 => x"82b9d80c",
          6092 => x"87c09eb4",
          6093 => x"0882b9dc",
          6094 => x"0c87c09e",
          6095 => x"b80882b9",
          6096 => x"e00c87c0",
          6097 => x"9ebc0882",
          6098 => x"b9e40c87",
          6099 => x"c09ec008",
          6100 => x"82b9e80c",
          6101 => x"87c09ec4",
          6102 => x"0882b9ec",
          6103 => x"0c87c09e",
          6104 => x"80085170",
          6105 => x"82b9f023",
          6106 => x"87c09e84",
          6107 => x"0882b9f4",
          6108 => x"0c87c09e",
          6109 => x"880882b9",
          6110 => x"f80c87c0",
          6111 => x"9e8c0882",
          6112 => x"b9fc0c81",
          6113 => x"0b82ba80",
          6114 => x"34800b87",
          6115 => x"c09e9008",
          6116 => x"7084800a",
          6117 => x"06515252",
          6118 => x"70802e83",
          6119 => x"38815271",
          6120 => x"82ba8134",
          6121 => x"800b87c0",
          6122 => x"9e900870",
          6123 => x"88800a06",
          6124 => x"51525270",
          6125 => x"802e8338",
          6126 => x"81527182",
          6127 => x"ba823480",
          6128 => x"0b87c09e",
          6129 => x"90087090",
          6130 => x"800a0651",
          6131 => x"52527080",
          6132 => x"2e833881",
          6133 => x"527182ba",
          6134 => x"8334800b",
          6135 => x"87c09e90",
          6136 => x"08708880",
          6137 => x"80065152",
          6138 => x"5270802e",
          6139 => x"83388152",
          6140 => x"7182ba84",
          6141 => x"34800b87",
          6142 => x"c09e9008",
          6143 => x"70a08080",
          6144 => x"06515252",
          6145 => x"70802e83",
          6146 => x"38815271",
          6147 => x"82ba8534",
          6148 => x"800b87c0",
          6149 => x"9e900870",
          6150 => x"90808006",
          6151 => x"51525270",
          6152 => x"802e8338",
          6153 => x"81527182",
          6154 => x"ba863480",
          6155 => x"0b87c09e",
          6156 => x"90087084",
          6157 => x"80800651",
          6158 => x"52527080",
          6159 => x"2e833881",
          6160 => x"527182ba",
          6161 => x"8734800b",
          6162 => x"87c09e90",
          6163 => x"08708280",
          6164 => x"80065152",
          6165 => x"5270802e",
          6166 => x"83388152",
          6167 => x"7182ba88",
          6168 => x"34800b87",
          6169 => x"c09e9008",
          6170 => x"70818080",
          6171 => x"06515252",
          6172 => x"70802e83",
          6173 => x"38815271",
          6174 => x"82ba8934",
          6175 => x"800b87c0",
          6176 => x"9e900870",
          6177 => x"80c08006",
          6178 => x"51525270",
          6179 => x"802e8338",
          6180 => x"81527182",
          6181 => x"ba8a3480",
          6182 => x"0b87c09e",
          6183 => x"900870a0",
          6184 => x"80065152",
          6185 => x"5270802e",
          6186 => x"83388152",
          6187 => x"7182ba8b",
          6188 => x"3487c09e",
          6189 => x"90087098",
          6190 => x"8006708a",
          6191 => x"2a515151",
          6192 => x"7082ba8c",
          6193 => x"34800b87",
          6194 => x"c09e9008",
          6195 => x"70848006",
          6196 => x"51525270",
          6197 => x"802e8338",
          6198 => x"81527182",
          6199 => x"ba8d3487",
          6200 => x"c09e9008",
          6201 => x"7083f006",
          6202 => x"70842a51",
          6203 => x"51517082",
          6204 => x"ba8e3480",
          6205 => x"0b87c09e",
          6206 => x"90087088",
          6207 => x"06515252",
          6208 => x"70802e83",
          6209 => x"38815271",
          6210 => x"82ba8f34",
          6211 => x"87c09e90",
          6212 => x"08708706",
          6213 => x"51517082",
          6214 => x"ba903483",
          6215 => x"3d0d04fb",
          6216 => x"3d0d82aa",
          6217 => x"d051ffb8",
          6218 => x"da3f82ba",
          6219 => x"80335473",
          6220 => x"802e8938",
          6221 => x"82aae451",
          6222 => x"ffb8c83f",
          6223 => x"82aaf851",
          6224 => x"ffb8c03f",
          6225 => x"82ba8233",
          6226 => x"5473802e",
          6227 => x"943882b9",
          6228 => x"dc0882b9",
          6229 => x"e0081154",
          6230 => x"5282ab90",
          6231 => x"51ff90f6",
          6232 => x"3f82ba87",
          6233 => x"33547380",
          6234 => x"2e943882",
          6235 => x"b9d40882",
          6236 => x"b9d80811",
          6237 => x"545282ab",
          6238 => x"ac51ff90",
          6239 => x"d93f82ba",
          6240 => x"84335473",
          6241 => x"802e9438",
          6242 => x"82b9bc08",
          6243 => x"82b9c008",
          6244 => x"11545282",
          6245 => x"abc851ff",
          6246 => x"90bc3f82",
          6247 => x"ba853354",
          6248 => x"73802e94",
          6249 => x"3882b9c4",
          6250 => x"0882b9c8",
          6251 => x"08115452",
          6252 => x"82abe451",
          6253 => x"ff909f3f",
          6254 => x"82ba8633",
          6255 => x"5473802e",
          6256 => x"943882b9",
          6257 => x"cc0882b9",
          6258 => x"d0081154",
          6259 => x"5282ac80",
          6260 => x"51ff9082",
          6261 => x"3f82ba8b",
          6262 => x"33547380",
          6263 => x"2e8e3882",
          6264 => x"ba8c3352",
          6265 => x"82ac9c51",
          6266 => x"ff8feb3f",
          6267 => x"82ba8f33",
          6268 => x"5473802e",
          6269 => x"8e3882ba",
          6270 => x"90335282",
          6271 => x"acbc51ff",
          6272 => x"8fd43f82",
          6273 => x"ba8d3354",
          6274 => x"73802e8e",
          6275 => x"3882ba8e",
          6276 => x"335282ac",
          6277 => x"dc51ff8f",
          6278 => x"bd3f82ba",
          6279 => x"81335473",
          6280 => x"802e8938",
          6281 => x"82acfc51",
          6282 => x"ffb6d83f",
          6283 => x"82ba8333",
          6284 => x"5473802e",
          6285 => x"893882ad",
          6286 => x"9051ffb6",
          6287 => x"c63f82ba",
          6288 => x"88335473",
          6289 => x"802e8938",
          6290 => x"82ad9c51",
          6291 => x"ffb6b43f",
          6292 => x"82ba8933",
          6293 => x"5473802e",
          6294 => x"893882ad",
          6295 => x"a851ffb6",
          6296 => x"a23f82ba",
          6297 => x"8a335473",
          6298 => x"802e8938",
          6299 => x"82adb451",
          6300 => x"ffb6903f",
          6301 => x"82adc051",
          6302 => x"ffb6883f",
          6303 => x"82b9e408",
          6304 => x"5282adcc",
          6305 => x"51ff8ece",
          6306 => x"3f82b9e8",
          6307 => x"085282ad",
          6308 => x"f451ff8e",
          6309 => x"c13f82b9",
          6310 => x"ec085282",
          6311 => x"ae9c51ff",
          6312 => x"8eb43f82",
          6313 => x"aec451ff",
          6314 => x"b5d93f82",
          6315 => x"b9f02252",
          6316 => x"82aecc51",
          6317 => x"ff8e9f3f",
          6318 => x"82b9f408",
          6319 => x"56bd84c0",
          6320 => x"527551cc",
          6321 => x"de3f82bb",
          6322 => x"9808bd84",
          6323 => x"c0297671",
          6324 => x"31545482",
          6325 => x"bb980852",
          6326 => x"82aef451",
          6327 => x"ff8df73f",
          6328 => x"82ba8733",
          6329 => x"5473802e",
          6330 => x"a93882b9",
          6331 => x"f80856bd",
          6332 => x"84c05275",
          6333 => x"51ccac3f",
          6334 => x"82bb9808",
          6335 => x"bd84c029",
          6336 => x"76713154",
          6337 => x"5482bb98",
          6338 => x"085282af",
          6339 => x"a051ff8d",
          6340 => x"c53f82ba",
          6341 => x"82335473",
          6342 => x"802ea938",
          6343 => x"82b9fc08",
          6344 => x"56bd84c0",
          6345 => x"527551cb",
          6346 => x"fa3f82bb",
          6347 => x"9808bd84",
          6348 => x"c0297671",
          6349 => x"31545482",
          6350 => x"bb980852",
          6351 => x"82afcc51",
          6352 => x"ff8d933f",
          6353 => x"82a7b051",
          6354 => x"ffb4b83f",
          6355 => x"873d0d04",
          6356 => x"fe3d0d02",
          6357 => x"920533ff",
          6358 => x"05527184",
          6359 => x"26aa3871",
          6360 => x"8429829a",
          6361 => x"80055271",
          6362 => x"080482af",
          6363 => x"f8519d39",
          6364 => x"82b08051",
          6365 => x"973982b0",
          6366 => x"88519139",
          6367 => x"82b09051",
          6368 => x"8b3982b0",
          6369 => x"94518539",
          6370 => x"82b09c51",
          6371 => x"ffb3f43f",
          6372 => x"843d0d04",
          6373 => x"7188800c",
          6374 => x"04ff3d0d",
          6375 => x"87c09684",
          6376 => x"70085252",
          6377 => x"80720c70",
          6378 => x"74077082",
          6379 => x"ba940c72",
          6380 => x"0c833d0d",
          6381 => x"04ff3d0d",
          6382 => x"87c09684",
          6383 => x"700882ba",
          6384 => x"940c5280",
          6385 => x"720c7309",
          6386 => x"7082ba94",
          6387 => x"08067082",
          6388 => x"ba940c73",
          6389 => x"0c51833d",
          6390 => x"0d04800b",
          6391 => x"87c09684",
          6392 => x"0c0482ba",
          6393 => x"940887c0",
          6394 => x"96840c04",
          6395 => x"fd3d0d76",
          6396 => x"982b7098",
          6397 => x"2c79982b",
          6398 => x"70982c72",
          6399 => x"10137082",
          6400 => x"2b515351",
          6401 => x"54515180",
          6402 => x"0b82b0a8",
          6403 => x"12335553",
          6404 => x"7174259c",
          6405 => x"3882b0a4",
          6406 => x"11081202",
          6407 => x"84059705",
          6408 => x"33713352",
          6409 => x"52527072",
          6410 => x"2e098106",
          6411 => x"83388153",
          6412 => x"7282bb98",
          6413 => x"0c853d0d",
          6414 => x"04fc3d0d",
          6415 => x"78028405",
          6416 => x"9f053371",
          6417 => x"33545553",
          6418 => x"71802ea2",
          6419 => x"388851ff",
          6420 => x"b5d33fa0",
          6421 => x"51ffb5cd",
          6422 => x"3f8851ff",
          6423 => x"b5c73f72",
          6424 => x"33ff0552",
          6425 => x"71733471",
          6426 => x"81ff0652",
          6427 => x"db397651",
          6428 => x"ffb2903f",
          6429 => x"73733486",
          6430 => x"3d0d04f6",
          6431 => x"3d0d7c02",
          6432 => x"8405b705",
          6433 => x"33028805",
          6434 => x"bb053382",
          6435 => x"baf03370",
          6436 => x"842982ba",
          6437 => x"98057008",
          6438 => x"5159595a",
          6439 => x"58597480",
          6440 => x"2e863874",
          6441 => x"519ab53f",
          6442 => x"82baf033",
          6443 => x"70842982",
          6444 => x"ba980581",
          6445 => x"19705458",
          6446 => x"565a9db6",
          6447 => x"3f82bb98",
          6448 => x"08750c82",
          6449 => x"baf03370",
          6450 => x"842982ba",
          6451 => x"98057008",
          6452 => x"51565a74",
          6453 => x"802ea738",
          6454 => x"75537852",
          6455 => x"7451ffbf",
          6456 => x"a43f82ba",
          6457 => x"f0338105",
          6458 => x"557482ba",
          6459 => x"f0347481",
          6460 => x"ff065593",
          6461 => x"75278738",
          6462 => x"800b82ba",
          6463 => x"f0347780",
          6464 => x"2eb63882",
          6465 => x"baec0856",
          6466 => x"75802eac",
          6467 => x"3882bae8",
          6468 => x"335574a4",
          6469 => x"388c3dfc",
          6470 => x"05547653",
          6471 => x"78527551",
          6472 => x"80d9c33f",
          6473 => x"82baec08",
          6474 => x"528a5181",
          6475 => x"8ed03f82",
          6476 => x"baec0851",
          6477 => x"80dda03f",
          6478 => x"8c3d0d04",
          6479 => x"fd3d0d82",
          6480 => x"ba985393",
          6481 => x"54720852",
          6482 => x"71802e89",
          6483 => x"38715199",
          6484 => x"8b3f8073",
          6485 => x"0cff1484",
          6486 => x"14545473",
          6487 => x"8025e638",
          6488 => x"800b82ba",
          6489 => x"f03482ba",
          6490 => x"ec085271",
          6491 => x"802e9538",
          6492 => x"715180de",
          6493 => x"803f82ba",
          6494 => x"ec085198",
          6495 => x"df3f800b",
          6496 => x"82baec0c",
          6497 => x"853d0d04",
          6498 => x"dc3d0d81",
          6499 => x"57805282",
          6500 => x"baec0851",
          6501 => x"80e2ed3f",
          6502 => x"82bb9808",
          6503 => x"80d33882",
          6504 => x"baec0853",
          6505 => x"80f85288",
          6506 => x"3d705256",
          6507 => x"818bbb3f",
          6508 => x"82bb9808",
          6509 => x"802eba38",
          6510 => x"7551ffbb",
          6511 => x"e83f82bb",
          6512 => x"98085580",
          6513 => x"0b82bb98",
          6514 => x"08259d38",
          6515 => x"82bb9808",
          6516 => x"ff057017",
          6517 => x"55558074",
          6518 => x"34755376",
          6519 => x"52811782",
          6520 => x"b3985257",
          6521 => x"ff87ef3f",
          6522 => x"74ff2e09",
          6523 => x"8106ffaf",
          6524 => x"38a63d0d",
          6525 => x"04d93d0d",
          6526 => x"aa3d08ad",
          6527 => x"3d085a5a",
          6528 => x"81705858",
          6529 => x"805282ba",
          6530 => x"ec085180",
          6531 => x"e1f63f82",
          6532 => x"bb980881",
          6533 => x"9538ff0b",
          6534 => x"82baec08",
          6535 => x"545580f8",
          6536 => x"528b3d70",
          6537 => x"5256818a",
          6538 => x"c13f82bb",
          6539 => x"9808802e",
          6540 => x"a5387551",
          6541 => x"ffbaee3f",
          6542 => x"82bb9808",
          6543 => x"81185855",
          6544 => x"800b82bb",
          6545 => x"9808258e",
          6546 => x"3882bb98",
          6547 => x"08ff0570",
          6548 => x"17555580",
          6549 => x"74347409",
          6550 => x"70307072",
          6551 => x"079f2a51",
          6552 => x"55557877",
          6553 => x"2e853873",
          6554 => x"ffac3882",
          6555 => x"baec088c",
          6556 => x"11085351",
          6557 => x"80e18d3f",
          6558 => x"82bb9808",
          6559 => x"802e8938",
          6560 => x"82b3a451",
          6561 => x"ffadfc3f",
          6562 => x"78772e09",
          6563 => x"81069b38",
          6564 => x"75527951",
          6565 => x"ffbafc3f",
          6566 => x"7951ffba",
          6567 => x"883fab3d",
          6568 => x"085482bb",
          6569 => x"98087434",
          6570 => x"80587782",
          6571 => x"bb980ca9",
          6572 => x"3d0d04f6",
          6573 => x"3d0d7c7e",
          6574 => x"715c7172",
          6575 => x"3357595a",
          6576 => x"5873a02e",
          6577 => x"098106a2",
          6578 => x"38783378",
          6579 => x"05567776",
          6580 => x"27983881",
          6581 => x"17705b70",
          6582 => x"71335658",
          6583 => x"5573a02e",
          6584 => x"09810686",
          6585 => x"38757526",
          6586 => x"ea388054",
          6587 => x"73882982",
          6588 => x"baf40570",
          6589 => x"085255ff",
          6590 => x"b9ab3f82",
          6591 => x"bb980853",
          6592 => x"79527408",
          6593 => x"51ffbcaa",
          6594 => x"3f82bb98",
          6595 => x"0880c638",
          6596 => x"84153355",
          6597 => x"74812e88",
          6598 => x"3874822e",
          6599 => x"8838b639",
          6600 => x"fce63fad",
          6601 => x"39811a5a",
          6602 => x"8c3dfc11",
          6603 => x"53f80551",
          6604 => x"ffa6ff3f",
          6605 => x"82bb9808",
          6606 => x"802e9a38",
          6607 => x"ff1b5378",
          6608 => x"527751fd",
          6609 => x"b03f82bb",
          6610 => x"980881ff",
          6611 => x"06557485",
          6612 => x"38745491",
          6613 => x"39811470",
          6614 => x"81ff0651",
          6615 => x"54827427",
          6616 => x"ff8a3880",
          6617 => x"547382bb",
          6618 => x"980c8c3d",
          6619 => x"0d04d33d",
          6620 => x"0db03d08",
          6621 => x"b23d08b4",
          6622 => x"3d08595f",
          6623 => x"5a800baf",
          6624 => x"3d3482ba",
          6625 => x"f03382ba",
          6626 => x"ec08555b",
          6627 => x"7381cb38",
          6628 => x"7382bae8",
          6629 => x"33555573",
          6630 => x"83388155",
          6631 => x"76802e81",
          6632 => x"bc388170",
          6633 => x"76065556",
          6634 => x"73802e81",
          6635 => x"ad38a851",
          6636 => x"97c03f82",
          6637 => x"bb980882",
          6638 => x"baec0c82",
          6639 => x"bb980880",
          6640 => x"2e819238",
          6641 => x"93537652",
          6642 => x"82bb9808",
          6643 => x"5180ccb4",
          6644 => x"3f82bb98",
          6645 => x"08802e8c",
          6646 => x"3882b3d0",
          6647 => x"51ffaba3",
          6648 => x"3f80f739",
          6649 => x"82bb9808",
          6650 => x"5b82baec",
          6651 => x"085380f8",
          6652 => x"52903d70",
          6653 => x"52548186",
          6654 => x"f13f82bb",
          6655 => x"98085682",
          6656 => x"bb980874",
          6657 => x"2e098106",
          6658 => x"80d03882",
          6659 => x"bb980851",
          6660 => x"ffb7923f",
          6661 => x"82bb9808",
          6662 => x"55800b82",
          6663 => x"bb980825",
          6664 => x"a93882bb",
          6665 => x"9808ff05",
          6666 => x"70175555",
          6667 => x"80743480",
          6668 => x"537481ff",
          6669 => x"06527551",
          6670 => x"f8c13f81",
          6671 => x"1b7081ff",
          6672 => x"065c5493",
          6673 => x"7b278338",
          6674 => x"805b74ff",
          6675 => x"2e098106",
          6676 => x"ff973886",
          6677 => x"397582ba",
          6678 => x"e834768c",
          6679 => x"3882baec",
          6680 => x"08802e84",
          6681 => x"38f9d53f",
          6682 => x"8f3d5dec",
          6683 => x"903f82bb",
          6684 => x"9808982b",
          6685 => x"70982c51",
          6686 => x"5978ff2e",
          6687 => x"ee387881",
          6688 => x"ff0682d2",
          6689 => x"c4337098",
          6690 => x"2b70982c",
          6691 => x"82d2c033",
          6692 => x"70982b70",
          6693 => x"972c7198",
          6694 => x"2c057084",
          6695 => x"2982b0a4",
          6696 => x"05700815",
          6697 => x"70335151",
          6698 => x"51515959",
          6699 => x"51595d58",
          6700 => x"81567378",
          6701 => x"2e80e938",
          6702 => x"777427b4",
          6703 => x"38748180",
          6704 => x"0a2981ff",
          6705 => x"0a057098",
          6706 => x"2c515580",
          6707 => x"752480ce",
          6708 => x"38765374",
          6709 => x"527751f6",
          6710 => x"933f82bb",
          6711 => x"980881ff",
          6712 => x"06547380",
          6713 => x"2ed73874",
          6714 => x"82d2c034",
          6715 => x"8156b139",
          6716 => x"7481800a",
          6717 => x"2981800a",
          6718 => x"0570982c",
          6719 => x"7081ff06",
          6720 => x"56515573",
          6721 => x"95269738",
          6722 => x"76537452",
          6723 => x"7751f5dc",
          6724 => x"3f82bb98",
          6725 => x"0881ff06",
          6726 => x"5473cc38",
          6727 => x"d3398056",
          6728 => x"75802e80",
          6729 => x"ca38811c",
          6730 => x"557482d2",
          6731 => x"c4347498",
          6732 => x"2b70982c",
          6733 => x"82d2c033",
          6734 => x"70982b70",
          6735 => x"982c7010",
          6736 => x"1170822b",
          6737 => x"82b0a811",
          6738 => x"335e5151",
          6739 => x"51575851",
          6740 => x"5574772e",
          6741 => x"098106fe",
          6742 => x"923882b0",
          6743 => x"ac14087d",
          6744 => x"0c800b82",
          6745 => x"d2c43480",
          6746 => x"0b82d2c0",
          6747 => x"34923975",
          6748 => x"82d2c434",
          6749 => x"7582d2c0",
          6750 => x"3478af3d",
          6751 => x"34757d0c",
          6752 => x"7e547395",
          6753 => x"26fde138",
          6754 => x"73842982",
          6755 => x"9a940554",
          6756 => x"73080482",
          6757 => x"d2cc3354",
          6758 => x"737e2efd",
          6759 => x"cb3882d2",
          6760 => x"c8335573",
          6761 => x"7527ab38",
          6762 => x"74982b70",
          6763 => x"982c5155",
          6764 => x"7375249e",
          6765 => x"38741a54",
          6766 => x"73338115",
          6767 => x"34748180",
          6768 => x"0a2981ff",
          6769 => x"0a057098",
          6770 => x"2c82d2cc",
          6771 => x"33565155",
          6772 => x"df3982d2",
          6773 => x"cc338111",
          6774 => x"56547482",
          6775 => x"d2cc3473",
          6776 => x"1a54ae3d",
          6777 => x"33743482",
          6778 => x"d2c83354",
          6779 => x"737e2589",
          6780 => x"38811454",
          6781 => x"7382d2c8",
          6782 => x"3482d2cc",
          6783 => x"33708180",
          6784 => x"0a2981ff",
          6785 => x"0a057098",
          6786 => x"2c82d2c8",
          6787 => x"335a5156",
          6788 => x"56747725",
          6789 => x"a338741a",
          6790 => x"70335254",
          6791 => x"ffaa863f",
          6792 => x"7481800a",
          6793 => x"2981800a",
          6794 => x"0570982c",
          6795 => x"82d2c833",
          6796 => x"56515573",
          6797 => x"7524df38",
          6798 => x"82d2cc33",
          6799 => x"70982b70",
          6800 => x"982c82d2",
          6801 => x"c8335a51",
          6802 => x"56567477",
          6803 => x"25fc9938",
          6804 => x"8851ffa9",
          6805 => x"d03f7481",
          6806 => x"800a2981",
          6807 => x"800a0570",
          6808 => x"982c82d2",
          6809 => x"c8335651",
          6810 => x"55737524",
          6811 => x"e338fbf8",
          6812 => x"39837a34",
          6813 => x"800b811b",
          6814 => x"3482d2cc",
          6815 => x"53805282",
          6816 => x"a98851f3",
          6817 => x"b43f81e4",
          6818 => x"3982d2cc",
          6819 => x"337081ff",
          6820 => x"06555573",
          6821 => x"802efbd0",
          6822 => x"3882d2c8",
          6823 => x"33ff0554",
          6824 => x"7382d2c8",
          6825 => x"34ff1554",
          6826 => x"7382d2cc",
          6827 => x"348851ff",
          6828 => x"a8f33f82",
          6829 => x"d2cc3370",
          6830 => x"982b7098",
          6831 => x"2c82d2c8",
          6832 => x"33575156",
          6833 => x"57747425",
          6834 => x"a838741a",
          6835 => x"54811433",
          6836 => x"74347333",
          6837 => x"51ffa8cd",
          6838 => x"3f748180",
          6839 => x"0a298180",
          6840 => x"0a057098",
          6841 => x"2c82d2c8",
          6842 => x"33585155",
          6843 => x"757524da",
          6844 => x"38a051ff",
          6845 => x"a8af3f82",
          6846 => x"d2cc3370",
          6847 => x"982b7098",
          6848 => x"2c82d2c8",
          6849 => x"33575156",
          6850 => x"57747424",
          6851 => x"fada3888",
          6852 => x"51ffa891",
          6853 => x"3f748180",
          6854 => x"0a298180",
          6855 => x"0a057098",
          6856 => x"2c82d2c8",
          6857 => x"33585155",
          6858 => x"757525e3",
          6859 => x"38fab939",
          6860 => x"82d2c833",
          6861 => x"7a055480",
          6862 => x"74348a51",
          6863 => x"ffa7e63f",
          6864 => x"82d2c852",
          6865 => x"7951f6eb",
          6866 => x"3f82bb98",
          6867 => x"0881ff06",
          6868 => x"54739638",
          6869 => x"82d2c833",
          6870 => x"5473802e",
          6871 => x"8f388153",
          6872 => x"73527951",
          6873 => x"f2953f84",
          6874 => x"39807a34",
          6875 => x"800b82d2",
          6876 => x"cc34800b",
          6877 => x"82d2c834",
          6878 => x"7982bb98",
          6879 => x"0caf3d0d",
          6880 => x"0482d2cc",
          6881 => x"33547380",
          6882 => x"2ef9dd38",
          6883 => x"8851ffa7",
          6884 => x"943f82d2",
          6885 => x"cc33ff05",
          6886 => x"547382d2",
          6887 => x"cc347381",
          6888 => x"ff0654e2",
          6889 => x"3982d2cc",
          6890 => x"3382d2c8",
          6891 => x"33555573",
          6892 => x"752ef9b4",
          6893 => x"38ff1454",
          6894 => x"7382d2c8",
          6895 => x"3474982b",
          6896 => x"70982c75",
          6897 => x"81ff0656",
          6898 => x"51557474",
          6899 => x"25a83874",
          6900 => x"1a548114",
          6901 => x"33743473",
          6902 => x"3351ffa6",
          6903 => x"c83f7481",
          6904 => x"800a2981",
          6905 => x"800a0570",
          6906 => x"982c82d2",
          6907 => x"c8335851",
          6908 => x"55757524",
          6909 => x"da38a051",
          6910 => x"ffa6aa3f",
          6911 => x"82d2cc33",
          6912 => x"70982b70",
          6913 => x"982c82d2",
          6914 => x"c8335751",
          6915 => x"56577474",
          6916 => x"24f8d538",
          6917 => x"8851ffa6",
          6918 => x"8c3f7481",
          6919 => x"800a2981",
          6920 => x"800a0570",
          6921 => x"982c82d2",
          6922 => x"c8335851",
          6923 => x"55757525",
          6924 => x"e338f8b4",
          6925 => x"3982d2cc",
          6926 => x"337081ff",
          6927 => x"0682d2c8",
          6928 => x"33595654",
          6929 => x"747727f8",
          6930 => x"9f388114",
          6931 => x"547382d2",
          6932 => x"cc34741a",
          6933 => x"70335254",
          6934 => x"ffa5ca3f",
          6935 => x"82d2cc33",
          6936 => x"7081ff06",
          6937 => x"82d2c833",
          6938 => x"58565475",
          6939 => x"7526db38",
          6940 => x"f7f63982",
          6941 => x"d2cc5380",
          6942 => x"5282a988",
          6943 => x"51efba3f",
          6944 => x"800b82d2",
          6945 => x"cc34800b",
          6946 => x"82d2c834",
          6947 => x"f7da397a",
          6948 => x"b03882ba",
          6949 => x"e4085574",
          6950 => x"802ea638",
          6951 => x"7451ffae",
          6952 => x"843f82bb",
          6953 => x"980882d2",
          6954 => x"c83482bb",
          6955 => x"980881ff",
          6956 => x"06810553",
          6957 => x"74527951",
          6958 => x"ffafca3f",
          6959 => x"935b81c0",
          6960 => x"397a8429",
          6961 => x"82ba9805",
          6962 => x"fc110856",
          6963 => x"5474802e",
          6964 => x"a7387451",
          6965 => x"ffadce3f",
          6966 => x"82bb9808",
          6967 => x"82d2c834",
          6968 => x"82bb9808",
          6969 => x"81ff0681",
          6970 => x"05537452",
          6971 => x"7951ffaf",
          6972 => x"943fff1b",
          6973 => x"5480fa39",
          6974 => x"73085574",
          6975 => x"802ef6e8",
          6976 => x"387451ff",
          6977 => x"ad9f3f99",
          6978 => x"397a932e",
          6979 => x"098106ae",
          6980 => x"3882ba98",
          6981 => x"08557480",
          6982 => x"2ea43874",
          6983 => x"51ffad85",
          6984 => x"3f82bb98",
          6985 => x"0882d2c8",
          6986 => x"3482bb98",
          6987 => x"0881ff06",
          6988 => x"81055374",
          6989 => x"527951ff",
          6990 => x"aecb3f80",
          6991 => x"c3397a84",
          6992 => x"2982ba9c",
          6993 => x"05700856",
          6994 => x"5474802e",
          6995 => x"ab387451",
          6996 => x"ffacd23f",
          6997 => x"82bb9808",
          6998 => x"82d2c834",
          6999 => x"82bb9808",
          7000 => x"81ff0681",
          7001 => x"05537452",
          7002 => x"7951ffae",
          7003 => x"983f811b",
          7004 => x"547381ff",
          7005 => x"065b8939",
          7006 => x"7482d2c8",
          7007 => x"34747a34",
          7008 => x"82d2cc53",
          7009 => x"82d2c833",
          7010 => x"527951ed",
          7011 => x"ac3ff5d8",
          7012 => x"3982d2cc",
          7013 => x"337081ff",
          7014 => x"0682d2c8",
          7015 => x"33595654",
          7016 => x"747727f5",
          7017 => x"c3388114",
          7018 => x"547382d2",
          7019 => x"cc34741a",
          7020 => x"70335254",
          7021 => x"ffa2ee3f",
          7022 => x"f5ae3982",
          7023 => x"d2cc3354",
          7024 => x"73802ef5",
          7025 => x"a3388851",
          7026 => x"ffa2da3f",
          7027 => x"82d2cc33",
          7028 => x"ff055473",
          7029 => x"82d2cc34",
          7030 => x"f58e39f9",
          7031 => x"3d0d83c0",
          7032 => x"800b82bb",
          7033 => x"900c8480",
          7034 => x"0b82bb8c",
          7035 => x"23a08053",
          7036 => x"805283c0",
          7037 => x"8051ffb2",
          7038 => x"8d3f82bb",
          7039 => x"90085480",
          7040 => x"58777434",
          7041 => x"81577681",
          7042 => x"153482bb",
          7043 => x"90085477",
          7044 => x"84153476",
          7045 => x"85153482",
          7046 => x"bb900854",
          7047 => x"77861534",
          7048 => x"76871534",
          7049 => x"82bb9008",
          7050 => x"82bb8c22",
          7051 => x"ff05fe80",
          7052 => x"80077083",
          7053 => x"ffff0670",
          7054 => x"882a5851",
          7055 => x"55567488",
          7056 => x"17347389",
          7057 => x"173482bb",
          7058 => x"8c227088",
          7059 => x"2982bb90",
          7060 => x"0805f811",
          7061 => x"51555577",
          7062 => x"82153476",
          7063 => x"83153489",
          7064 => x"3d0d04ff",
          7065 => x"3d0d7352",
          7066 => x"81518472",
          7067 => x"278f38fb",
          7068 => x"12832a82",
          7069 => x"117083ff",
          7070 => x"ff065151",
          7071 => x"517082bb",
          7072 => x"980c833d",
          7073 => x"0d04f93d",
          7074 => x"0d02a605",
          7075 => x"22028405",
          7076 => x"aa052271",
          7077 => x"0582bb90",
          7078 => x"0871832b",
          7079 => x"71117483",
          7080 => x"2b731170",
          7081 => x"33811233",
          7082 => x"71882b07",
          7083 => x"02a405ae",
          7084 => x"05227181",
          7085 => x"ffff0607",
          7086 => x"70882a53",
          7087 => x"51525954",
          7088 => x"5b5b5753",
          7089 => x"54557177",
          7090 => x"34708118",
          7091 => x"3482bb90",
          7092 => x"08147588",
          7093 => x"2a525470",
          7094 => x"82153474",
          7095 => x"83153482",
          7096 => x"bb900870",
          7097 => x"17703381",
          7098 => x"12337188",
          7099 => x"2b077083",
          7100 => x"2b8ffff8",
          7101 => x"06515256",
          7102 => x"52710573",
          7103 => x"83ffff06",
          7104 => x"70882a54",
          7105 => x"54517182",
          7106 => x"12347281",
          7107 => x"ff065372",
          7108 => x"83123482",
          7109 => x"bb900816",
          7110 => x"56717634",
          7111 => x"72811734",
          7112 => x"893d0d04",
          7113 => x"fb3d0d82",
          7114 => x"bb900802",
          7115 => x"84059e05",
          7116 => x"2270832b",
          7117 => x"72118611",
          7118 => x"33871233",
          7119 => x"718b2b71",
          7120 => x"832b0758",
          7121 => x"5b595255",
          7122 => x"52720584",
          7123 => x"12338513",
          7124 => x"3371882b",
          7125 => x"0770882a",
          7126 => x"54565652",
          7127 => x"70841334",
          7128 => x"73851334",
          7129 => x"82bb9008",
          7130 => x"70148411",
          7131 => x"33851233",
          7132 => x"718b2b71",
          7133 => x"832b0756",
          7134 => x"59575272",
          7135 => x"05861233",
          7136 => x"87133371",
          7137 => x"882b0770",
          7138 => x"882a5456",
          7139 => x"56527086",
          7140 => x"13347387",
          7141 => x"133482bb",
          7142 => x"90081370",
          7143 => x"33811233",
          7144 => x"71882b07",
          7145 => x"7081ffff",
          7146 => x"0670882a",
          7147 => x"53515353",
          7148 => x"53717334",
          7149 => x"70811434",
          7150 => x"873d0d04",
          7151 => x"fa3d0d02",
          7152 => x"a2052282",
          7153 => x"bb900871",
          7154 => x"832b7111",
          7155 => x"70338112",
          7156 => x"3371882b",
          7157 => x"07708829",
          7158 => x"15703381",
          7159 => x"12337198",
          7160 => x"2b71902b",
          7161 => x"07535f53",
          7162 => x"55525a56",
          7163 => x"57535471",
          7164 => x"802580f6",
          7165 => x"387251fe",
          7166 => x"ab3f82bb",
          7167 => x"90087016",
          7168 => x"70338112",
          7169 => x"33718b2b",
          7170 => x"71832b07",
          7171 => x"74117033",
          7172 => x"81123371",
          7173 => x"882b0770",
          7174 => x"832b8fff",
          7175 => x"f8065152",
          7176 => x"5451535a",
          7177 => x"58537205",
          7178 => x"74882a54",
          7179 => x"52728213",
          7180 => x"34738313",
          7181 => x"3482bb90",
          7182 => x"08701670",
          7183 => x"33811233",
          7184 => x"718b2b71",
          7185 => x"832b0756",
          7186 => x"59575572",
          7187 => x"05703381",
          7188 => x"12337188",
          7189 => x"2b077081",
          7190 => x"ffff0670",
          7191 => x"882a5751",
          7192 => x"52585272",
          7193 => x"74347181",
          7194 => x"1534883d",
          7195 => x"0d04fb3d",
          7196 => x"0d82bb90",
          7197 => x"08028405",
          7198 => x"9e052270",
          7199 => x"832b7211",
          7200 => x"82113383",
          7201 => x"1233718b",
          7202 => x"2b71832b",
          7203 => x"07595b59",
          7204 => x"52565273",
          7205 => x"05713381",
          7206 => x"13337188",
          7207 => x"2b07028c",
          7208 => x"05a20522",
          7209 => x"71077088",
          7210 => x"2a535153",
          7211 => x"53537173",
          7212 => x"34708114",
          7213 => x"3482bb90",
          7214 => x"08701570",
          7215 => x"33811233",
          7216 => x"718b2b71",
          7217 => x"832b0756",
          7218 => x"59575272",
          7219 => x"05821233",
          7220 => x"83133371",
          7221 => x"882b0770",
          7222 => x"882a5455",
          7223 => x"56527082",
          7224 => x"13347283",
          7225 => x"133482bb",
          7226 => x"90081482",
          7227 => x"11338312",
          7228 => x"3371882b",
          7229 => x"0782bb98",
          7230 => x"0c525487",
          7231 => x"3d0d04f7",
          7232 => x"3d0d7b82",
          7233 => x"bb900831",
          7234 => x"832a7083",
          7235 => x"ffff0670",
          7236 => x"535753fd",
          7237 => x"a73f82bb",
          7238 => x"90087683",
          7239 => x"2b711182",
          7240 => x"11338312",
          7241 => x"33718b2b",
          7242 => x"71832b07",
          7243 => x"75117033",
          7244 => x"81123371",
          7245 => x"982b7190",
          7246 => x"2b075342",
          7247 => x"4051535b",
          7248 => x"58555954",
          7249 => x"7280258d",
          7250 => x"38828080",
          7251 => x"527551fe",
          7252 => x"9d3f8184",
          7253 => x"39841433",
          7254 => x"85153371",
          7255 => x"8b2b7183",
          7256 => x"2b077611",
          7257 => x"79882a53",
          7258 => x"51555855",
          7259 => x"76861434",
          7260 => x"7581ff06",
          7261 => x"56758714",
          7262 => x"3482bb90",
          7263 => x"08701984",
          7264 => x"12338513",
          7265 => x"3371882b",
          7266 => x"0770882a",
          7267 => x"54575b56",
          7268 => x"53728416",
          7269 => x"34738516",
          7270 => x"3482bb90",
          7271 => x"08185380",
          7272 => x"0b861434",
          7273 => x"800b8714",
          7274 => x"3482bb90",
          7275 => x"08537684",
          7276 => x"14347585",
          7277 => x"143482bb",
          7278 => x"90081870",
          7279 => x"33811233",
          7280 => x"71882b07",
          7281 => x"70828080",
          7282 => x"0770882a",
          7283 => x"53515556",
          7284 => x"54747434",
          7285 => x"72811534",
          7286 => x"8b3d0d04",
          7287 => x"ff3d0d73",
          7288 => x"5282bb90",
          7289 => x"088438f7",
          7290 => x"f23f7180",
          7291 => x"2e863871",
          7292 => x"51fe8c3f",
          7293 => x"833d0d04",
          7294 => x"f53d0d80",
          7295 => x"7e5258f8",
          7296 => x"e23f82bb",
          7297 => x"980883ff",
          7298 => x"ff0682bb",
          7299 => x"90088411",
          7300 => x"33851233",
          7301 => x"71882b07",
          7302 => x"705f5956",
          7303 => x"585a81ff",
          7304 => x"ff597578",
          7305 => x"2e80cb38",
          7306 => x"75882917",
          7307 => x"70338112",
          7308 => x"3371882b",
          7309 => x"077081ff",
          7310 => x"ff067931",
          7311 => x"7083ffff",
          7312 => x"06707f27",
          7313 => x"52535156",
          7314 => x"59557779",
          7315 => x"278a3873",
          7316 => x"802e8538",
          7317 => x"75785a5b",
          7318 => x"84153385",
          7319 => x"16337188",
          7320 => x"2b075754",
          7321 => x"75c23878",
          7322 => x"81ffff2e",
          7323 => x"85387a79",
          7324 => x"59568076",
          7325 => x"832b82bb",
          7326 => x"90081170",
          7327 => x"33811233",
          7328 => x"71882b07",
          7329 => x"7081ffff",
          7330 => x"0651525a",
          7331 => x"565c5573",
          7332 => x"752e8338",
          7333 => x"81558054",
          7334 => x"79782681",
          7335 => x"cc387454",
          7336 => x"74802e81",
          7337 => x"c438777a",
          7338 => x"2e098106",
          7339 => x"89387551",
          7340 => x"f8f23f81",
          7341 => x"ac398280",
          7342 => x"80537952",
          7343 => x"7551f7c6",
          7344 => x"3f82bb90",
          7345 => x"08701c86",
          7346 => x"11338712",
          7347 => x"33718b2b",
          7348 => x"71832b07",
          7349 => x"535a5e55",
          7350 => x"74057a17",
          7351 => x"7083ffff",
          7352 => x"0670882a",
          7353 => x"5c595654",
          7354 => x"78841534",
          7355 => x"7681ff06",
          7356 => x"57768515",
          7357 => x"3482bb90",
          7358 => x"0875832b",
          7359 => x"7111721e",
          7360 => x"86113387",
          7361 => x"12337188",
          7362 => x"2b077088",
          7363 => x"2a535b5e",
          7364 => x"535a5654",
          7365 => x"73861934",
          7366 => x"75871934",
          7367 => x"82bb9008",
          7368 => x"701c8411",
          7369 => x"33851233",
          7370 => x"718b2b71",
          7371 => x"832b0753",
          7372 => x"5d5a5574",
          7373 => x"05547886",
          7374 => x"15347687",
          7375 => x"153482bb",
          7376 => x"90087016",
          7377 => x"711d8411",
          7378 => x"33851233",
          7379 => x"71882b07",
          7380 => x"70882a53",
          7381 => x"5a5f5256",
          7382 => x"54738416",
          7383 => x"34758516",
          7384 => x"3482bb90",
          7385 => x"081b8405",
          7386 => x"547382bb",
          7387 => x"980c8d3d",
          7388 => x"0d04fe3d",
          7389 => x"0d745282",
          7390 => x"bb900884",
          7391 => x"38f4dc3f",
          7392 => x"71537180",
          7393 => x"2e8b3871",
          7394 => x"51fced3f",
          7395 => x"82bb9808",
          7396 => x"537282bb",
          7397 => x"980c843d",
          7398 => x"0d04ee3d",
          7399 => x"0d646640",
          7400 => x"5c807042",
          7401 => x"4082bb90",
          7402 => x"08602e09",
          7403 => x"81068438",
          7404 => x"f4a93f7b",
          7405 => x"8e387e51",
          7406 => x"ffb83f82",
          7407 => x"bb980854",
          7408 => x"83c7397e",
          7409 => x"8b387b51",
          7410 => x"fc923f7e",
          7411 => x"5483ba39",
          7412 => x"7e51f58f",
          7413 => x"3f82bb98",
          7414 => x"0883ffff",
          7415 => x"0682bb90",
          7416 => x"087d7131",
          7417 => x"832a7083",
          7418 => x"ffff0670",
          7419 => x"832b7311",
          7420 => x"70338112",
          7421 => x"3371882b",
          7422 => x"07707531",
          7423 => x"7083ffff",
          7424 => x"06708829",
          7425 => x"fc057388",
          7426 => x"291a7033",
          7427 => x"81123371",
          7428 => x"882b0770",
          7429 => x"902b5344",
          7430 => x"4e534841",
          7431 => x"525c545b",
          7432 => x"415c565b",
          7433 => x"5b738025",
          7434 => x"8f387681",
          7435 => x"ffff0675",
          7436 => x"317083ff",
          7437 => x"ff064254",
          7438 => x"82163383",
          7439 => x"17337188",
          7440 => x"2b077088",
          7441 => x"291c7033",
          7442 => x"81123371",
          7443 => x"982b7190",
          7444 => x"2b075347",
          7445 => x"45525654",
          7446 => x"7380258b",
          7447 => x"38787531",
          7448 => x"7083ffff",
          7449 => x"06415477",
          7450 => x"7b2781fe",
          7451 => x"38601854",
          7452 => x"737b2e09",
          7453 => x"81068f38",
          7454 => x"7851f6c0",
          7455 => x"3f7a83ff",
          7456 => x"ff065881",
          7457 => x"e5397f8e",
          7458 => x"387a7424",
          7459 => x"89387851",
          7460 => x"f6aa3f81",
          7461 => x"a5397f18",
          7462 => x"557a7524",
          7463 => x"80c83879",
          7464 => x"1d821133",
          7465 => x"83123371",
          7466 => x"882b0753",
          7467 => x"5754f4f4",
          7468 => x"3f805278",
          7469 => x"51f7b73f",
          7470 => x"82bb9808",
          7471 => x"83ffff06",
          7472 => x"7e547c53",
          7473 => x"70832b82",
          7474 => x"bb900811",
          7475 => x"84055355",
          7476 => x"59ff9ae7",
          7477 => x"3f82bb90",
          7478 => x"08148405",
          7479 => x"7583ffff",
          7480 => x"06595c81",
          7481 => x"85396015",
          7482 => x"547a7424",
          7483 => x"80d43878",
          7484 => x"51f5c93f",
          7485 => x"82bb9008",
          7486 => x"1d821133",
          7487 => x"83123371",
          7488 => x"882b0753",
          7489 => x"4354f49c",
          7490 => x"3f805278",
          7491 => x"51f6df3f",
          7492 => x"82bb9808",
          7493 => x"83ffff06",
          7494 => x"7e547c53",
          7495 => x"70832b82",
          7496 => x"bb900811",
          7497 => x"84055355",
          7498 => x"59ff9a8f",
          7499 => x"3f82bb90",
          7500 => x"08148405",
          7501 => x"60620519",
          7502 => x"555c7383",
          7503 => x"ffff0658",
          7504 => x"a9397b7f",
          7505 => x"5254f9b0",
          7506 => x"3f82bb98",
          7507 => x"085c82bb",
          7508 => x"9808802e",
          7509 => x"93387d53",
          7510 => x"735282bb",
          7511 => x"980851ff",
          7512 => x"9ea33f73",
          7513 => x"51f7983f",
          7514 => x"7a587a78",
          7515 => x"27993880",
          7516 => x"537a5278",
          7517 => x"51f28f3f",
          7518 => x"7a19832b",
          7519 => x"82bb9008",
          7520 => x"05840551",
          7521 => x"f6f93f7b",
          7522 => x"547382bb",
          7523 => x"980c943d",
          7524 => x"0d04fc3d",
          7525 => x"0d777729",
          7526 => x"705254fb",
          7527 => x"d53f82bb",
          7528 => x"98085582",
          7529 => x"bb980880",
          7530 => x"2e8e3873",
          7531 => x"53805282",
          7532 => x"bb980851",
          7533 => x"ffa2cf3f",
          7534 => x"7482bb98",
          7535 => x"0c863d0d",
          7536 => x"04ff3d0d",
          7537 => x"028f0533",
          7538 => x"51815270",
          7539 => x"72268738",
          7540 => x"82bb9411",
          7541 => x"33527182",
          7542 => x"bb980c83",
          7543 => x"3d0d04fc",
          7544 => x"3d0d029b",
          7545 => x"05330284",
          7546 => x"059f0533",
          7547 => x"56538351",
          7548 => x"72812680",
          7549 => x"e0387284",
          7550 => x"2b87c092",
          7551 => x"8c115351",
          7552 => x"88547480",
          7553 => x"2e843881",
          7554 => x"88547372",
          7555 => x"0c87c092",
          7556 => x"8c115181",
          7557 => x"710c850b",
          7558 => x"87c0988c",
          7559 => x"0c705271",
          7560 => x"08708206",
          7561 => x"51517080",
          7562 => x"2e8a3887",
          7563 => x"c0988c08",
          7564 => x"5170ec38",
          7565 => x"7108fc80",
          7566 => x"80065271",
          7567 => x"923887c0",
          7568 => x"988c0851",
          7569 => x"70802e87",
          7570 => x"387182bb",
          7571 => x"94143482",
          7572 => x"bb941333",
          7573 => x"517082bb",
          7574 => x"980c863d",
          7575 => x"0d04f33d",
          7576 => x"0d606264",
          7577 => x"028c05bf",
          7578 => x"05335740",
          7579 => x"585b8374",
          7580 => x"525afecd",
          7581 => x"3f82bb98",
          7582 => x"0881067a",
          7583 => x"54527181",
          7584 => x"be387172",
          7585 => x"75842b87",
          7586 => x"c0928011",
          7587 => x"87c0928c",
          7588 => x"1287c092",
          7589 => x"8413415a",
          7590 => x"40575a58",
          7591 => x"850b87c0",
          7592 => x"988c0c76",
          7593 => x"7d0c8476",
          7594 => x"0c750870",
          7595 => x"852a7081",
          7596 => x"06515354",
          7597 => x"71802e8e",
          7598 => x"387b0852",
          7599 => x"717b7081",
          7600 => x"055d3481",
          7601 => x"19598074",
          7602 => x"a2065353",
          7603 => x"71732e83",
          7604 => x"38815378",
          7605 => x"83ff268f",
          7606 => x"3872802e",
          7607 => x"8a3887c0",
          7608 => x"988c0852",
          7609 => x"71c33887",
          7610 => x"c0988c08",
          7611 => x"5271802e",
          7612 => x"87387884",
          7613 => x"802e9938",
          7614 => x"81760c87",
          7615 => x"c0928c15",
          7616 => x"53720870",
          7617 => x"82065152",
          7618 => x"71f738ff",
          7619 => x"1a5a8d39",
          7620 => x"84801781",
          7621 => x"197081ff",
          7622 => x"065a5357",
          7623 => x"79802e90",
          7624 => x"3873fc80",
          7625 => x"80065271",
          7626 => x"87387d78",
          7627 => x"26feed38",
          7628 => x"73fc8080",
          7629 => x"06527180",
          7630 => x"2e833881",
          7631 => x"52715372",
          7632 => x"82bb980c",
          7633 => x"8f3d0d04",
          7634 => x"f33d0d60",
          7635 => x"6264028c",
          7636 => x"05bf0533",
          7637 => x"5740585b",
          7638 => x"83598074",
          7639 => x"5258fce1",
          7640 => x"3f82bb98",
          7641 => x"08810679",
          7642 => x"54527178",
          7643 => x"2e098106",
          7644 => x"81b13877",
          7645 => x"74842b87",
          7646 => x"c0928011",
          7647 => x"87c0928c",
          7648 => x"1287c092",
          7649 => x"84134059",
          7650 => x"5f565a85",
          7651 => x"0b87c098",
          7652 => x"8c0c767d",
          7653 => x"0c82760c",
          7654 => x"80587508",
          7655 => x"70842a70",
          7656 => x"81065153",
          7657 => x"5471802e",
          7658 => x"8c387a70",
          7659 => x"81055c33",
          7660 => x"7c0c8118",
          7661 => x"5873812a",
          7662 => x"70810651",
          7663 => x"5271802e",
          7664 => x"8a3887c0",
          7665 => x"988c0852",
          7666 => x"71d03887",
          7667 => x"c0988c08",
          7668 => x"5271802e",
          7669 => x"87387784",
          7670 => x"802e9938",
          7671 => x"81760c87",
          7672 => x"c0928c15",
          7673 => x"53720870",
          7674 => x"82065152",
          7675 => x"71f738ff",
          7676 => x"19598d39",
          7677 => x"811a7081",
          7678 => x"ff068480",
          7679 => x"19595b52",
          7680 => x"78802e90",
          7681 => x"3873fc80",
          7682 => x"80065271",
          7683 => x"87387d7a",
          7684 => x"26fef838",
          7685 => x"73fc8080",
          7686 => x"06527180",
          7687 => x"2e833881",
          7688 => x"52715372",
          7689 => x"82bb980c",
          7690 => x"8f3d0d04",
          7691 => x"fa3d0d7a",
          7692 => x"028405a3",
          7693 => x"05330288",
          7694 => x"05a70533",
          7695 => x"71545456",
          7696 => x"57fafe3f",
          7697 => x"82bb9808",
          7698 => x"81065383",
          7699 => x"547280fe",
          7700 => x"38850b87",
          7701 => x"c0988c0c",
          7702 => x"81567176",
          7703 => x"2e80dc38",
          7704 => x"71762493",
          7705 => x"3874842b",
          7706 => x"87c0928c",
          7707 => x"11545471",
          7708 => x"802e8d38",
          7709 => x"80d43971",
          7710 => x"832e80c6",
          7711 => x"3880cb39",
          7712 => x"72087081",
          7713 => x"2a708106",
          7714 => x"51515271",
          7715 => x"802e8a38",
          7716 => x"87c0988c",
          7717 => x"085271e8",
          7718 => x"3887c098",
          7719 => x"8c085271",
          7720 => x"96388173",
          7721 => x"0c87c092",
          7722 => x"8c145372",
          7723 => x"08708206",
          7724 => x"515271f7",
          7725 => x"38963980",
          7726 => x"56923988",
          7727 => x"800a770c",
          7728 => x"85398180",
          7729 => x"770c7256",
          7730 => x"83398456",
          7731 => x"75547382",
          7732 => x"bb980c88",
          7733 => x"3d0d04fe",
          7734 => x"3d0d7481",
          7735 => x"11337133",
          7736 => x"71882b07",
          7737 => x"82bb980c",
          7738 => x"5351843d",
          7739 => x"0d04fd3d",
          7740 => x"0d758311",
          7741 => x"33821233",
          7742 => x"71902b71",
          7743 => x"882b0781",
          7744 => x"14337072",
          7745 => x"07882b75",
          7746 => x"33710782",
          7747 => x"bb980c52",
          7748 => x"53545654",
          7749 => x"52853d0d",
          7750 => x"04ff3d0d",
          7751 => x"73028405",
          7752 => x"92052252",
          7753 => x"52707270",
          7754 => x"81055434",
          7755 => x"70882a51",
          7756 => x"70723483",
          7757 => x"3d0d04ff",
          7758 => x"3d0d7375",
          7759 => x"52527072",
          7760 => x"70810554",
          7761 => x"3470882a",
          7762 => x"51707270",
          7763 => x"81055434",
          7764 => x"70882a51",
          7765 => x"70727081",
          7766 => x"05543470",
          7767 => x"882a5170",
          7768 => x"7234833d",
          7769 => x"0d04fe3d",
          7770 => x"0d767577",
          7771 => x"54545170",
          7772 => x"802e9238",
          7773 => x"71708105",
          7774 => x"53337370",
          7775 => x"81055534",
          7776 => x"ff1151eb",
          7777 => x"39843d0d",
          7778 => x"04fe3d0d",
          7779 => x"75777654",
          7780 => x"52537272",
          7781 => x"70810554",
          7782 => x"34ff1151",
          7783 => x"70f43884",
          7784 => x"3d0d04fc",
          7785 => x"3d0d7877",
          7786 => x"79565653",
          7787 => x"74708105",
          7788 => x"56337470",
          7789 => x"81055633",
          7790 => x"717131ff",
          7791 => x"16565252",
          7792 => x"5272802e",
          7793 => x"86387180",
          7794 => x"2ee23871",
          7795 => x"82bb980c",
          7796 => x"863d0d04",
          7797 => x"fe3d0d74",
          7798 => x"76545189",
          7799 => x"3971732e",
          7800 => x"8a388111",
          7801 => x"51703352",
          7802 => x"71f33870",
          7803 => x"3382bb98",
          7804 => x"0c843d0d",
          7805 => x"04800b82",
          7806 => x"bb980c04",
          7807 => x"800b82bb",
          7808 => x"980c04f7",
          7809 => x"3d0d7b56",
          7810 => x"800b8317",
          7811 => x"33565a74",
          7812 => x"7a2e80d6",
          7813 => x"388154b0",
          7814 => x"160853b4",
          7815 => x"16705381",
          7816 => x"17335259",
          7817 => x"faa23f82",
          7818 => x"bb98087a",
          7819 => x"2e098106",
          7820 => x"b73882bb",
          7821 => x"98088317",
          7822 => x"34b01608",
          7823 => x"70a41808",
          7824 => x"319c1808",
          7825 => x"59565874",
          7826 => x"77279f38",
          7827 => x"82163355",
          7828 => x"74822e09",
          7829 => x"81069338",
          7830 => x"81547618",
          7831 => x"53785281",
          7832 => x"163351f9",
          7833 => x"e33f8339",
          7834 => x"815a7982",
          7835 => x"bb980c8b",
          7836 => x"3d0d04fa",
          7837 => x"3d0d787a",
          7838 => x"56568057",
          7839 => x"74b01708",
          7840 => x"2eaf3875",
          7841 => x"51fefc3f",
          7842 => x"82bb9808",
          7843 => x"5782bb98",
          7844 => x"089f3881",
          7845 => x"547453b4",
          7846 => x"16528116",
          7847 => x"3351f7be",
          7848 => x"3f82bb98",
          7849 => x"08802e85",
          7850 => x"38ff5581",
          7851 => x"5774b017",
          7852 => x"0c7682bb",
          7853 => x"980c883d",
          7854 => x"0d04f83d",
          7855 => x"0d7a7052",
          7856 => x"57fec03f",
          7857 => x"82bb9808",
          7858 => x"5882bb98",
          7859 => x"08819138",
          7860 => x"76335574",
          7861 => x"832e0981",
          7862 => x"0680f038",
          7863 => x"84173359",
          7864 => x"78812e09",
          7865 => x"810680e3",
          7866 => x"38848053",
          7867 => x"82bb9808",
          7868 => x"52b41770",
          7869 => x"5256fd91",
          7870 => x"3f82d4d5",
          7871 => x"5284b217",
          7872 => x"51fc963f",
          7873 => x"848b85a4",
          7874 => x"d2527551",
          7875 => x"fca93f86",
          7876 => x"8a85e4f2",
          7877 => x"52849817",
          7878 => x"51fc9c3f",
          7879 => x"90170852",
          7880 => x"849c1751",
          7881 => x"fc913f8c",
          7882 => x"17085284",
          7883 => x"a01751fc",
          7884 => x"863fa017",
          7885 => x"08810570",
          7886 => x"b0190c79",
          7887 => x"55537552",
          7888 => x"81173351",
          7889 => x"f8823f77",
          7890 => x"84183480",
          7891 => x"53805281",
          7892 => x"173351f9",
          7893 => x"d73f82bb",
          7894 => x"9808802e",
          7895 => x"83388158",
          7896 => x"7782bb98",
          7897 => x"0c8a3d0d",
          7898 => x"04fb3d0d",
          7899 => x"77fe1a98",
          7900 => x"1208fe05",
          7901 => x"55565480",
          7902 => x"56747327",
          7903 => x"8d388a14",
          7904 => x"22757129",
          7905 => x"ac160805",
          7906 => x"57537582",
          7907 => x"bb980c87",
          7908 => x"3d0d04f9",
          7909 => x"3d0d7a7a",
          7910 => x"70085654",
          7911 => x"57817727",
          7912 => x"81df3876",
          7913 => x"98150827",
          7914 => x"81d738ff",
          7915 => x"74335458",
          7916 => x"72822e80",
          7917 => x"f5387282",
          7918 => x"24893872",
          7919 => x"812e8d38",
          7920 => x"81bf3972",
          7921 => x"832e818e",
          7922 => x"3881b639",
          7923 => x"76812a17",
          7924 => x"70892aa4",
          7925 => x"16080553",
          7926 => x"745255fd",
          7927 => x"963f82bb",
          7928 => x"9808819f",
          7929 => x"387483ff",
          7930 => x"0614b411",
          7931 => x"33811770",
          7932 => x"892aa418",
          7933 => x"08055576",
          7934 => x"54575753",
          7935 => x"fcf53f82",
          7936 => x"bb980880",
          7937 => x"fe387483",
          7938 => x"ff0614b4",
          7939 => x"11337088",
          7940 => x"2b780779",
          7941 => x"81067184",
          7942 => x"2a5c5258",
          7943 => x"51537280",
          7944 => x"e238759f",
          7945 => x"ff065880",
          7946 => x"da397688",
          7947 => x"2aa41508",
          7948 => x"05527351",
          7949 => x"fcbd3f82",
          7950 => x"bb980880",
          7951 => x"c6387610",
          7952 => x"83fe0674",
          7953 => x"05b40551",
          7954 => x"f98d3f82",
          7955 => x"bb980883",
          7956 => x"ffff0658",
          7957 => x"ae397687",
          7958 => x"2aa41508",
          7959 => x"05527351",
          7960 => x"fc913f82",
          7961 => x"bb98089b",
          7962 => x"3876822b",
          7963 => x"83fc0674",
          7964 => x"05b40551",
          7965 => x"f8f83f82",
          7966 => x"bb9808f0",
          7967 => x"0a065883",
          7968 => x"39815877",
          7969 => x"82bb980c",
          7970 => x"893d0d04",
          7971 => x"f83d0d7a",
          7972 => x"7c7e5a58",
          7973 => x"56825981",
          7974 => x"7727829e",
          7975 => x"38769817",
          7976 => x"08278296",
          7977 => x"38753353",
          7978 => x"72792e81",
          7979 => x"9d387279",
          7980 => x"24893872",
          7981 => x"812e8d38",
          7982 => x"82803972",
          7983 => x"832e81b8",
          7984 => x"3881f739",
          7985 => x"76812a17",
          7986 => x"70892aa4",
          7987 => x"18080553",
          7988 => x"765255fb",
          7989 => x"9e3f82bb",
          7990 => x"98085982",
          7991 => x"bb980881",
          7992 => x"d9387483",
          7993 => x"ff0616b4",
          7994 => x"05811678",
          7995 => x"81065956",
          7996 => x"54775376",
          7997 => x"802e8f38",
          7998 => x"77842b9f",
          7999 => x"f0067433",
          8000 => x"8f067107",
          8001 => x"51537274",
          8002 => x"34810b83",
          8003 => x"17347489",
          8004 => x"2aa41708",
          8005 => x"05527551",
          8006 => x"fad93f82",
          8007 => x"bb980859",
          8008 => x"82bb9808",
          8009 => x"81943874",
          8010 => x"83ff0616",
          8011 => x"b4057884",
          8012 => x"2a545476",
          8013 => x"8f387788",
          8014 => x"2a743381",
          8015 => x"f006718f",
          8016 => x"06075153",
          8017 => x"72743480",
          8018 => x"ec397688",
          8019 => x"2aa41708",
          8020 => x"05527551",
          8021 => x"fa9d3f82",
          8022 => x"bb980859",
          8023 => x"82bb9808",
          8024 => x"80d83877",
          8025 => x"83ffff06",
          8026 => x"52761083",
          8027 => x"fe067605",
          8028 => x"b40551f7",
          8029 => x"a43fbe39",
          8030 => x"76872aa4",
          8031 => x"17080552",
          8032 => x"7551f9ef",
          8033 => x"3f82bb98",
          8034 => x"085982bb",
          8035 => x"9808ab38",
          8036 => x"77f00a06",
          8037 => x"77822b83",
          8038 => x"fc067018",
          8039 => x"b4057054",
          8040 => x"515454f6",
          8041 => x"c93f82bb",
          8042 => x"98088f0a",
          8043 => x"06740752",
          8044 => x"7251f783",
          8045 => x"3f810b83",
          8046 => x"17347882",
          8047 => x"bb980c8a",
          8048 => x"3d0d04f8",
          8049 => x"3d0d7a7c",
          8050 => x"7e720859",
          8051 => x"56565981",
          8052 => x"7527a438",
          8053 => x"74981708",
          8054 => x"279d3873",
          8055 => x"802eaa38",
          8056 => x"ff537352",
          8057 => x"7551fda4",
          8058 => x"3f82bb98",
          8059 => x"085482bb",
          8060 => x"980880f2",
          8061 => x"38933982",
          8062 => x"5480eb39",
          8063 => x"815480e6",
          8064 => x"3982bb98",
          8065 => x"085480de",
          8066 => x"39745278",
          8067 => x"51fb843f",
          8068 => x"82bb9808",
          8069 => x"5882bb98",
          8070 => x"08802e80",
          8071 => x"c73882bb",
          8072 => x"9808812e",
          8073 => x"d23882bb",
          8074 => x"9808ff2e",
          8075 => x"cf388053",
          8076 => x"74527551",
          8077 => x"fcd63f82",
          8078 => x"bb9808c5",
          8079 => x"38981608",
          8080 => x"fe119018",
          8081 => x"08575557",
          8082 => x"74742790",
          8083 => x"38811590",
          8084 => x"170c8416",
          8085 => x"33810754",
          8086 => x"73841734",
          8087 => x"77557678",
          8088 => x"26ffa638",
          8089 => x"80547382",
          8090 => x"bb980c8a",
          8091 => x"3d0d04f6",
          8092 => x"3d0d7c7e",
          8093 => x"7108595b",
          8094 => x"5b799538",
          8095 => x"8c170858",
          8096 => x"77802e88",
          8097 => x"38981708",
          8098 => x"7826b238",
          8099 => x"8158ae39",
          8100 => x"79527a51",
          8101 => x"f9fd3f81",
          8102 => x"557482bb",
          8103 => x"98082782",
          8104 => x"e03882bb",
          8105 => x"98085582",
          8106 => x"bb9808ff",
          8107 => x"2e82d238",
          8108 => x"98170882",
          8109 => x"bb980826",
          8110 => x"82c73879",
          8111 => x"58901708",
          8112 => x"70565473",
          8113 => x"802e82b9",
          8114 => x"38777a2e",
          8115 => x"09810680",
          8116 => x"e238811a",
          8117 => x"56981708",
          8118 => x"76268338",
          8119 => x"82567552",
          8120 => x"7a51f9af",
          8121 => x"3f805982",
          8122 => x"bb980881",
          8123 => x"2e098106",
          8124 => x"863882bb",
          8125 => x"98085982",
          8126 => x"bb980809",
          8127 => x"70307072",
          8128 => x"07802570",
          8129 => x"7c0782bb",
          8130 => x"98085451",
          8131 => x"51555573",
          8132 => x"81ef3882",
          8133 => x"bb980880",
          8134 => x"2e95388c",
          8135 => x"17085481",
          8136 => x"74279038",
          8137 => x"73981808",
          8138 => x"27893873",
          8139 => x"58853975",
          8140 => x"80db3877",
          8141 => x"56811656",
          8142 => x"98170876",
          8143 => x"26893882",
          8144 => x"56757826",
          8145 => x"81ac3875",
          8146 => x"527a51f8",
          8147 => x"c63f82bb",
          8148 => x"9808802e",
          8149 => x"b8388059",
          8150 => x"82bb9808",
          8151 => x"812e0981",
          8152 => x"06863882",
          8153 => x"bb980859",
          8154 => x"82bb9808",
          8155 => x"09703070",
          8156 => x"72078025",
          8157 => x"707c0751",
          8158 => x"51555573",
          8159 => x"80f83875",
          8160 => x"782e0981",
          8161 => x"06ffae38",
          8162 => x"735580f5",
          8163 => x"39ff5375",
          8164 => x"527651f9",
          8165 => x"f73f82bb",
          8166 => x"980882bb",
          8167 => x"98083070",
          8168 => x"82bb9808",
          8169 => x"07802551",
          8170 => x"55557980",
          8171 => x"2e943873",
          8172 => x"802e8f38",
          8173 => x"75537952",
          8174 => x"7651f9d0",
          8175 => x"3f82bb98",
          8176 => x"085574a5",
          8177 => x"38758c18",
          8178 => x"0c981708",
          8179 => x"fe059018",
          8180 => x"08565474",
          8181 => x"74268638",
          8182 => x"ff159018",
          8183 => x"0c841733",
          8184 => x"81075473",
          8185 => x"84183497",
          8186 => x"39ff5674",
          8187 => x"812e9038",
          8188 => x"8c398055",
          8189 => x"8c3982bb",
          8190 => x"98085585",
          8191 => x"39815675",
          8192 => x"557482bb",
          8193 => x"980c8c3d",
          8194 => x"0d04f83d",
          8195 => x"0d7a7052",
          8196 => x"55f3f03f",
          8197 => x"82bb9808",
          8198 => x"58815682",
          8199 => x"bb980880",
          8200 => x"d8387b52",
          8201 => x"7451f6c1",
          8202 => x"3f82bb98",
          8203 => x"0882bb98",
          8204 => x"08b0170c",
          8205 => x"59848053",
          8206 => x"7752b415",
          8207 => x"705257f2",
          8208 => x"c83f7756",
          8209 => x"84398116",
          8210 => x"568a1522",
          8211 => x"58757827",
          8212 => x"97388154",
          8213 => x"75195376",
          8214 => x"52811533",
          8215 => x"51ede93f",
          8216 => x"82bb9808",
          8217 => x"802edf38",
          8218 => x"8a152276",
          8219 => x"32703070",
          8220 => x"7207709f",
          8221 => x"2a535156",
          8222 => x"567582bb",
          8223 => x"980c8a3d",
          8224 => x"0d04f83d",
          8225 => x"0d7a7c71",
          8226 => x"08585657",
          8227 => x"74f0800a",
          8228 => x"2680f138",
          8229 => x"749f0653",
          8230 => x"7280e938",
          8231 => x"7490180c",
          8232 => x"88170854",
          8233 => x"73aa3875",
          8234 => x"33538273",
          8235 => x"278838a8",
          8236 => x"16085473",
          8237 => x"9b387485",
          8238 => x"2a53820b",
          8239 => x"8817225a",
          8240 => x"58727927",
          8241 => x"80fe38a8",
          8242 => x"16089818",
          8243 => x"0c80cd39",
          8244 => x"8a162270",
          8245 => x"892b5458",
          8246 => x"727526b2",
          8247 => x"38735276",
          8248 => x"51f5b03f",
          8249 => x"82bb9808",
          8250 => x"5482bb98",
          8251 => x"08ff2ebd",
          8252 => x"38810b82",
          8253 => x"bb980827",
          8254 => x"8b389816",
          8255 => x"0882bb98",
          8256 => x"08268538",
          8257 => x"8258bd39",
          8258 => x"74733155",
          8259 => x"cb397352",
          8260 => x"7551f4d5",
          8261 => x"3f82bb98",
          8262 => x"0898180c",
          8263 => x"7394180c",
          8264 => x"98170853",
          8265 => x"82587280",
          8266 => x"2e9a3885",
          8267 => x"39815894",
          8268 => x"3974892a",
          8269 => x"1398180c",
          8270 => x"7483ff06",
          8271 => x"16b4059c",
          8272 => x"180c8058",
          8273 => x"7782bb98",
          8274 => x"0c8a3d0d",
          8275 => x"04f83d0d",
          8276 => x"7a700890",
          8277 => x"1208a005",
          8278 => x"595754f0",
          8279 => x"800a7727",
          8280 => x"8638800b",
          8281 => x"98150c98",
          8282 => x"14085384",
          8283 => x"5572802e",
          8284 => x"81cb3876",
          8285 => x"83ff0658",
          8286 => x"7781b538",
          8287 => x"81139815",
          8288 => x"0c941408",
          8289 => x"55749238",
          8290 => x"76852a88",
          8291 => x"17225653",
          8292 => x"74732681",
          8293 => x"9b3880c0",
          8294 => x"398a1622",
          8295 => x"ff057789",
          8296 => x"2a065372",
          8297 => x"818a3874",
          8298 => x"527351f3",
          8299 => x"e63f82bb",
          8300 => x"98085382",
          8301 => x"55810b82",
          8302 => x"bb980827",
          8303 => x"80ff3881",
          8304 => x"5582bb98",
          8305 => x"08ff2e80",
          8306 => x"f4389816",
          8307 => x"0882bb98",
          8308 => x"082680ca",
          8309 => x"387b8a38",
          8310 => x"7798150c",
          8311 => x"845580dd",
          8312 => x"39941408",
          8313 => x"527351f9",
          8314 => x"863f82bb",
          8315 => x"98085387",
          8316 => x"5582bb98",
          8317 => x"08802e80",
          8318 => x"c4388255",
          8319 => x"82bb9808",
          8320 => x"812eba38",
          8321 => x"815582bb",
          8322 => x"9808ff2e",
          8323 => x"b03882bb",
          8324 => x"98085275",
          8325 => x"51fbf33f",
          8326 => x"82bb9808",
          8327 => x"a0387294",
          8328 => x"150c7252",
          8329 => x"7551f2c1",
          8330 => x"3f82bb98",
          8331 => x"0898150c",
          8332 => x"7690150c",
          8333 => x"7716b405",
          8334 => x"9c150c80",
          8335 => x"557482bb",
          8336 => x"980c8a3d",
          8337 => x"0d04f73d",
          8338 => x"0d7b7d71",
          8339 => x"085b5b57",
          8340 => x"80527651",
          8341 => x"fcac3f82",
          8342 => x"bb980854",
          8343 => x"82bb9808",
          8344 => x"80ec3882",
          8345 => x"bb980856",
          8346 => x"98170852",
          8347 => x"7851f083",
          8348 => x"3f82bb98",
          8349 => x"085482bb",
          8350 => x"980880d2",
          8351 => x"3882bb98",
          8352 => x"089c1808",
          8353 => x"70335154",
          8354 => x"587281e5",
          8355 => x"2e098106",
          8356 => x"83388158",
          8357 => x"82bb9808",
          8358 => x"55728338",
          8359 => x"81557775",
          8360 => x"07537280",
          8361 => x"2e8e3881",
          8362 => x"1656757a",
          8363 => x"2e098106",
          8364 => x"8838a539",
          8365 => x"82bb9808",
          8366 => x"56815276",
          8367 => x"51fd8e3f",
          8368 => x"82bb9808",
          8369 => x"5482bb98",
          8370 => x"08802eff",
          8371 => x"9b387384",
          8372 => x"2e098106",
          8373 => x"83388754",
          8374 => x"7382bb98",
          8375 => x"0c8b3d0d",
          8376 => x"04fd3d0d",
          8377 => x"769a1152",
          8378 => x"54ebec3f",
          8379 => x"82bb9808",
          8380 => x"83ffff06",
          8381 => x"76703351",
          8382 => x"53537183",
          8383 => x"2e098106",
          8384 => x"90389414",
          8385 => x"51ebd03f",
          8386 => x"82bb9808",
          8387 => x"902b7307",
          8388 => x"537282bb",
          8389 => x"980c853d",
          8390 => x"0d04fc3d",
          8391 => x"0d777970",
          8392 => x"83ffff06",
          8393 => x"549a1253",
          8394 => x"5555ebed",
          8395 => x"3f767033",
          8396 => x"51537283",
          8397 => x"2e098106",
          8398 => x"8b387390",
          8399 => x"2a529415",
          8400 => x"51ebd63f",
          8401 => x"863d0d04",
          8402 => x"f73d0d7b",
          8403 => x"7d5b5584",
          8404 => x"75085a58",
          8405 => x"98150880",
          8406 => x"2e818a38",
          8407 => x"98150852",
          8408 => x"7851ee8f",
          8409 => x"3f82bb98",
          8410 => x"085882bb",
          8411 => x"980880f5",
          8412 => x"389c1508",
          8413 => x"70335553",
          8414 => x"73863884",
          8415 => x"5880e639",
          8416 => x"8b133370",
          8417 => x"bf067081",
          8418 => x"ff065851",
          8419 => x"53728616",
          8420 => x"3482bb98",
          8421 => x"08537381",
          8422 => x"e52e8338",
          8423 => x"815373ae",
          8424 => x"2ea93881",
          8425 => x"70740654",
          8426 => x"5772802e",
          8427 => x"9e38758f",
          8428 => x"2e993882",
          8429 => x"bb980876",
          8430 => x"df065454",
          8431 => x"72882e09",
          8432 => x"81068338",
          8433 => x"7654737a",
          8434 => x"2ea03880",
          8435 => x"527451fa",
          8436 => x"fc3f82bb",
          8437 => x"98085882",
          8438 => x"bb980889",
          8439 => x"38981508",
          8440 => x"fefa3886",
          8441 => x"39800b98",
          8442 => x"160c7782",
          8443 => x"bb980c8b",
          8444 => x"3d0d04fb",
          8445 => x"3d0d7770",
          8446 => x"08575481",
          8447 => x"527351fc",
          8448 => x"c53f82bb",
          8449 => x"98085582",
          8450 => x"bb9808b4",
          8451 => x"38981408",
          8452 => x"527551ec",
          8453 => x"de3f82bb",
          8454 => x"98085582",
          8455 => x"bb9808a0",
          8456 => x"38a05382",
          8457 => x"bb980852",
          8458 => x"9c140851",
          8459 => x"eadb3f8b",
          8460 => x"53a01452",
          8461 => x"9c140851",
          8462 => x"eaac3f81",
          8463 => x"0b831734",
          8464 => x"7482bb98",
          8465 => x"0c873d0d",
          8466 => x"04fd3d0d",
          8467 => x"75700898",
          8468 => x"12085470",
          8469 => x"535553ec",
          8470 => x"9a3f82bb",
          8471 => x"98088d38",
          8472 => x"9c130853",
          8473 => x"e5733481",
          8474 => x"0b831534",
          8475 => x"853d0d04",
          8476 => x"fa3d0d78",
          8477 => x"7a575780",
          8478 => x"0b891734",
          8479 => x"98170880",
          8480 => x"2e818238",
          8481 => x"80708918",
          8482 => x"5555559c",
          8483 => x"17081470",
          8484 => x"33811656",
          8485 => x"515271a0",
          8486 => x"2ea83871",
          8487 => x"852e0981",
          8488 => x"06843881",
          8489 => x"e5527389",
          8490 => x"2e098106",
          8491 => x"8b38ae73",
          8492 => x"70810555",
          8493 => x"34811555",
          8494 => x"71737081",
          8495 => x"05553481",
          8496 => x"15558a74",
          8497 => x"27c53875",
          8498 => x"15880552",
          8499 => x"800b8113",
          8500 => x"349c1708",
          8501 => x"528b1233",
          8502 => x"8817349c",
          8503 => x"17089c11",
          8504 => x"5252e88a",
          8505 => x"3f82bb98",
          8506 => x"08760c96",
          8507 => x"1251e7e7",
          8508 => x"3f82bb98",
          8509 => x"08861723",
          8510 => x"981251e7",
          8511 => x"da3f82bb",
          8512 => x"98088417",
          8513 => x"23883d0d",
          8514 => x"04f33d0d",
          8515 => x"7f70085e",
          8516 => x"5b806170",
          8517 => x"33515555",
          8518 => x"73af2e83",
          8519 => x"38815573",
          8520 => x"80dc2e91",
          8521 => x"3874802e",
          8522 => x"8c38941d",
          8523 => x"08881c0c",
          8524 => x"aa398115",
          8525 => x"41806170",
          8526 => x"33565656",
          8527 => x"73af2e09",
          8528 => x"81068338",
          8529 => x"81567380",
          8530 => x"dc327030",
          8531 => x"70802578",
          8532 => x"07515154",
          8533 => x"73dc3873",
          8534 => x"881c0c60",
          8535 => x"70335154",
          8536 => x"739f2696",
          8537 => x"38ff800b",
          8538 => x"ab1c3480",
          8539 => x"527a51f6",
          8540 => x"913f82bb",
          8541 => x"98085585",
          8542 => x"9839913d",
          8543 => x"61a01d5c",
          8544 => x"5a5e8b53",
          8545 => x"a0527951",
          8546 => x"e7ff3f80",
          8547 => x"70595788",
          8548 => x"7933555c",
          8549 => x"73ae2e09",
          8550 => x"810680d4",
          8551 => x"38781870",
          8552 => x"33811a71",
          8553 => x"ae327030",
          8554 => x"709f2a73",
          8555 => x"82260751",
          8556 => x"51535a57",
          8557 => x"54738c38",
          8558 => x"79175475",
          8559 => x"74348117",
          8560 => x"57db3975",
          8561 => x"af327030",
          8562 => x"709f2a51",
          8563 => x"51547580",
          8564 => x"dc2e8c38",
          8565 => x"73802e87",
          8566 => x"3875a026",
          8567 => x"82bd3877",
          8568 => x"197e0ca4",
          8569 => x"54a07627",
          8570 => x"82bd38a0",
          8571 => x"5482b839",
          8572 => x"78187033",
          8573 => x"811a5a57",
          8574 => x"54a07627",
          8575 => x"81fc3875",
          8576 => x"af327030",
          8577 => x"7780dc32",
          8578 => x"70307280",
          8579 => x"25718025",
          8580 => x"07515156",
          8581 => x"51557380",
          8582 => x"2eac3884",
          8583 => x"39811858",
          8584 => x"80781a70",
          8585 => x"33515555",
          8586 => x"73af2e09",
          8587 => x"81068338",
          8588 => x"81557380",
          8589 => x"dc327030",
          8590 => x"70802577",
          8591 => x"07515154",
          8592 => x"73db3881",
          8593 => x"b53975ae",
          8594 => x"2e098106",
          8595 => x"83388154",
          8596 => x"767c2774",
          8597 => x"07547380",
          8598 => x"2ea2387b",
          8599 => x"8b327030",
          8600 => x"77ae3270",
          8601 => x"30728025",
          8602 => x"719f2a07",
          8603 => x"53515651",
          8604 => x"557481a7",
          8605 => x"3888578b",
          8606 => x"5cfef539",
          8607 => x"75982b54",
          8608 => x"7380258c",
          8609 => x"387580ff",
          8610 => x"0682b4e0",
          8611 => x"11335754",
          8612 => x"7551e6e1",
          8613 => x"3f82bb98",
          8614 => x"08802eb2",
          8615 => x"38781870",
          8616 => x"33811a71",
          8617 => x"545a5654",
          8618 => x"e6d23f82",
          8619 => x"bb980880",
          8620 => x"2e80e838",
          8621 => x"ff1c5476",
          8622 => x"742780df",
          8623 => x"38791754",
          8624 => x"75743481",
          8625 => x"177a1155",
          8626 => x"57747434",
          8627 => x"a7397552",
          8628 => x"82b48051",
          8629 => x"e5fe3f82",
          8630 => x"bb9808bf",
          8631 => x"38ff9f16",
          8632 => x"54739926",
          8633 => x"8938e016",
          8634 => x"7081ff06",
          8635 => x"57547917",
          8636 => x"54757434",
          8637 => x"811757fd",
          8638 => x"f7397719",
          8639 => x"7e0c7680",
          8640 => x"2e993879",
          8641 => x"33547381",
          8642 => x"e52e0981",
          8643 => x"06843885",
          8644 => x"7a348454",
          8645 => x"a076278f",
          8646 => x"388b3986",
          8647 => x"5581f239",
          8648 => x"845680f3",
          8649 => x"39805473",
          8650 => x"8b1b3480",
          8651 => x"7b085852",
          8652 => x"7a51f2ce",
          8653 => x"3f82bb98",
          8654 => x"085682bb",
          8655 => x"980880d7",
          8656 => x"38981b08",
          8657 => x"527651e6",
          8658 => x"aa3f82bb",
          8659 => x"98085682",
          8660 => x"bb980880",
          8661 => x"c2389c1b",
          8662 => x"08703355",
          8663 => x"5573802e",
          8664 => x"ffbe388b",
          8665 => x"1533bf06",
          8666 => x"5473861c",
          8667 => x"348b1533",
          8668 => x"70832a70",
          8669 => x"81065155",
          8670 => x"58739238",
          8671 => x"8b537952",
          8672 => x"7451e49f",
          8673 => x"3f82bb98",
          8674 => x"08802e8b",
          8675 => x"3875527a",
          8676 => x"51f3ba3f",
          8677 => x"ff9f3975",
          8678 => x"ab1c3357",
          8679 => x"5574802e",
          8680 => x"bb387484",
          8681 => x"2e098106",
          8682 => x"80e73875",
          8683 => x"852a7081",
          8684 => x"0677822a",
          8685 => x"58515473",
          8686 => x"802e9638",
          8687 => x"75810654",
          8688 => x"73802efb",
          8689 => x"b538ff80",
          8690 => x"0bab1c34",
          8691 => x"805580c1",
          8692 => x"39758106",
          8693 => x"5473ba38",
          8694 => x"8555b639",
          8695 => x"75822a70",
          8696 => x"81065154",
          8697 => x"73ab3886",
          8698 => x"1b337084",
          8699 => x"2a708106",
          8700 => x"51555573",
          8701 => x"802ee138",
          8702 => x"901b0883",
          8703 => x"ff061db4",
          8704 => x"05527c51",
          8705 => x"f5db3f82",
          8706 => x"bb980888",
          8707 => x"1c0cfaea",
          8708 => x"397482bb",
          8709 => x"980c8f3d",
          8710 => x"0d04f63d",
          8711 => x"0d7c5bff",
          8712 => x"7b087071",
          8713 => x"7355595c",
          8714 => x"55597380",
          8715 => x"2e81c638",
          8716 => x"75708105",
          8717 => x"573370a0",
          8718 => x"26525271",
          8719 => x"ba2e8d38",
          8720 => x"70ee3871",
          8721 => x"ba2e0981",
          8722 => x"0681a538",
          8723 => x"7333d011",
          8724 => x"7081ff06",
          8725 => x"51525370",
          8726 => x"89269138",
          8727 => x"82147381",
          8728 => x"ff06d005",
          8729 => x"56527176",
          8730 => x"2e80f738",
          8731 => x"800b82b4",
          8732 => x"d0595577",
          8733 => x"087a5557",
          8734 => x"76708105",
          8735 => x"58337470",
          8736 => x"81055633",
          8737 => x"ff9f1253",
          8738 => x"53537099",
          8739 => x"268938e0",
          8740 => x"137081ff",
          8741 => x"065451ff",
          8742 => x"9f125170",
          8743 => x"99268938",
          8744 => x"e0127081",
          8745 => x"ff065351",
          8746 => x"7230709f",
          8747 => x"2a515172",
          8748 => x"722e0981",
          8749 => x"06853870",
          8750 => x"ffbe3872",
          8751 => x"30747732",
          8752 => x"70307072",
          8753 => x"079f2a73",
          8754 => x"9f2a0753",
          8755 => x"54545170",
          8756 => x"802e8f38",
          8757 => x"81158419",
          8758 => x"59558375",
          8759 => x"25ff9438",
          8760 => x"8b397483",
          8761 => x"24863874",
          8762 => x"767c0c59",
          8763 => x"78518639",
          8764 => x"82d2e433",
          8765 => x"517082bb",
          8766 => x"980c8c3d",
          8767 => x"0d04fa3d",
          8768 => x"0d785680",
          8769 => x"0b831734",
          8770 => x"ff0bb017",
          8771 => x"0c795275",
          8772 => x"51e2e03f",
          8773 => x"845582bb",
          8774 => x"98088180",
          8775 => x"3884b216",
          8776 => x"51dfb43f",
          8777 => x"82bb9808",
          8778 => x"83ffff06",
          8779 => x"54835573",
          8780 => x"82d4d52e",
          8781 => x"09810680",
          8782 => x"e338800b",
          8783 => x"b4173356",
          8784 => x"577481e9",
          8785 => x"2e098106",
          8786 => x"83388157",
          8787 => x"7481eb32",
          8788 => x"70307080",
          8789 => x"25790751",
          8790 => x"5154738a",
          8791 => x"387481e8",
          8792 => x"2e098106",
          8793 => x"b5388353",
          8794 => x"82b49052",
          8795 => x"80ea1651",
          8796 => x"e0b13f82",
          8797 => x"bb980855",
          8798 => x"82bb9808",
          8799 => x"802e9d38",
          8800 => x"855382b4",
          8801 => x"94528186",
          8802 => x"1651e097",
          8803 => x"3f82bb98",
          8804 => x"085582bb",
          8805 => x"9808802e",
          8806 => x"83388255",
          8807 => x"7482bb98",
          8808 => x"0c883d0d",
          8809 => x"04f23d0d",
          8810 => x"61028405",
          8811 => x"80cb0533",
          8812 => x"58558075",
          8813 => x"0c6051fc",
          8814 => x"e13f82bb",
          8815 => x"9808588b",
          8816 => x"56800b82",
          8817 => x"bb980824",
          8818 => x"86fc3882",
          8819 => x"bb980884",
          8820 => x"2982d2d0",
          8821 => x"05700855",
          8822 => x"538c5673",
          8823 => x"802e86e6",
          8824 => x"3873750c",
          8825 => x"7681fe06",
          8826 => x"74335457",
          8827 => x"72802eae",
          8828 => x"38811433",
          8829 => x"51d7ca3f",
          8830 => x"82bb9808",
          8831 => x"81ff0670",
          8832 => x"81065455",
          8833 => x"72983876",
          8834 => x"802e86b8",
          8835 => x"3874822a",
          8836 => x"70810651",
          8837 => x"538a5672",
          8838 => x"86ac3886",
          8839 => x"a7398074",
          8840 => x"34778115",
          8841 => x"34815281",
          8842 => x"143351d7",
          8843 => x"b23f82bb",
          8844 => x"980881ff",
          8845 => x"06708106",
          8846 => x"54558356",
          8847 => x"72868738",
          8848 => x"76802e8f",
          8849 => x"3874822a",
          8850 => x"70810651",
          8851 => x"538a5672",
          8852 => x"85f43880",
          8853 => x"70537452",
          8854 => x"5bfda33f",
          8855 => x"82bb9808",
          8856 => x"81ff0657",
          8857 => x"76822e09",
          8858 => x"810680e2",
          8859 => x"388c3d74",
          8860 => x"56588356",
          8861 => x"83f61533",
          8862 => x"70585372",
          8863 => x"802e8d38",
          8864 => x"83fa1551",
          8865 => x"dce83f82",
          8866 => x"bb980857",
          8867 => x"76787084",
          8868 => x"055a0cff",
          8869 => x"16901656",
          8870 => x"56758025",
          8871 => x"d738800b",
          8872 => x"8d3d5456",
          8873 => x"72708405",
          8874 => x"54085b83",
          8875 => x"577a802e",
          8876 => x"95387a52",
          8877 => x"7351fcc6",
          8878 => x"3f82bb98",
          8879 => x"0881ff06",
          8880 => x"57817727",
          8881 => x"89388116",
          8882 => x"56837627",
          8883 => x"d7388156",
          8884 => x"76842e84",
          8885 => x"f1388d56",
          8886 => x"76812684",
          8887 => x"e938bf14",
          8888 => x"51dbf43f",
          8889 => x"82bb9808",
          8890 => x"83ffff06",
          8891 => x"53728480",
          8892 => x"2e098106",
          8893 => x"84d03880",
          8894 => x"ca1451db",
          8895 => x"da3f82bb",
          8896 => x"980883ff",
          8897 => x"ff065877",
          8898 => x"8d3880d8",
          8899 => x"1451dbde",
          8900 => x"3f82bb98",
          8901 => x"0858779c",
          8902 => x"150c80c4",
          8903 => x"14338215",
          8904 => x"3480c414",
          8905 => x"33ff1170",
          8906 => x"81ff0651",
          8907 => x"54558d56",
          8908 => x"72812684",
          8909 => x"91387481",
          8910 => x"ff067871",
          8911 => x"2980c116",
          8912 => x"33525953",
          8913 => x"728a1523",
          8914 => x"72802e8b",
          8915 => x"38ff1373",
          8916 => x"06537280",
          8917 => x"2e86388d",
          8918 => x"5683eb39",
          8919 => x"80c51451",
          8920 => x"daf53f82",
          8921 => x"bb980853",
          8922 => x"82bb9808",
          8923 => x"88152372",
          8924 => x"8f06578d",
          8925 => x"567683ce",
          8926 => x"3880c714",
          8927 => x"51dad83f",
          8928 => x"82bb9808",
          8929 => x"83ffff06",
          8930 => x"55748d38",
          8931 => x"80d41451",
          8932 => x"dadc3f82",
          8933 => x"bb980855",
          8934 => x"80c21451",
          8935 => x"dab93f82",
          8936 => x"bb980883",
          8937 => x"ffff0653",
          8938 => x"8d567280",
          8939 => x"2e839738",
          8940 => x"88142278",
          8941 => x"1471842a",
          8942 => x"055a5a78",
          8943 => x"75268386",
          8944 => x"388a1422",
          8945 => x"52747931",
          8946 => x"51fefad7",
          8947 => x"3f82bb98",
          8948 => x"085582bb",
          8949 => x"9808802e",
          8950 => x"82ec3882",
          8951 => x"bb980880",
          8952 => x"fffffff5",
          8953 => x"26833883",
          8954 => x"577483ff",
          8955 => x"f5268338",
          8956 => x"8257749f",
          8957 => x"f5268538",
          8958 => x"81578939",
          8959 => x"8d567680",
          8960 => x"2e82c338",
          8961 => x"82157098",
          8962 => x"160c7ba0",
          8963 => x"160c731c",
          8964 => x"70a4170c",
          8965 => x"7a1dac17",
          8966 => x"0c545576",
          8967 => x"832e0981",
          8968 => x"06af3880",
          8969 => x"de1451d9",
          8970 => x"ae3f82bb",
          8971 => x"980883ff",
          8972 => x"ff06538d",
          8973 => x"5672828e",
          8974 => x"3879828a",
          8975 => x"3880e014",
          8976 => x"51d9ab3f",
          8977 => x"82bb9808",
          8978 => x"a8150c74",
          8979 => x"822b53a2",
          8980 => x"398d5679",
          8981 => x"802e81ee",
          8982 => x"387713a8",
          8983 => x"150c7415",
          8984 => x"5376822e",
          8985 => x"8d387410",
          8986 => x"1570812a",
          8987 => x"76810605",
          8988 => x"515383ff",
          8989 => x"13892a53",
          8990 => x"8d56729c",
          8991 => x"15082681",
          8992 => x"c538ff0b",
          8993 => x"90150cff",
          8994 => x"0b8c150c",
          8995 => x"ff800b84",
          8996 => x"15347683",
          8997 => x"2e098106",
          8998 => x"81923880",
          8999 => x"e41451d8",
          9000 => x"b63f82bb",
          9001 => x"980883ff",
          9002 => x"ff065372",
          9003 => x"812e0981",
          9004 => x"0680f938",
          9005 => x"811b5273",
          9006 => x"51dbb83f",
          9007 => x"82bb9808",
          9008 => x"80ea3882",
          9009 => x"bb980884",
          9010 => x"153484b2",
          9011 => x"1451d887",
          9012 => x"3f82bb98",
          9013 => x"0883ffff",
          9014 => x"06537282",
          9015 => x"d4d52e09",
          9016 => x"810680c8",
          9017 => x"38b41451",
          9018 => x"d8843f82",
          9019 => x"bb980884",
          9020 => x"8b85a4d2",
          9021 => x"2e098106",
          9022 => x"b3388498",
          9023 => x"1451d7ee",
          9024 => x"3f82bb98",
          9025 => x"08868a85",
          9026 => x"e4f22e09",
          9027 => x"81069d38",
          9028 => x"849c1451",
          9029 => x"d7d83f82",
          9030 => x"bb980890",
          9031 => x"150c84a0",
          9032 => x"1451d7ca",
          9033 => x"3f82bb98",
          9034 => x"088c150c",
          9035 => x"76743482",
          9036 => x"d2e02281",
          9037 => x"05537282",
          9038 => x"d2e02372",
          9039 => x"86152380",
          9040 => x"0b94150c",
          9041 => x"80567582",
          9042 => x"bb980c90",
          9043 => x"3d0d04fb",
          9044 => x"3d0d7754",
          9045 => x"89557380",
          9046 => x"2eb93873",
          9047 => x"08537280",
          9048 => x"2eb13872",
          9049 => x"33527180",
          9050 => x"2ea93886",
          9051 => x"13228415",
          9052 => x"22575271",
          9053 => x"762e0981",
          9054 => x"06993881",
          9055 => x"133351d0",
          9056 => x"c03f82bb",
          9057 => x"98088106",
          9058 => x"52718838",
          9059 => x"71740854",
          9060 => x"55833980",
          9061 => x"53787371",
          9062 => x"0c527482",
          9063 => x"bb980c87",
          9064 => x"3d0d04fa",
          9065 => x"3d0d02ab",
          9066 => x"05337a58",
          9067 => x"893dfc05",
          9068 => x"5256f4e6",
          9069 => x"3f8b5480",
          9070 => x"0b82bb98",
          9071 => x"0824bc38",
          9072 => x"82bb9808",
          9073 => x"842982d2",
          9074 => x"d0057008",
          9075 => x"55557380",
          9076 => x"2e843880",
          9077 => x"74347854",
          9078 => x"73802e84",
          9079 => x"38807434",
          9080 => x"78750c75",
          9081 => x"5475802e",
          9082 => x"92388053",
          9083 => x"893d7053",
          9084 => x"840551f7",
          9085 => x"b03f82bb",
          9086 => x"98085473",
          9087 => x"82bb980c",
          9088 => x"883d0d04",
          9089 => x"eb3d0d67",
          9090 => x"02840580",
          9091 => x"e7053359",
          9092 => x"59895478",
          9093 => x"802e84c8",
          9094 => x"3877bf06",
          9095 => x"7054983d",
          9096 => x"d0055399",
          9097 => x"3d840552",
          9098 => x"58f6fa3f",
          9099 => x"82bb9808",
          9100 => x"5582bb98",
          9101 => x"0884a438",
          9102 => x"7a5c6852",
          9103 => x"8c3d7052",
          9104 => x"56edc63f",
          9105 => x"82bb9808",
          9106 => x"5582bb98",
          9107 => x"08923802",
          9108 => x"80d70533",
          9109 => x"70982b55",
          9110 => x"57738025",
          9111 => x"83388655",
          9112 => x"779c0654",
          9113 => x"73802e81",
          9114 => x"ab387480",
          9115 => x"2e953874",
          9116 => x"842e0981",
          9117 => x"06aa3875",
          9118 => x"51eaf83f",
          9119 => x"82bb9808",
          9120 => x"559e3902",
          9121 => x"b2053391",
          9122 => x"06547381",
          9123 => x"b8387782",
          9124 => x"2a708106",
          9125 => x"51547380",
          9126 => x"2e8e3888",
          9127 => x"5583bc39",
          9128 => x"77880758",
          9129 => x"7483b438",
          9130 => x"77832a70",
          9131 => x"81065154",
          9132 => x"73802e81",
          9133 => x"af386252",
          9134 => x"7a51e8a5",
          9135 => x"3f82bb98",
          9136 => x"08568288",
          9137 => x"b20a5262",
          9138 => x"8e0551d4",
          9139 => x"ea3f6254",
          9140 => x"a00b8b15",
          9141 => x"34805362",
          9142 => x"527a51e8",
          9143 => x"bd3f8052",
          9144 => x"629c0551",
          9145 => x"d4d13f7a",
          9146 => x"54810b83",
          9147 => x"15347580",
          9148 => x"2e80f138",
          9149 => x"7ab01108",
          9150 => x"51548053",
          9151 => x"7552973d",
          9152 => x"d40551dd",
          9153 => x"be3f82bb",
          9154 => x"98085582",
          9155 => x"bb980882",
          9156 => x"ca38b739",
          9157 => x"7482c438",
          9158 => x"02b20533",
          9159 => x"70842a70",
          9160 => x"81065155",
          9161 => x"5673802e",
          9162 => x"86388455",
          9163 => x"82ad3977",
          9164 => x"812a7081",
          9165 => x"06515473",
          9166 => x"802ea938",
          9167 => x"75810654",
          9168 => x"73802ea0",
          9169 => x"38875582",
          9170 => x"92397352",
          9171 => x"7a51d6a3",
          9172 => x"3f82bb98",
          9173 => x"087bff18",
          9174 => x"8c120c55",
          9175 => x"5582bb98",
          9176 => x"0881f838",
          9177 => x"77832a70",
          9178 => x"81065154",
          9179 => x"73802e86",
          9180 => x"387780c0",
          9181 => x"07587ab0",
          9182 => x"1108a01b",
          9183 => x"0c63a41b",
          9184 => x"0c635370",
          9185 => x"5257e6d9",
          9186 => x"3f82bb98",
          9187 => x"0882bb98",
          9188 => x"08881b0c",
          9189 => x"639c0552",
          9190 => x"5ad2d33f",
          9191 => x"82bb9808",
          9192 => x"82bb9808",
          9193 => x"8c1b0c77",
          9194 => x"7a0c5686",
          9195 => x"1722841a",
          9196 => x"2377901a",
          9197 => x"34800b91",
          9198 => x"1a34800b",
          9199 => x"9c1a0c80",
          9200 => x"0b941a0c",
          9201 => x"77852a70",
          9202 => x"81065154",
          9203 => x"73802e81",
          9204 => x"8d3882bb",
          9205 => x"9808802e",
          9206 => x"81843882",
          9207 => x"bb980894",
          9208 => x"1a0c8a17",
          9209 => x"2270892b",
          9210 => x"7b525957",
          9211 => x"a8397652",
          9212 => x"7851d79f",
          9213 => x"3f82bb98",
          9214 => x"085782bb",
          9215 => x"98088126",
          9216 => x"83388255",
          9217 => x"82bb9808",
          9218 => x"ff2e0981",
          9219 => x"06833879",
          9220 => x"55757831",
          9221 => x"56743070",
          9222 => x"76078025",
          9223 => x"51547776",
          9224 => x"278a3881",
          9225 => x"70750655",
          9226 => x"5a73c338",
          9227 => x"76981a0c",
          9228 => x"74a93875",
          9229 => x"83ff0654",
          9230 => x"73802ea2",
          9231 => x"3876527a",
          9232 => x"51d6a63f",
          9233 => x"82bb9808",
          9234 => x"85388255",
          9235 => x"8e397589",
          9236 => x"2a82bb98",
          9237 => x"08059c1a",
          9238 => x"0c843980",
          9239 => x"790c7454",
          9240 => x"7382bb98",
          9241 => x"0c973d0d",
          9242 => x"04f23d0d",
          9243 => x"60636564",
          9244 => x"40405d59",
          9245 => x"807e0c90",
          9246 => x"3dfc0552",
          9247 => x"7851f9cf",
          9248 => x"3f82bb98",
          9249 => x"085582bb",
          9250 => x"98088a38",
          9251 => x"91193355",
          9252 => x"74802e86",
          9253 => x"38745682",
          9254 => x"c4399019",
          9255 => x"33810655",
          9256 => x"87567480",
          9257 => x"2e82b638",
          9258 => x"9539820b",
          9259 => x"911a3482",
          9260 => x"5682aa39",
          9261 => x"810b911a",
          9262 => x"34815682",
          9263 => x"a0398c19",
          9264 => x"08941a08",
          9265 => x"3155747c",
          9266 => x"27833874",
          9267 => x"5c7b802e",
          9268 => x"82893894",
          9269 => x"19087083",
          9270 => x"ff065656",
          9271 => x"7481b238",
          9272 => x"7e8a1122",
          9273 => x"ff057789",
          9274 => x"2a065b55",
          9275 => x"79a83875",
          9276 => x"87388819",
          9277 => x"08558f39",
          9278 => x"98190852",
          9279 => x"7851d593",
          9280 => x"3f82bb98",
          9281 => x"08558175",
          9282 => x"27ff9f38",
          9283 => x"74ff2eff",
          9284 => x"a3387498",
          9285 => x"1a0c9819",
          9286 => x"08527e51",
          9287 => x"d4cb3f82",
          9288 => x"bb980880",
          9289 => x"2eff8338",
          9290 => x"82bb9808",
          9291 => x"1a7c892a",
          9292 => x"59577780",
          9293 => x"2e80d638",
          9294 => x"771a7f8a",
          9295 => x"1122585c",
          9296 => x"55757527",
          9297 => x"8538757a",
          9298 => x"31587754",
          9299 => x"76537c52",
          9300 => x"811b3351",
          9301 => x"ca883f82",
          9302 => x"bb9808fe",
          9303 => x"d7387e83",
          9304 => x"11335656",
          9305 => x"74802e9f",
          9306 => x"38b01608",
          9307 => x"77315574",
          9308 => x"78279438",
          9309 => x"848053b4",
          9310 => x"1652b016",
          9311 => x"08773189",
          9312 => x"2b7d0551",
          9313 => x"cfe03f77",
          9314 => x"892b56b9",
          9315 => x"39769c1a",
          9316 => x"0c941908",
          9317 => x"83ff0684",
          9318 => x"80713157",
          9319 => x"557b7627",
          9320 => x"83387b56",
          9321 => x"9c190852",
          9322 => x"7e51d1c7",
          9323 => x"3f82bb98",
          9324 => x"08fe8138",
          9325 => x"75539419",
          9326 => x"0883ff06",
          9327 => x"1fb40552",
          9328 => x"7c51cfa2",
          9329 => x"3f7b7631",
          9330 => x"7e08177f",
          9331 => x"0c761e94",
          9332 => x"1b081894",
          9333 => x"1c0c5e5c",
          9334 => x"fdf33980",
          9335 => x"567582bb",
          9336 => x"980c903d",
          9337 => x"0d04f23d",
          9338 => x"0d606365",
          9339 => x"6440405d",
          9340 => x"58807e0c",
          9341 => x"903dfc05",
          9342 => x"527751f6",
          9343 => x"d23f82bb",
          9344 => x"98085582",
          9345 => x"bb98088a",
          9346 => x"38911833",
          9347 => x"5574802e",
          9348 => x"86387456",
          9349 => x"83b83990",
          9350 => x"18337081",
          9351 => x"2a708106",
          9352 => x"51565687",
          9353 => x"5674802e",
          9354 => x"83a43895",
          9355 => x"39820b91",
          9356 => x"19348256",
          9357 => x"83983981",
          9358 => x"0b911934",
          9359 => x"8156838e",
          9360 => x"39941808",
          9361 => x"7c115656",
          9362 => x"74762784",
          9363 => x"3875095c",
          9364 => x"7b802e82",
          9365 => x"ec389418",
          9366 => x"087083ff",
          9367 => x"06565674",
          9368 => x"81fd387e",
          9369 => x"8a1122ff",
          9370 => x"0577892a",
          9371 => x"065c557a",
          9372 => x"bf38758c",
          9373 => x"38881808",
          9374 => x"55749c38",
          9375 => x"7a528539",
          9376 => x"98180852",
          9377 => x"7751d7e7",
          9378 => x"3f82bb98",
          9379 => x"085582bb",
          9380 => x"9808802e",
          9381 => x"82ab3874",
          9382 => x"812eff91",
          9383 => x"3874ff2e",
          9384 => x"ff953874",
          9385 => x"98190c88",
          9386 => x"18088538",
          9387 => x"7488190c",
          9388 => x"7e55b015",
          9389 => x"089c1908",
          9390 => x"2e098106",
          9391 => x"8d387451",
          9392 => x"cec13f82",
          9393 => x"bb9808fe",
          9394 => x"ee389818",
          9395 => x"08527e51",
          9396 => x"d1973f82",
          9397 => x"bb980880",
          9398 => x"2efed238",
          9399 => x"82bb9808",
          9400 => x"1b7c892a",
          9401 => x"5a577880",
          9402 => x"2e80d538",
          9403 => x"781b7f8a",
          9404 => x"1122585b",
          9405 => x"55757527",
          9406 => x"8538757b",
          9407 => x"31597854",
          9408 => x"76537c52",
          9409 => x"811a3351",
          9410 => x"c8be3f82",
          9411 => x"bb9808fe",
          9412 => x"a6387eb0",
          9413 => x"11087831",
          9414 => x"56567479",
          9415 => x"279b3884",
          9416 => x"8053b016",
          9417 => x"08773189",
          9418 => x"2b7d0552",
          9419 => x"b41651cc",
          9420 => x"b53f7e55",
          9421 => x"800b8316",
          9422 => x"3478892b",
          9423 => x"5680db39",
          9424 => x"8c180894",
          9425 => x"19082693",
          9426 => x"387e51cd",
          9427 => x"b63f82bb",
          9428 => x"9808fde3",
          9429 => x"387e77b0",
          9430 => x"120c5576",
          9431 => x"9c190c94",
          9432 => x"180883ff",
          9433 => x"06848071",
          9434 => x"3157557b",
          9435 => x"76278338",
          9436 => x"7b569c18",
          9437 => x"08527e51",
          9438 => x"cdf93f82",
          9439 => x"bb9808fd",
          9440 => x"b6387553",
          9441 => x"7c529418",
          9442 => x"0883ff06",
          9443 => x"1fb40551",
          9444 => x"cbd43f7e",
          9445 => x"55810b83",
          9446 => x"16347b76",
          9447 => x"317e0817",
          9448 => x"7f0c761e",
          9449 => x"941a0818",
          9450 => x"70941c0c",
          9451 => x"8c1b0858",
          9452 => x"585e5c74",
          9453 => x"76278338",
          9454 => x"7555748c",
          9455 => x"190cfd90",
          9456 => x"39901833",
          9457 => x"80c00755",
          9458 => x"74901934",
          9459 => x"80567582",
          9460 => x"bb980c90",
          9461 => x"3d0d04f8",
          9462 => x"3d0d7a8b",
          9463 => x"3dfc0553",
          9464 => x"705256f2",
          9465 => x"ea3f82bb",
          9466 => x"98085782",
          9467 => x"bb980880",
          9468 => x"fb389016",
          9469 => x"3370862a",
          9470 => x"70810651",
          9471 => x"55557380",
          9472 => x"2e80e938",
          9473 => x"a0160852",
          9474 => x"7851cce7",
          9475 => x"3f82bb98",
          9476 => x"085782bb",
          9477 => x"980880d4",
          9478 => x"38a41608",
          9479 => x"8b1133a0",
          9480 => x"07555573",
          9481 => x"8b163488",
          9482 => x"16085374",
          9483 => x"52750851",
          9484 => x"dde83f8c",
          9485 => x"1608529c",
          9486 => x"1551c9fb",
          9487 => x"3f8288b2",
          9488 => x"0a529615",
          9489 => x"51c9f03f",
          9490 => x"76529215",
          9491 => x"51c9ca3f",
          9492 => x"7854810b",
          9493 => x"83153478",
          9494 => x"51ccdf3f",
          9495 => x"82bb9808",
          9496 => x"90173381",
          9497 => x"bf065557",
          9498 => x"73901734",
          9499 => x"7682bb98",
          9500 => x"0c8a3d0d",
          9501 => x"04fc3d0d",
          9502 => x"76705254",
          9503 => x"fed93f82",
          9504 => x"bb980853",
          9505 => x"82bb9808",
          9506 => x"9c38863d",
          9507 => x"fc055273",
          9508 => x"51f1bc3f",
          9509 => x"82bb9808",
          9510 => x"5382bb98",
          9511 => x"08873882",
          9512 => x"bb980874",
          9513 => x"0c7282bb",
          9514 => x"980c863d",
          9515 => x"0d04ff3d",
          9516 => x"0d843d51",
          9517 => x"e6e43f8b",
          9518 => x"52800b82",
          9519 => x"bb980824",
          9520 => x"8b3882bb",
          9521 => x"980882d2",
          9522 => x"e4348052",
          9523 => x"7182bb98",
          9524 => x"0c833d0d",
          9525 => x"04ef3d0d",
          9526 => x"8053933d",
          9527 => x"d0055294",
          9528 => x"3d51e9c1",
          9529 => x"3f82bb98",
          9530 => x"085582bb",
          9531 => x"980880e0",
          9532 => x"38765863",
          9533 => x"52933dd4",
          9534 => x"0551e08d",
          9535 => x"3f82bb98",
          9536 => x"085582bb",
          9537 => x"9808bc38",
          9538 => x"0280c705",
          9539 => x"3370982b",
          9540 => x"55567380",
          9541 => x"25893876",
          9542 => x"7a94120c",
          9543 => x"54b23902",
          9544 => x"a2053370",
          9545 => x"842a7081",
          9546 => x"06515556",
          9547 => x"73802e9e",
          9548 => x"38767f53",
          9549 => x"705254db",
          9550 => x"a83f82bb",
          9551 => x"98089415",
          9552 => x"0c8e3982",
          9553 => x"bb980884",
          9554 => x"2e098106",
          9555 => x"83388555",
          9556 => x"7482bb98",
          9557 => x"0c933d0d",
          9558 => x"04e43d0d",
          9559 => x"6f6f5b5b",
          9560 => x"807a3480",
          9561 => x"539e3dff",
          9562 => x"b805529f",
          9563 => x"3d51e8b5",
          9564 => x"3f82bb98",
          9565 => x"085782bb",
          9566 => x"980882fc",
          9567 => x"387b437a",
          9568 => x"7c941108",
          9569 => x"47555864",
          9570 => x"5473802e",
          9571 => x"81ed38a0",
          9572 => x"52933d70",
          9573 => x"5255d5ea",
          9574 => x"3f82bb98",
          9575 => x"085782bb",
          9576 => x"980882d4",
          9577 => x"3868527b",
          9578 => x"51c9c83f",
          9579 => x"82bb9808",
          9580 => x"5782bb98",
          9581 => x"0882c138",
          9582 => x"69527b51",
          9583 => x"daa33f82",
          9584 => x"bb980845",
          9585 => x"76527451",
          9586 => x"d5b83f82",
          9587 => x"bb980857",
          9588 => x"82bb9808",
          9589 => x"82a23880",
          9590 => x"527451da",
          9591 => x"eb3f82bb",
          9592 => x"98085782",
          9593 => x"bb9808a4",
          9594 => x"3869527b",
          9595 => x"51d9f23f",
          9596 => x"7382bb98",
          9597 => x"082ea638",
          9598 => x"76527451",
          9599 => x"d6cf3f82",
          9600 => x"bb980857",
          9601 => x"82bb9808",
          9602 => x"802ecc38",
          9603 => x"76842e09",
          9604 => x"81068638",
          9605 => x"825781e0",
          9606 => x"397681dc",
          9607 => x"389e3dff",
          9608 => x"bc055274",
          9609 => x"51dcc93f",
          9610 => x"76903d78",
          9611 => x"11811133",
          9612 => x"51565a56",
          9613 => x"73802e91",
          9614 => x"3802b905",
          9615 => x"55811681",
          9616 => x"16703356",
          9617 => x"565673f5",
          9618 => x"38811654",
          9619 => x"73782681",
          9620 => x"90387580",
          9621 => x"2e993878",
          9622 => x"16810555",
          9623 => x"ff186f11",
          9624 => x"ff18ff18",
          9625 => x"58585558",
          9626 => x"74337434",
          9627 => x"75ee38ff",
          9628 => x"186f1155",
          9629 => x"58af7434",
          9630 => x"fe8d3977",
          9631 => x"7b2e0981",
          9632 => x"068a38ff",
          9633 => x"186f1155",
          9634 => x"58af7434",
          9635 => x"800b82d2",
          9636 => x"e4337084",
          9637 => x"2982b4d0",
          9638 => x"05700870",
          9639 => x"33525c56",
          9640 => x"56567376",
          9641 => x"2e8d3881",
          9642 => x"16701a70",
          9643 => x"33515556",
          9644 => x"73f53882",
          9645 => x"16547378",
          9646 => x"26a73880",
          9647 => x"55747627",
          9648 => x"91387419",
          9649 => x"5473337a",
          9650 => x"7081055c",
          9651 => x"34811555",
          9652 => x"ec39ba7a",
          9653 => x"7081055c",
          9654 => x"3474ff2e",
          9655 => x"09810685",
          9656 => x"38915794",
          9657 => x"396e1881",
          9658 => x"19595473",
          9659 => x"337a7081",
          9660 => x"055c347a",
          9661 => x"7826ee38",
          9662 => x"807a3476",
          9663 => x"82bb980c",
          9664 => x"9e3d0d04",
          9665 => x"f73d0d7b",
          9666 => x"7d8d3dfc",
          9667 => x"05547153",
          9668 => x"5755ecbb",
          9669 => x"3f82bb98",
          9670 => x"085382bb",
          9671 => x"980882fa",
          9672 => x"38911533",
          9673 => x"537282f2",
          9674 => x"388c1508",
          9675 => x"54737627",
          9676 => x"92389015",
          9677 => x"3370812a",
          9678 => x"70810651",
          9679 => x"54577283",
          9680 => x"38735694",
          9681 => x"15085480",
          9682 => x"7094170c",
          9683 => x"5875782e",
          9684 => x"82973879",
          9685 => x"8a112270",
          9686 => x"892b5951",
          9687 => x"5373782e",
          9688 => x"b7387652",
          9689 => x"ff1651fe",
          9690 => x"e3b93f82",
          9691 => x"bb9808ff",
          9692 => x"15785470",
          9693 => x"535553fe",
          9694 => x"e3a93f82",
          9695 => x"bb980873",
          9696 => x"26963876",
          9697 => x"30707506",
          9698 => x"7094180c",
          9699 => x"77713198",
          9700 => x"18085758",
          9701 => x"5153b139",
          9702 => x"88150854",
          9703 => x"73a63873",
          9704 => x"527451cd",
          9705 => x"ca3f82bb",
          9706 => x"98085482",
          9707 => x"bb980881",
          9708 => x"2e819a38",
          9709 => x"82bb9808",
          9710 => x"ff2e819b",
          9711 => x"3882bb98",
          9712 => x"0888160c",
          9713 => x"7398160c",
          9714 => x"73802e81",
          9715 => x"9c387676",
          9716 => x"2780dc38",
          9717 => x"75773194",
          9718 => x"16081894",
          9719 => x"170c9016",
          9720 => x"3370812a",
          9721 => x"70810651",
          9722 => x"555a5672",
          9723 => x"802e9a38",
          9724 => x"73527451",
          9725 => x"ccf93f82",
          9726 => x"bb980854",
          9727 => x"82bb9808",
          9728 => x"943882bb",
          9729 => x"980856a7",
          9730 => x"39735274",
          9731 => x"51c7843f",
          9732 => x"82bb9808",
          9733 => x"5473ff2e",
          9734 => x"be388174",
          9735 => x"27af3879",
          9736 => x"53739814",
          9737 => x"0827a638",
          9738 => x"7398160c",
          9739 => x"ffa03994",
          9740 => x"15081694",
          9741 => x"160c7583",
          9742 => x"ff065372",
          9743 => x"802eaa38",
          9744 => x"73527951",
          9745 => x"c6a33f82",
          9746 => x"bb980894",
          9747 => x"38820b91",
          9748 => x"16348253",
          9749 => x"80c43981",
          9750 => x"0b911634",
          9751 => x"8153bb39",
          9752 => x"75892a82",
          9753 => x"bb980805",
          9754 => x"58941508",
          9755 => x"548c1508",
          9756 => x"74279038",
          9757 => x"738c160c",
          9758 => x"90153380",
          9759 => x"c0075372",
          9760 => x"90163473",
          9761 => x"83ff0653",
          9762 => x"72802e8c",
          9763 => x"38779c16",
          9764 => x"082e8538",
          9765 => x"779c160c",
          9766 => x"80537282",
          9767 => x"bb980c8b",
          9768 => x"3d0d04f9",
          9769 => x"3d0d7956",
          9770 => x"89547580",
          9771 => x"2e818a38",
          9772 => x"8053893d",
          9773 => x"fc05528a",
          9774 => x"3d840551",
          9775 => x"e1e73f82",
          9776 => x"bb980855",
          9777 => x"82bb9808",
          9778 => x"80ea3877",
          9779 => x"760c7a52",
          9780 => x"7551d8b5",
          9781 => x"3f82bb98",
          9782 => x"085582bb",
          9783 => x"980880c3",
          9784 => x"38ab1633",
          9785 => x"70982b55",
          9786 => x"57807424",
          9787 => x"a2388616",
          9788 => x"3370842a",
          9789 => x"70810651",
          9790 => x"55577380",
          9791 => x"2ead389c",
          9792 => x"16085277",
          9793 => x"51d3da3f",
          9794 => x"82bb9808",
          9795 => x"88170c77",
          9796 => x"54861422",
          9797 => x"84172374",
          9798 => x"527551ce",
          9799 => x"e53f82bb",
          9800 => x"98085574",
          9801 => x"842e0981",
          9802 => x"06853885",
          9803 => x"55863974",
          9804 => x"802e8438",
          9805 => x"80760c74",
          9806 => x"547382bb",
          9807 => x"980c893d",
          9808 => x"0d04fc3d",
          9809 => x"0d76873d",
          9810 => x"fc055370",
          9811 => x"5253e7ff",
          9812 => x"3f82bb98",
          9813 => x"08873882",
          9814 => x"bb980873",
          9815 => x"0c863d0d",
          9816 => x"04fb3d0d",
          9817 => x"7779893d",
          9818 => x"fc055471",
          9819 => x"535654e7",
          9820 => x"de3f82bb",
          9821 => x"98085382",
          9822 => x"bb980880",
          9823 => x"df387493",
          9824 => x"3882bb98",
          9825 => x"08527351",
          9826 => x"cdf83f82",
          9827 => x"bb980853",
          9828 => x"80ca3982",
          9829 => x"bb980852",
          9830 => x"7351d3ac",
          9831 => x"3f82bb98",
          9832 => x"085382bb",
          9833 => x"9808842e",
          9834 => x"09810685",
          9835 => x"38805387",
          9836 => x"3982bb98",
          9837 => x"08a63874",
          9838 => x"527351d5",
          9839 => x"b33f7252",
          9840 => x"7351cf89",
          9841 => x"3f82bb98",
          9842 => x"08843270",
          9843 => x"30707207",
          9844 => x"9f2c7082",
          9845 => x"bb980806",
          9846 => x"51515454",
          9847 => x"7282bb98",
          9848 => x"0c873d0d",
          9849 => x"04ee3d0d",
          9850 => x"65578053",
          9851 => x"893d7053",
          9852 => x"963d5256",
          9853 => x"dfaf3f82",
          9854 => x"bb980855",
          9855 => x"82bb9808",
          9856 => x"b2386452",
          9857 => x"7551d681",
          9858 => x"3f82bb98",
          9859 => x"085582bb",
          9860 => x"9808a038",
          9861 => x"0280cb05",
          9862 => x"3370982b",
          9863 => x"55587380",
          9864 => x"25853886",
          9865 => x"558d3976",
          9866 => x"802e8838",
          9867 => x"76527551",
          9868 => x"d4be3f74",
          9869 => x"82bb980c",
          9870 => x"943d0d04",
          9871 => x"f03d0d63",
          9872 => x"65555c80",
          9873 => x"53923dec",
          9874 => x"0552933d",
          9875 => x"51ded63f",
          9876 => x"82bb9808",
          9877 => x"5b82bb98",
          9878 => x"08828038",
          9879 => x"7c740c73",
          9880 => x"08981108",
          9881 => x"fe119013",
          9882 => x"08595658",
          9883 => x"55757426",
          9884 => x"9138757c",
          9885 => x"0c81e439",
          9886 => x"815b81cc",
          9887 => x"39825b81",
          9888 => x"c73982bb",
          9889 => x"98087533",
          9890 => x"55597381",
          9891 => x"2e098106",
          9892 => x"bf388275",
          9893 => x"5f577652",
          9894 => x"923df005",
          9895 => x"51c1f43f",
          9896 => x"82bb9808",
          9897 => x"ff2ed138",
          9898 => x"82bb9808",
          9899 => x"812ece38",
          9900 => x"82bb9808",
          9901 => x"307082bb",
          9902 => x"98080780",
          9903 => x"257a0581",
          9904 => x"197f5359",
          9905 => x"5a549814",
          9906 => x"087726ca",
          9907 => x"3880f939",
          9908 => x"a4150882",
          9909 => x"bb980857",
          9910 => x"58759838",
          9911 => x"77528118",
          9912 => x"7d5258ff",
          9913 => x"bf8d3f82",
          9914 => x"bb98085b",
          9915 => x"82bb9808",
          9916 => x"80d6387c",
          9917 => x"70337712",
          9918 => x"ff1a5d52",
          9919 => x"56547482",
          9920 => x"2e098106",
          9921 => x"9e38b414",
          9922 => x"51ffbbcb",
          9923 => x"3f82bb98",
          9924 => x"0883ffff",
          9925 => x"06703070",
          9926 => x"80251b82",
          9927 => x"19595b51",
          9928 => x"549b39b4",
          9929 => x"1451ffbb",
          9930 => x"c53f82bb",
          9931 => x"9808f00a",
          9932 => x"06703070",
          9933 => x"80251b84",
          9934 => x"19595b51",
          9935 => x"547583ff",
          9936 => x"067a5856",
          9937 => x"79ff9238",
          9938 => x"787c0c7c",
          9939 => x"7990120c",
          9940 => x"84113381",
          9941 => x"07565474",
          9942 => x"8415347a",
          9943 => x"82bb980c",
          9944 => x"923d0d04",
          9945 => x"f93d0d79",
          9946 => x"8a3dfc05",
          9947 => x"53705257",
          9948 => x"e3dd3f82",
          9949 => x"bb980856",
          9950 => x"82bb9808",
          9951 => x"81a83891",
          9952 => x"17335675",
          9953 => x"81a03890",
          9954 => x"17337081",
          9955 => x"2a708106",
          9956 => x"51555587",
          9957 => x"5573802e",
          9958 => x"818e3894",
          9959 => x"17085473",
          9960 => x"8c180827",
          9961 => x"81803873",
          9962 => x"9b3882bb",
          9963 => x"98085388",
          9964 => x"17085276",
          9965 => x"51c48c3f",
          9966 => x"82bb9808",
          9967 => x"7488190c",
          9968 => x"5680c939",
          9969 => x"98170852",
          9970 => x"7651ffbf",
          9971 => x"c63f82bb",
          9972 => x"9808ff2e",
          9973 => x"09810683",
          9974 => x"38815682",
          9975 => x"bb980881",
          9976 => x"2e098106",
          9977 => x"85388256",
          9978 => x"a33975a0",
          9979 => x"38775482",
          9980 => x"bb980898",
          9981 => x"15082794",
          9982 => x"38981708",
          9983 => x"5382bb98",
          9984 => x"08527651",
          9985 => x"c3bd3f82",
          9986 => x"bb980856",
          9987 => x"9417088c",
          9988 => x"180c9017",
          9989 => x"3380c007",
          9990 => x"54739018",
          9991 => x"3475802e",
          9992 => x"85387591",
          9993 => x"18347555",
          9994 => x"7482bb98",
          9995 => x"0c893d0d",
          9996 => x"04e23d0d",
          9997 => x"8253a03d",
          9998 => x"ffa40552",
          9999 => x"a13d51da",
         10000 => x"e43f82bb",
         10001 => x"98085582",
         10002 => x"bb980881",
         10003 => x"f5387845",
         10004 => x"a13d0852",
         10005 => x"953d7052",
         10006 => x"58d1ae3f",
         10007 => x"82bb9808",
         10008 => x"5582bb98",
         10009 => x"0881db38",
         10010 => x"0280fb05",
         10011 => x"3370852a",
         10012 => x"70810651",
         10013 => x"55568655",
         10014 => x"7381c738",
         10015 => x"75982b54",
         10016 => x"80742481",
         10017 => x"bd380280",
         10018 => x"d6053370",
         10019 => x"81065854",
         10020 => x"87557681",
         10021 => x"ad386b52",
         10022 => x"7851ccc5",
         10023 => x"3f82bb98",
         10024 => x"0874842a",
         10025 => x"70810651",
         10026 => x"55567380",
         10027 => x"2e80d438",
         10028 => x"785482bb",
         10029 => x"98089415",
         10030 => x"082e8186",
         10031 => x"38735a82",
         10032 => x"bb98085c",
         10033 => x"76528a3d",
         10034 => x"705254c7",
         10035 => x"b53f82bb",
         10036 => x"98085582",
         10037 => x"bb980880",
         10038 => x"e93882bb",
         10039 => x"98085273",
         10040 => x"51cce53f",
         10041 => x"82bb9808",
         10042 => x"5582bb98",
         10043 => x"08863887",
         10044 => x"5580cf39",
         10045 => x"82bb9808",
         10046 => x"842e8838",
         10047 => x"82bb9808",
         10048 => x"80c03877",
         10049 => x"51cec23f",
         10050 => x"82bb9808",
         10051 => x"82bb9808",
         10052 => x"307082bb",
         10053 => x"98080780",
         10054 => x"25515555",
         10055 => x"75802e94",
         10056 => x"3873802e",
         10057 => x"8f388053",
         10058 => x"75527751",
         10059 => x"c1953f82",
         10060 => x"bb980855",
         10061 => x"748c3878",
         10062 => x"51ffbafe",
         10063 => x"3f82bb98",
         10064 => x"08557482",
         10065 => x"bb980ca0",
         10066 => x"3d0d04e9",
         10067 => x"3d0d8253",
         10068 => x"993dc005",
         10069 => x"529a3d51",
         10070 => x"d8cb3f82",
         10071 => x"bb980854",
         10072 => x"82bb9808",
         10073 => x"82b03878",
         10074 => x"5e69528e",
         10075 => x"3d705258",
         10076 => x"cf973f82",
         10077 => x"bb980854",
         10078 => x"82bb9808",
         10079 => x"86388854",
         10080 => x"82943982",
         10081 => x"bb980884",
         10082 => x"2e098106",
         10083 => x"82883802",
         10084 => x"80df0533",
         10085 => x"70852a81",
         10086 => x"06515586",
         10087 => x"547481f6",
         10088 => x"38785a74",
         10089 => x"528a3d70",
         10090 => x"5257c1c3",
         10091 => x"3f82bb98",
         10092 => x"08755556",
         10093 => x"82bb9808",
         10094 => x"83388754",
         10095 => x"82bb9808",
         10096 => x"812e0981",
         10097 => x"06833882",
         10098 => x"5482bb98",
         10099 => x"08ff2e09",
         10100 => x"81068638",
         10101 => x"815481b4",
         10102 => x"397381b0",
         10103 => x"3882bb98",
         10104 => x"08527851",
         10105 => x"c4a43f82",
         10106 => x"bb980854",
         10107 => x"82bb9808",
         10108 => x"819a388b",
         10109 => x"53a052b4",
         10110 => x"1951ffb7",
         10111 => x"8c3f7854",
         10112 => x"ae0bb415",
         10113 => x"34785490",
         10114 => x"0bbf1534",
         10115 => x"8288b20a",
         10116 => x"5280ca19",
         10117 => x"51ffb69f",
         10118 => x"3f755378",
         10119 => x"b4115351",
         10120 => x"c9f83fa0",
         10121 => x"5378b411",
         10122 => x"5380d405",
         10123 => x"51ffb6b6",
         10124 => x"3f7854ae",
         10125 => x"0b80d515",
         10126 => x"347f5378",
         10127 => x"80d41153",
         10128 => x"51c9d73f",
         10129 => x"7854810b",
         10130 => x"83153477",
         10131 => x"51cba43f",
         10132 => x"82bb9808",
         10133 => x"5482bb98",
         10134 => x"08b23882",
         10135 => x"88b20a52",
         10136 => x"64960551",
         10137 => x"ffb5d03f",
         10138 => x"75536452",
         10139 => x"7851c9aa",
         10140 => x"3f645490",
         10141 => x"0b8b1534",
         10142 => x"7854810b",
         10143 => x"83153478",
         10144 => x"51ffb8b6",
         10145 => x"3f82bb98",
         10146 => x"08548b39",
         10147 => x"80537552",
         10148 => x"7651ffbe",
         10149 => x"ae3f7382",
         10150 => x"bb980c99",
         10151 => x"3d0d04da",
         10152 => x"3d0da93d",
         10153 => x"840551d2",
         10154 => x"f13f8253",
         10155 => x"a83dff84",
         10156 => x"0552a93d",
         10157 => x"51d5ee3f",
         10158 => x"82bb9808",
         10159 => x"5582bb98",
         10160 => x"0882d338",
         10161 => x"784da93d",
         10162 => x"08529d3d",
         10163 => x"705258cc",
         10164 => x"b83f82bb",
         10165 => x"98085582",
         10166 => x"bb980882",
         10167 => x"b9380281",
         10168 => x"9b053381",
         10169 => x"a0065486",
         10170 => x"557382aa",
         10171 => x"38a053a4",
         10172 => x"3d0852a8",
         10173 => x"3dff8805",
         10174 => x"51ffb4ea",
         10175 => x"3fac5377",
         10176 => x"52923d70",
         10177 => x"5254ffb4",
         10178 => x"dd3faa3d",
         10179 => x"08527351",
         10180 => x"cbf73f82",
         10181 => x"bb980855",
         10182 => x"82bb9808",
         10183 => x"9538636f",
         10184 => x"2e098106",
         10185 => x"883865a2",
         10186 => x"3d082e92",
         10187 => x"38885581",
         10188 => x"e53982bb",
         10189 => x"9808842e",
         10190 => x"09810681",
         10191 => x"b8387351",
         10192 => x"c9b13f82",
         10193 => x"bb980855",
         10194 => x"82bb9808",
         10195 => x"81c83868",
         10196 => x"569353a8",
         10197 => x"3dff9505",
         10198 => x"528d1651",
         10199 => x"ffb4873f",
         10200 => x"02af0533",
         10201 => x"8b17348b",
         10202 => x"16337084",
         10203 => x"2a708106",
         10204 => x"51555573",
         10205 => x"893874a0",
         10206 => x"0754738b",
         10207 => x"17347854",
         10208 => x"810b8315",
         10209 => x"348b1633",
         10210 => x"70842a70",
         10211 => x"81065155",
         10212 => x"5573802e",
         10213 => x"80e5386e",
         10214 => x"642e80df",
         10215 => x"38755278",
         10216 => x"51c6be3f",
         10217 => x"82bb9808",
         10218 => x"527851ff",
         10219 => x"b7bb3f82",
         10220 => x"5582bb98",
         10221 => x"08802e80",
         10222 => x"dd3882bb",
         10223 => x"98085278",
         10224 => x"51ffb5af",
         10225 => x"3f82bb98",
         10226 => x"087980d4",
         10227 => x"11585855",
         10228 => x"82bb9808",
         10229 => x"80c03881",
         10230 => x"16335473",
         10231 => x"ae2e0981",
         10232 => x"06993863",
         10233 => x"53755276",
         10234 => x"51c6af3f",
         10235 => x"7854810b",
         10236 => x"83153487",
         10237 => x"3982bb98",
         10238 => x"089c3877",
         10239 => x"51c8ca3f",
         10240 => x"82bb9808",
         10241 => x"5582bb98",
         10242 => x"088c3878",
         10243 => x"51ffb5aa",
         10244 => x"3f82bb98",
         10245 => x"08557482",
         10246 => x"bb980ca8",
         10247 => x"3d0d04ed",
         10248 => x"3d0d0280",
         10249 => x"db053302",
         10250 => x"840580df",
         10251 => x"05335757",
         10252 => x"8253953d",
         10253 => x"d0055296",
         10254 => x"3d51d2e9",
         10255 => x"3f82bb98",
         10256 => x"085582bb",
         10257 => x"980880cf",
         10258 => x"38785a65",
         10259 => x"52953dd4",
         10260 => x"0551c9b5",
         10261 => x"3f82bb98",
         10262 => x"085582bb",
         10263 => x"9808b838",
         10264 => x"0280cf05",
         10265 => x"3381a006",
         10266 => x"54865573",
         10267 => x"aa3875a7",
         10268 => x"06617109",
         10269 => x"8b123371",
         10270 => x"067a7406",
         10271 => x"07515755",
         10272 => x"56748b15",
         10273 => x"34785481",
         10274 => x"0b831534",
         10275 => x"7851ffb4",
         10276 => x"a93f82bb",
         10277 => x"98085574",
         10278 => x"82bb980c",
         10279 => x"953d0d04",
         10280 => x"ef3d0d64",
         10281 => x"56825393",
         10282 => x"3dd00552",
         10283 => x"943d51d1",
         10284 => x"f43f82bb",
         10285 => x"98085582",
         10286 => x"bb980880",
         10287 => x"cb387658",
         10288 => x"6352933d",
         10289 => x"d40551c8",
         10290 => x"c03f82bb",
         10291 => x"98085582",
         10292 => x"bb9808b4",
         10293 => x"380280c7",
         10294 => x"053381a0",
         10295 => x"06548655",
         10296 => x"73a63884",
         10297 => x"16228617",
         10298 => x"2271902b",
         10299 => x"07535496",
         10300 => x"1f51ffb0",
         10301 => x"c23f7654",
         10302 => x"810b8315",
         10303 => x"347651ff",
         10304 => x"b3b83f82",
         10305 => x"bb980855",
         10306 => x"7482bb98",
         10307 => x"0c933d0d",
         10308 => x"04ea3d0d",
         10309 => x"696b5c5a",
         10310 => x"8053983d",
         10311 => x"d0055299",
         10312 => x"3d51d181",
         10313 => x"3f82bb98",
         10314 => x"0882bb98",
         10315 => x"08307082",
         10316 => x"bb980807",
         10317 => x"80255155",
         10318 => x"5779802e",
         10319 => x"81853881",
         10320 => x"70750655",
         10321 => x"5573802e",
         10322 => x"80f9387b",
         10323 => x"5d805f80",
         10324 => x"528d3d70",
         10325 => x"5254ffbe",
         10326 => x"a93f82bb",
         10327 => x"98085782",
         10328 => x"bb980880",
         10329 => x"d1387452",
         10330 => x"7351c3dc",
         10331 => x"3f82bb98",
         10332 => x"085782bb",
         10333 => x"9808bf38",
         10334 => x"82bb9808",
         10335 => x"82bb9808",
         10336 => x"655b5956",
         10337 => x"78188119",
         10338 => x"7b185659",
         10339 => x"55743374",
         10340 => x"34811656",
         10341 => x"8a7827ec",
         10342 => x"388b5675",
         10343 => x"1a548074",
         10344 => x"3475802e",
         10345 => x"9e38ff16",
         10346 => x"701b7033",
         10347 => x"51555673",
         10348 => x"a02ee838",
         10349 => x"8e397684",
         10350 => x"2e098106",
         10351 => x"8638807a",
         10352 => x"34805776",
         10353 => x"30707807",
         10354 => x"80255154",
         10355 => x"7a802e80",
         10356 => x"c1387380",
         10357 => x"2ebc387b",
         10358 => x"a0110853",
         10359 => x"51ffb193",
         10360 => x"3f82bb98",
         10361 => x"085782bb",
         10362 => x"9808a738",
         10363 => x"7b703355",
         10364 => x"5580c356",
         10365 => x"73832e8b",
         10366 => x"3880e456",
         10367 => x"73842e83",
         10368 => x"38a75675",
         10369 => x"15b40551",
         10370 => x"ffade33f",
         10371 => x"82bb9808",
         10372 => x"7b0c7682",
         10373 => x"bb980c98",
         10374 => x"3d0d04e6",
         10375 => x"3d0d8253",
         10376 => x"9c3dffb8",
         10377 => x"05529d3d",
         10378 => x"51cefa3f",
         10379 => x"82bb9808",
         10380 => x"82bb9808",
         10381 => x"565482bb",
         10382 => x"98088398",
         10383 => x"388b53a0",
         10384 => x"528b3d70",
         10385 => x"5259ffae",
         10386 => x"c03f736d",
         10387 => x"70337081",
         10388 => x"ff065257",
         10389 => x"55579f74",
         10390 => x"2781bc38",
         10391 => x"78587481",
         10392 => x"ff066d81",
         10393 => x"054e7052",
         10394 => x"55ffaf89",
         10395 => x"3f82bb98",
         10396 => x"08802ea5",
         10397 => x"386c7033",
         10398 => x"70535754",
         10399 => x"ffaefd3f",
         10400 => x"82bb9808",
         10401 => x"802e8d38",
         10402 => x"74882b76",
         10403 => x"076d8105",
         10404 => x"4e558639",
         10405 => x"82bb9808",
         10406 => x"55ff9f15",
         10407 => x"7083ffff",
         10408 => x"06515473",
         10409 => x"99268a38",
         10410 => x"e0157083",
         10411 => x"ffff0656",
         10412 => x"5480ff75",
         10413 => x"27873882",
         10414 => x"b3e01533",
         10415 => x"5574802e",
         10416 => x"a3387452",
         10417 => x"82b5e051",
         10418 => x"ffae893f",
         10419 => x"82bb9808",
         10420 => x"933881ff",
         10421 => x"75278838",
         10422 => x"76892688",
         10423 => x"388b398a",
         10424 => x"77278638",
         10425 => x"865581ec",
         10426 => x"3981ff75",
         10427 => x"278f3874",
         10428 => x"882a5473",
         10429 => x"78708105",
         10430 => x"5a348117",
         10431 => x"57747870",
         10432 => x"81055a34",
         10433 => x"81176d70",
         10434 => x"337081ff",
         10435 => x"06525755",
         10436 => x"57739f26",
         10437 => x"fec8388b",
         10438 => x"3d335486",
         10439 => x"557381e5",
         10440 => x"2e81b138",
         10441 => x"76802e99",
         10442 => x"3802a705",
         10443 => x"55761570",
         10444 => x"33515473",
         10445 => x"a02e0981",
         10446 => x"068738ff",
         10447 => x"175776ed",
         10448 => x"38794180",
         10449 => x"43805291",
         10450 => x"3d705255",
         10451 => x"ffbab33f",
         10452 => x"82bb9808",
         10453 => x"5482bb98",
         10454 => x"0880f738",
         10455 => x"81527451",
         10456 => x"ffbfe53f",
         10457 => x"82bb9808",
         10458 => x"5482bb98",
         10459 => x"088d3876",
         10460 => x"80c43867",
         10461 => x"54e57434",
         10462 => x"80c63982",
         10463 => x"bb980884",
         10464 => x"2e098106",
         10465 => x"80cc3880",
         10466 => x"5476742e",
         10467 => x"80c43881",
         10468 => x"527451ff",
         10469 => x"bdb03f82",
         10470 => x"bb980854",
         10471 => x"82bb9808",
         10472 => x"b138a053",
         10473 => x"82bb9808",
         10474 => x"526751ff",
         10475 => x"abdb3f67",
         10476 => x"54880b8b",
         10477 => x"15348b53",
         10478 => x"78526751",
         10479 => x"ffaba73f",
         10480 => x"7954810b",
         10481 => x"83153479",
         10482 => x"51ffadee",
         10483 => x"3f82bb98",
         10484 => x"08547355",
         10485 => x"7482bb98",
         10486 => x"0c9c3d0d",
         10487 => x"04f23d0d",
         10488 => x"60620288",
         10489 => x"0580cb05",
         10490 => x"33933dfc",
         10491 => x"05557254",
         10492 => x"405e5ad2",
         10493 => x"da3f82bb",
         10494 => x"98085882",
         10495 => x"bb980882",
         10496 => x"bd38911a",
         10497 => x"33587782",
         10498 => x"b5387c80",
         10499 => x"2e97388c",
         10500 => x"1a085978",
         10501 => x"9038901a",
         10502 => x"3370812a",
         10503 => x"70810651",
         10504 => x"55557390",
         10505 => x"38875482",
         10506 => x"97398258",
         10507 => x"82903981",
         10508 => x"58828b39",
         10509 => x"7e8a1122",
         10510 => x"70892b70",
         10511 => x"557f5456",
         10512 => x"5656fec9",
         10513 => x"de3fff14",
         10514 => x"7d067030",
         10515 => x"7072079f",
         10516 => x"2a82bb98",
         10517 => x"08058c19",
         10518 => x"087c405a",
         10519 => x"5d555581",
         10520 => x"77278838",
         10521 => x"98160877",
         10522 => x"26833882",
         10523 => x"57767756",
         10524 => x"59805674",
         10525 => x"527951ff",
         10526 => x"ae993f81",
         10527 => x"157f5555",
         10528 => x"98140875",
         10529 => x"26833882",
         10530 => x"5582bb98",
         10531 => x"08812eff",
         10532 => x"993882bb",
         10533 => x"9808ff2e",
         10534 => x"ff953882",
         10535 => x"bb98088e",
         10536 => x"38811656",
         10537 => x"757b2e09",
         10538 => x"81068738",
         10539 => x"93397459",
         10540 => x"80567477",
         10541 => x"2e098106",
         10542 => x"ffb93887",
         10543 => x"5880ff39",
         10544 => x"7d802eba",
         10545 => x"38787b55",
         10546 => x"557a802e",
         10547 => x"b4388115",
         10548 => x"5673812e",
         10549 => x"09810683",
         10550 => x"38ff5675",
         10551 => x"5374527e",
         10552 => x"51ffafa8",
         10553 => x"3f82bb98",
         10554 => x"085882bb",
         10555 => x"980880ce",
         10556 => x"38748116",
         10557 => x"ff165656",
         10558 => x"5c73d338",
         10559 => x"8439ff19",
         10560 => x"5c7e7c8c",
         10561 => x"120c557d",
         10562 => x"802eb338",
         10563 => x"78881b0c",
         10564 => x"7c8c1b0c",
         10565 => x"901a3380",
         10566 => x"c0075473",
         10567 => x"901b3498",
         10568 => x"1508fe05",
         10569 => x"90160857",
         10570 => x"54757426",
         10571 => x"9138757b",
         10572 => x"3190160c",
         10573 => x"84153381",
         10574 => x"07547384",
         10575 => x"16347754",
         10576 => x"7382bb98",
         10577 => x"0c903d0d",
         10578 => x"04e93d0d",
         10579 => x"6b6d0288",
         10580 => x"0580eb05",
         10581 => x"339d3d54",
         10582 => x"5a5c59c5",
         10583 => x"bd3f8b56",
         10584 => x"800b82bb",
         10585 => x"9808248b",
         10586 => x"f83882bb",
         10587 => x"98088429",
         10588 => x"82d2d005",
         10589 => x"70085155",
         10590 => x"74802e84",
         10591 => x"38807534",
         10592 => x"82bb9808",
         10593 => x"81ff065f",
         10594 => x"81527e51",
         10595 => x"ffa0d03f",
         10596 => x"82bb9808",
         10597 => x"81ff0670",
         10598 => x"81065657",
         10599 => x"8356748b",
         10600 => x"c0387682",
         10601 => x"2a708106",
         10602 => x"51558a56",
         10603 => x"748bb238",
         10604 => x"993dfc05",
         10605 => x"5383527e",
         10606 => x"51ffa4f0",
         10607 => x"3f82bb98",
         10608 => x"08993867",
         10609 => x"5574802e",
         10610 => x"92387482",
         10611 => x"8080268b",
         10612 => x"38ff1575",
         10613 => x"06557480",
         10614 => x"2e833881",
         10615 => x"4878802e",
         10616 => x"87388480",
         10617 => x"79269238",
         10618 => x"7881800a",
         10619 => x"268b38ff",
         10620 => x"19790655",
         10621 => x"74802e86",
         10622 => x"3893568a",
         10623 => x"e4397889",
         10624 => x"2a6e892a",
         10625 => x"70892b77",
         10626 => x"59484359",
         10627 => x"7a833881",
         10628 => x"56613070",
         10629 => x"80257707",
         10630 => x"51559156",
         10631 => x"748ac238",
         10632 => x"993df805",
         10633 => x"5381527e",
         10634 => x"51ffa480",
         10635 => x"3f815682",
         10636 => x"bb98088a",
         10637 => x"ac387783",
         10638 => x"2a707706",
         10639 => x"82bb9808",
         10640 => x"43564574",
         10641 => x"8338bf41",
         10642 => x"66558e56",
         10643 => x"6075268a",
         10644 => x"90387461",
         10645 => x"31704855",
         10646 => x"80ff7527",
         10647 => x"8a833893",
         10648 => x"56788180",
         10649 => x"2689fa38",
         10650 => x"77812a70",
         10651 => x"81065643",
         10652 => x"74802e95",
         10653 => x"38778706",
         10654 => x"5574822e",
         10655 => x"838d3877",
         10656 => x"81065574",
         10657 => x"802e8383",
         10658 => x"38778106",
         10659 => x"55935682",
         10660 => x"5e74802e",
         10661 => x"89cb3878",
         10662 => x"5a7d832e",
         10663 => x"09810680",
         10664 => x"e13878ae",
         10665 => x"3866912a",
         10666 => x"57810b82",
         10667 => x"b6842256",
         10668 => x"5a74802e",
         10669 => x"9d387477",
         10670 => x"26983882",
         10671 => x"b6845679",
         10672 => x"10821770",
         10673 => x"2257575a",
         10674 => x"74802e86",
         10675 => x"38767527",
         10676 => x"ee387952",
         10677 => x"6651fec4",
         10678 => x"ca3f82bb",
         10679 => x"98088429",
         10680 => x"84870570",
         10681 => x"892a5e55",
         10682 => x"a05c800b",
         10683 => x"82bb9808",
         10684 => x"fc808a05",
         10685 => x"5644fdff",
         10686 => x"f00a7527",
         10687 => x"80ec3888",
         10688 => x"d33978ae",
         10689 => x"38668c2a",
         10690 => x"57810b82",
         10691 => x"b5f42256",
         10692 => x"5a74802e",
         10693 => x"9d387477",
         10694 => x"26983882",
         10695 => x"b5f45679",
         10696 => x"10821770",
         10697 => x"2257575a",
         10698 => x"74802e86",
         10699 => x"38767527",
         10700 => x"ee387952",
         10701 => x"6651fec3",
         10702 => x"ea3f82bb",
         10703 => x"98081084",
         10704 => x"055782bb",
         10705 => x"98089ff5",
         10706 => x"26963881",
         10707 => x"0b82bb98",
         10708 => x"081082bb",
         10709 => x"98080571",
         10710 => x"11722a83",
         10711 => x"0559565e",
         10712 => x"83ff1789",
         10713 => x"2a5d815c",
         10714 => x"a044601c",
         10715 => x"7d116505",
         10716 => x"697012ff",
         10717 => x"05713070",
         10718 => x"72067431",
         10719 => x"5c525957",
         10720 => x"59407d83",
         10721 => x"2e098106",
         10722 => x"8938761c",
         10723 => x"6018415c",
         10724 => x"8439761d",
         10725 => x"5d799029",
         10726 => x"18706231",
         10727 => x"68585155",
         10728 => x"74762687",
         10729 => x"af38757c",
         10730 => x"317d317a",
         10731 => x"53706531",
         10732 => x"5255fec2",
         10733 => x"ee3f82bb",
         10734 => x"9808587d",
         10735 => x"832e0981",
         10736 => x"069b3882",
         10737 => x"bb980883",
         10738 => x"fff52680",
         10739 => x"dd387887",
         10740 => x"83387981",
         10741 => x"2a5978fd",
         10742 => x"be3886f8",
         10743 => x"397d822e",
         10744 => x"09810680",
         10745 => x"c53883ff",
         10746 => x"f50b82bb",
         10747 => x"980827a0",
         10748 => x"38788f38",
         10749 => x"791a5574",
         10750 => x"80c02686",
         10751 => x"387459fd",
         10752 => x"96396281",
         10753 => x"06557480",
         10754 => x"2e8f3883",
         10755 => x"5efd8839",
         10756 => x"82bb9808",
         10757 => x"9ff52692",
         10758 => x"387886b8",
         10759 => x"38791a59",
         10760 => x"81807927",
         10761 => x"fcf13886",
         10762 => x"ab398055",
         10763 => x"7d812e09",
         10764 => x"81068338",
         10765 => x"7d559ff5",
         10766 => x"78278b38",
         10767 => x"74810655",
         10768 => x"8e567486",
         10769 => x"9c388480",
         10770 => x"5380527a",
         10771 => x"51ffa2b9",
         10772 => x"3f8b5382",
         10773 => x"b49c527a",
         10774 => x"51ffa28a",
         10775 => x"3f848052",
         10776 => x"8b1b51ff",
         10777 => x"a1b33f79",
         10778 => x"8d1c347b",
         10779 => x"83ffff06",
         10780 => x"528e1b51",
         10781 => x"ffa1a23f",
         10782 => x"810b901c",
         10783 => x"347d8332",
         10784 => x"70307096",
         10785 => x"2a848006",
         10786 => x"54515591",
         10787 => x"1b51ffa1",
         10788 => x"883f6655",
         10789 => x"7483ffff",
         10790 => x"26903874",
         10791 => x"83ffff06",
         10792 => x"52931b51",
         10793 => x"ffa0f23f",
         10794 => x"8a397452",
         10795 => x"a01b51ff",
         10796 => x"a1853ff8",
         10797 => x"0b951c34",
         10798 => x"bf52981b",
         10799 => x"51ffa0d9",
         10800 => x"3f81ff52",
         10801 => x"9a1b51ff",
         10802 => x"a0cf3f60",
         10803 => x"529c1b51",
         10804 => x"ffa0e43f",
         10805 => x"7d832e09",
         10806 => x"810680cb",
         10807 => x"388288b2",
         10808 => x"0a5280c3",
         10809 => x"1b51ffa0",
         10810 => x"ce3f7c52",
         10811 => x"a41b51ff",
         10812 => x"a0c53f82",
         10813 => x"52ac1b51",
         10814 => x"ffa0bc3f",
         10815 => x"8152b01b",
         10816 => x"51ffa095",
         10817 => x"3f8652b2",
         10818 => x"1b51ffa0",
         10819 => x"8c3fff80",
         10820 => x"0b80c01c",
         10821 => x"34a90b80",
         10822 => x"c21c3493",
         10823 => x"5382b4a8",
         10824 => x"5280c71b",
         10825 => x"51ae3982",
         10826 => x"88b20a52",
         10827 => x"a71b51ff",
         10828 => x"a0853f7c",
         10829 => x"83ffff06",
         10830 => x"52961b51",
         10831 => x"ff9fda3f",
         10832 => x"ff800ba4",
         10833 => x"1c34a90b",
         10834 => x"a61c3493",
         10835 => x"5382b4bc",
         10836 => x"52ab1b51",
         10837 => x"ffa08f3f",
         10838 => x"82d4d552",
         10839 => x"83fe1b70",
         10840 => x"5259ff9f",
         10841 => x"b43f8154",
         10842 => x"60537a52",
         10843 => x"7e51ff9b",
         10844 => x"d73f8156",
         10845 => x"82bb9808",
         10846 => x"83e7387d",
         10847 => x"832e0981",
         10848 => x"0680ee38",
         10849 => x"75546086",
         10850 => x"05537a52",
         10851 => x"7e51ff9b",
         10852 => x"b73f8480",
         10853 => x"5380527a",
         10854 => x"51ff9fed",
         10855 => x"3f848b85",
         10856 => x"a4d2527a",
         10857 => x"51ff9f8f",
         10858 => x"3f868a85",
         10859 => x"e4f25283",
         10860 => x"e41b51ff",
         10861 => x"9f813fff",
         10862 => x"185283e8",
         10863 => x"1b51ff9e",
         10864 => x"f63f8252",
         10865 => x"83ec1b51",
         10866 => x"ff9eec3f",
         10867 => x"82d4d552",
         10868 => x"7851ff9e",
         10869 => x"c43f7554",
         10870 => x"60870553",
         10871 => x"7a527e51",
         10872 => x"ff9ae53f",
         10873 => x"75546016",
         10874 => x"537a527e",
         10875 => x"51ff9ad8",
         10876 => x"3f655380",
         10877 => x"527a51ff",
         10878 => x"9f8f3f7f",
         10879 => x"5680587d",
         10880 => x"832e0981",
         10881 => x"069a38f8",
         10882 => x"527a51ff",
         10883 => x"9ea93fff",
         10884 => x"52841b51",
         10885 => x"ff9ea03f",
         10886 => x"f00a5288",
         10887 => x"1b519139",
         10888 => x"87fffff8",
         10889 => x"557d812e",
         10890 => x"8338f855",
         10891 => x"74527a51",
         10892 => x"ff9e843f",
         10893 => x"7c556157",
         10894 => x"74622683",
         10895 => x"38745776",
         10896 => x"5475537a",
         10897 => x"527e51ff",
         10898 => x"99fe3f82",
         10899 => x"bb980882",
         10900 => x"87388480",
         10901 => x"5382bb98",
         10902 => x"08527a51",
         10903 => x"ff9eaa3f",
         10904 => x"76167578",
         10905 => x"31565674",
         10906 => x"cd388118",
         10907 => x"5877802e",
         10908 => x"ff8d3879",
         10909 => x"557d832e",
         10910 => x"83386355",
         10911 => x"61577462",
         10912 => x"26833874",
         10913 => x"57765475",
         10914 => x"537a527e",
         10915 => x"51ff99b8",
         10916 => x"3f82bb98",
         10917 => x"0881c138",
         10918 => x"76167578",
         10919 => x"31565674",
         10920 => x"db388c56",
         10921 => x"7d832e93",
         10922 => x"38865666",
         10923 => x"83ffff26",
         10924 => x"8a388456",
         10925 => x"7d822e83",
         10926 => x"38815664",
         10927 => x"81065877",
         10928 => x"80fe3884",
         10929 => x"80537752",
         10930 => x"7a51ff9d",
         10931 => x"bc3f82d4",
         10932 => x"d5527851",
         10933 => x"ff9cc23f",
         10934 => x"83be1b55",
         10935 => x"77753481",
         10936 => x"0b811634",
         10937 => x"810b8216",
         10938 => x"34778316",
         10939 => x"34758416",
         10940 => x"34606705",
         10941 => x"5680fdc1",
         10942 => x"527551fe",
         10943 => x"bca53ffe",
         10944 => x"0b851634",
         10945 => x"82bb9808",
         10946 => x"822abf07",
         10947 => x"56758616",
         10948 => x"3482bb98",
         10949 => x"08871634",
         10950 => x"605283c6",
         10951 => x"1b51ff9c",
         10952 => x"963f6652",
         10953 => x"83ca1b51",
         10954 => x"ff9c8c3f",
         10955 => x"81547753",
         10956 => x"7a527e51",
         10957 => x"ff98913f",
         10958 => x"815682bb",
         10959 => x"9808a238",
         10960 => x"80538052",
         10961 => x"7e51ff99",
         10962 => x"e33f8156",
         10963 => x"82bb9808",
         10964 => x"90388939",
         10965 => x"8e568a39",
         10966 => x"81568639",
         10967 => x"82bb9808",
         10968 => x"567582bb",
         10969 => x"980c993d",
         10970 => x"0d04f53d",
         10971 => x"0d7d605b",
         10972 => x"59807960",
         10973 => x"ff055a57",
         10974 => x"57767825",
         10975 => x"b4388d3d",
         10976 => x"f8115555",
         10977 => x"8153fc15",
         10978 => x"527951c9",
         10979 => x"dc3f7a81",
         10980 => x"2e098106",
         10981 => x"9c388c3d",
         10982 => x"3355748d",
         10983 => x"2edb3874",
         10984 => x"76708105",
         10985 => x"58348117",
         10986 => x"57748a2e",
         10987 => x"098106c9",
         10988 => x"38807634",
         10989 => x"78557683",
         10990 => x"38765574",
         10991 => x"82bb980c",
         10992 => x"8d3d0d04",
         10993 => x"f73d0d7b",
         10994 => x"028405b3",
         10995 => x"05335957",
         10996 => x"778a2e09",
         10997 => x"81068738",
         10998 => x"8d527651",
         10999 => x"e73f8417",
         11000 => x"08568076",
         11001 => x"24be3888",
         11002 => x"17087717",
         11003 => x"8c055659",
         11004 => x"77753481",
         11005 => x"1656bb76",
         11006 => x"25a1388b",
         11007 => x"3dfc0554",
         11008 => x"75538c17",
         11009 => x"52760851",
         11010 => x"cbdc3f79",
         11011 => x"76327030",
         11012 => x"7072079f",
         11013 => x"2a703053",
         11014 => x"51565675",
         11015 => x"84180c81",
         11016 => x"1988180c",
         11017 => x"8b3d0d04",
         11018 => x"f93d0d79",
         11019 => x"84110856",
         11020 => x"56807524",
         11021 => x"a738893d",
         11022 => x"fc055474",
         11023 => x"538c1652",
         11024 => x"750851cb",
         11025 => x"a13f82bb",
         11026 => x"98089138",
         11027 => x"84160878",
         11028 => x"2e098106",
         11029 => x"87388816",
         11030 => x"08558339",
         11031 => x"ff557482",
         11032 => x"bb980c89",
         11033 => x"3d0d04fd",
         11034 => x"3d0d7554",
         11035 => x"80cc5380",
         11036 => x"527351ff",
         11037 => x"9a933f76",
         11038 => x"740c853d",
         11039 => x"0d04ea3d",
         11040 => x"0d0280e3",
         11041 => x"05336a53",
         11042 => x"863d7053",
         11043 => x"5454d83f",
         11044 => x"73527251",
         11045 => x"feae3f72",
         11046 => x"51ff8d3f",
         11047 => x"983d0d04",
         11048 => x"00ffffff",
         11049 => x"ff00ffff",
         11050 => x"ffff00ff",
         11051 => x"ffffff00",
         11052 => x"00002ba8",
         11053 => x"00002b2c",
         11054 => x"00002b33",
         11055 => x"00002b3a",
         11056 => x"00002b41",
         11057 => x"00002b48",
         11058 => x"00002b4f",
         11059 => x"00002b56",
         11060 => x"00002b5d",
         11061 => x"00002b64",
         11062 => x"00002b6b",
         11063 => x"00002b72",
         11064 => x"00002b78",
         11065 => x"00002b7e",
         11066 => x"00002b84",
         11067 => x"00002b8a",
         11068 => x"00002b90",
         11069 => x"00002b96",
         11070 => x"00002b9c",
         11071 => x"00002ba2",
         11072 => x"0000436a",
         11073 => x"00004370",
         11074 => x"00004376",
         11075 => x"0000437c",
         11076 => x"00004382",
         11077 => x"00004993",
         11078 => x"00004a89",
         11079 => x"00004b81",
         11080 => x"00004dbb",
         11081 => x"00004a71",
         11082 => x"00004868",
         11083 => x"00004c35",
         11084 => x"00004d91",
         11085 => x"00004c73",
         11086 => x"00004d09",
         11087 => x"00004c8f",
         11088 => x"00004b30",
         11089 => x"00004868",
         11090 => x"00004b81",
         11091 => x"00004ba5",
         11092 => x"00004c35",
         11093 => x"00004868",
         11094 => x"00004868",
         11095 => x"00004c8f",
         11096 => x"00004d09",
         11097 => x"00004d91",
         11098 => x"00004dbb",
         11099 => x"00000e2f",
         11100 => x"00001718",
         11101 => x"00001718",
         11102 => x"00000e5e",
         11103 => x"00001718",
         11104 => x"00001718",
         11105 => x"00001718",
         11106 => x"00001718",
         11107 => x"00001718",
         11108 => x"00001718",
         11109 => x"00001718",
         11110 => x"00000e1b",
         11111 => x"00001718",
         11112 => x"00000e46",
         11113 => x"00000e76",
         11114 => x"00001718",
         11115 => x"00001718",
         11116 => x"00001718",
         11117 => x"00001718",
         11118 => x"00001718",
         11119 => x"00001718",
         11120 => x"00001718",
         11121 => x"00001718",
         11122 => x"00001718",
         11123 => x"00001718",
         11124 => x"00001718",
         11125 => x"00001718",
         11126 => x"00001718",
         11127 => x"00001718",
         11128 => x"00001718",
         11129 => x"00001718",
         11130 => x"00001718",
         11131 => x"00001718",
         11132 => x"00001718",
         11133 => x"00001718",
         11134 => x"00001718",
         11135 => x"00001718",
         11136 => x"00001718",
         11137 => x"00001718",
         11138 => x"00001718",
         11139 => x"00001718",
         11140 => x"00001718",
         11141 => x"00001718",
         11142 => x"00001718",
         11143 => x"00001718",
         11144 => x"00001718",
         11145 => x"00001718",
         11146 => x"00001718",
         11147 => x"00001718",
         11148 => x"00001718",
         11149 => x"00001718",
         11150 => x"00000fa6",
         11151 => x"00001718",
         11152 => x"00001718",
         11153 => x"00001718",
         11154 => x"00001718",
         11155 => x"00001114",
         11156 => x"00001718",
         11157 => x"00001718",
         11158 => x"00001718",
         11159 => x"00001718",
         11160 => x"00001718",
         11161 => x"00001718",
         11162 => x"00001718",
         11163 => x"00001718",
         11164 => x"00001718",
         11165 => x"00001718",
         11166 => x"00000ed6",
         11167 => x"0000103d",
         11168 => x"00000ead",
         11169 => x"00000ead",
         11170 => x"00000ead",
         11171 => x"00001718",
         11172 => x"0000103d",
         11173 => x"00001718",
         11174 => x"00001718",
         11175 => x"00000e96",
         11176 => x"00001718",
         11177 => x"00001718",
         11178 => x"000010ea",
         11179 => x"000010f5",
         11180 => x"00001718",
         11181 => x"00001718",
         11182 => x"00000f0f",
         11183 => x"00001718",
         11184 => x"0000111d",
         11185 => x"00001718",
         11186 => x"00001718",
         11187 => x"00001114",
         11188 => x"64696e69",
         11189 => x"74000000",
         11190 => x"64696f63",
         11191 => x"746c0000",
         11192 => x"66696e69",
         11193 => x"74000000",
         11194 => x"666c6f61",
         11195 => x"64000000",
         11196 => x"66657865",
         11197 => x"63000000",
         11198 => x"6d636c65",
         11199 => x"61720000",
         11200 => x"6d636f70",
         11201 => x"79000000",
         11202 => x"6d646966",
         11203 => x"66000000",
         11204 => x"6d64756d",
         11205 => x"70000000",
         11206 => x"6d656200",
         11207 => x"6d656800",
         11208 => x"6d657700",
         11209 => x"68696400",
         11210 => x"68696500",
         11211 => x"68666400",
         11212 => x"68666500",
         11213 => x"63616c6c",
         11214 => x"00000000",
         11215 => x"6a6d7000",
         11216 => x"72657374",
         11217 => x"61727400",
         11218 => x"72657365",
         11219 => x"74000000",
         11220 => x"696e666f",
         11221 => x"00000000",
         11222 => x"74657374",
         11223 => x"00000000",
         11224 => x"74626173",
         11225 => x"69630000",
         11226 => x"6d626173",
         11227 => x"69630000",
         11228 => x"6b696c6f",
         11229 => x"00000000",
         11230 => x"65640000",
         11231 => x"4469736b",
         11232 => x"20457272",
         11233 => x"6f720a00",
         11234 => x"496e7465",
         11235 => x"726e616c",
         11236 => x"20657272",
         11237 => x"6f722e0a",
         11238 => x"00000000",
         11239 => x"4469736b",
         11240 => x"206e6f74",
         11241 => x"20726561",
         11242 => x"64792e0a",
         11243 => x"00000000",
         11244 => x"4e6f2066",
         11245 => x"696c6520",
         11246 => x"666f756e",
         11247 => x"642e0a00",
         11248 => x"4e6f2070",
         11249 => x"61746820",
         11250 => x"666f756e",
         11251 => x"642e0a00",
         11252 => x"496e7661",
         11253 => x"6c696420",
         11254 => x"66696c65",
         11255 => x"6e616d65",
         11256 => x"2e0a0000",
         11257 => x"41636365",
         11258 => x"73732064",
         11259 => x"656e6965",
         11260 => x"642e0a00",
         11261 => x"46696c65",
         11262 => x"20616c72",
         11263 => x"65616479",
         11264 => x"20657869",
         11265 => x"7374732e",
         11266 => x"0a000000",
         11267 => x"46696c65",
         11268 => x"2068616e",
         11269 => x"646c6520",
         11270 => x"696e7661",
         11271 => x"6c69642e",
         11272 => x"0a000000",
         11273 => x"53442069",
         11274 => x"73207772",
         11275 => x"69746520",
         11276 => x"70726f74",
         11277 => x"65637465",
         11278 => x"642e0a00",
         11279 => x"44726976",
         11280 => x"65206e75",
         11281 => x"6d626572",
         11282 => x"20697320",
         11283 => x"696e7661",
         11284 => x"6c69642e",
         11285 => x"0a000000",
         11286 => x"4469736b",
         11287 => x"206e6f74",
         11288 => x"20656e61",
         11289 => x"626c6564",
         11290 => x"2e0a0000",
         11291 => x"4e6f2063",
         11292 => x"6f6d7061",
         11293 => x"7469626c",
         11294 => x"65206669",
         11295 => x"6c657379",
         11296 => x"7374656d",
         11297 => x"20666f75",
         11298 => x"6e64206f",
         11299 => x"6e206469",
         11300 => x"736b2e0a",
         11301 => x"00000000",
         11302 => x"466f726d",
         11303 => x"61742061",
         11304 => x"626f7274",
         11305 => x"65642e0a",
         11306 => x"00000000",
         11307 => x"54696d65",
         11308 => x"6f75742c",
         11309 => x"206f7065",
         11310 => x"72617469",
         11311 => x"6f6e2063",
         11312 => x"616e6365",
         11313 => x"6c6c6564",
         11314 => x"2e0a0000",
         11315 => x"46696c65",
         11316 => x"20697320",
         11317 => x"6c6f636b",
         11318 => x"65642e0a",
         11319 => x"00000000",
         11320 => x"496e7375",
         11321 => x"66666963",
         11322 => x"69656e74",
         11323 => x"206d656d",
         11324 => x"6f72792e",
         11325 => x"0a000000",
         11326 => x"546f6f20",
         11327 => x"6d616e79",
         11328 => x"206f7065",
         11329 => x"6e206669",
         11330 => x"6c65732e",
         11331 => x"0a000000",
         11332 => x"50617261",
         11333 => x"6d657465",
         11334 => x"72732069",
         11335 => x"6e636f72",
         11336 => x"72656374",
         11337 => x"2e0a0000",
         11338 => x"53756363",
         11339 => x"6573732e",
         11340 => x"0a000000",
         11341 => x"556e6b6e",
         11342 => x"6f776e20",
         11343 => x"6572726f",
         11344 => x"722e0a00",
         11345 => x"0a256c75",
         11346 => x"20627974",
         11347 => x"65732025",
         11348 => x"73206174",
         11349 => x"20256c75",
         11350 => x"20627974",
         11351 => x"65732f73",
         11352 => x"65632e0a",
         11353 => x"00000000",
         11354 => x"72656164",
         11355 => x"00000000",
         11356 => x"25303858",
         11357 => x"00000000",
         11358 => x"3a202000",
         11359 => x"25303458",
         11360 => x"00000000",
         11361 => x"20202020",
         11362 => x"20202020",
         11363 => x"00000000",
         11364 => x"25303258",
         11365 => x"00000000",
         11366 => x"20200000",
         11367 => x"207c0000",
         11368 => x"7c0d0a00",
         11369 => x"5a505554",
         11370 => x"41000000",
         11371 => x"0a2a2a20",
         11372 => x"25732028",
         11373 => x"00000000",
         11374 => x"30322f30",
         11375 => x"352f3230",
         11376 => x"32300000",
         11377 => x"76312e35",
         11378 => x"32000000",
         11379 => x"205a5055",
         11380 => x"2c207265",
         11381 => x"76202530",
         11382 => x"32782920",
         11383 => x"25732025",
         11384 => x"73202a2a",
         11385 => x"0a0a0000",
         11386 => x"5a505554",
         11387 => x"4120496e",
         11388 => x"74657272",
         11389 => x"75707420",
         11390 => x"48616e64",
         11391 => x"6c65720a",
         11392 => x"00000000",
         11393 => x"54696d65",
         11394 => x"7220696e",
         11395 => x"74657272",
         11396 => x"7570740a",
         11397 => x"00000000",
         11398 => x"50533220",
         11399 => x"696e7465",
         11400 => x"72727570",
         11401 => x"740a0000",
         11402 => x"494f4354",
         11403 => x"4c205244",
         11404 => x"20696e74",
         11405 => x"65727275",
         11406 => x"70740a00",
         11407 => x"494f4354",
         11408 => x"4c205752",
         11409 => x"20696e74",
         11410 => x"65727275",
         11411 => x"70740a00",
         11412 => x"55415254",
         11413 => x"30205258",
         11414 => x"20696e74",
         11415 => x"65727275",
         11416 => x"70740a00",
         11417 => x"55415254",
         11418 => x"30205458",
         11419 => x"20696e74",
         11420 => x"65727275",
         11421 => x"70740a00",
         11422 => x"55415254",
         11423 => x"31205258",
         11424 => x"20696e74",
         11425 => x"65727275",
         11426 => x"70740a00",
         11427 => x"55415254",
         11428 => x"31205458",
         11429 => x"20696e74",
         11430 => x"65727275",
         11431 => x"70740a00",
         11432 => x"53657474",
         11433 => x"696e6720",
         11434 => x"75702074",
         11435 => x"696d6572",
         11436 => x"2e2e2e0a",
         11437 => x"00000000",
         11438 => x"456e6162",
         11439 => x"6c696e67",
         11440 => x"2074696d",
         11441 => x"65722e2e",
         11442 => x"2e0a0000",
         11443 => x"6175746f",
         11444 => x"65786563",
         11445 => x"2e626174",
         11446 => x"00000000",
         11447 => x"7a707574",
         11448 => x"612e6873",
         11449 => x"74000000",
         11450 => x"303a0000",
         11451 => x"4661696c",
         11452 => x"65642074",
         11453 => x"6f20696e",
         11454 => x"69746961",
         11455 => x"6c697365",
         11456 => x"20736420",
         11457 => x"63617264",
         11458 => x"20302c20",
         11459 => x"706c6561",
         11460 => x"73652069",
         11461 => x"6e697420",
         11462 => x"6d616e75",
         11463 => x"616c6c79",
         11464 => x"2e000000",
         11465 => x"2a200000",
         11466 => x"42616420",
         11467 => x"6469736b",
         11468 => x"20696421",
         11469 => x"00000000",
         11470 => x"496e6974",
         11471 => x"69616c69",
         11472 => x"7365642e",
         11473 => x"0a000000",
         11474 => x"4661696c",
         11475 => x"65642074",
         11476 => x"6f20696e",
         11477 => x"69746961",
         11478 => x"6c697365",
         11479 => x"2e0a0000",
         11480 => x"72633d25",
         11481 => x"640a0000",
         11482 => x"25753a00",
         11483 => x"436c6561",
         11484 => x"72696e67",
         11485 => x"2e2e2e2e",
         11486 => x"00000000",
         11487 => x"436f7079",
         11488 => x"696e672e",
         11489 => x"2e2e0000",
         11490 => x"436f6d70",
         11491 => x"6172696e",
         11492 => x"672e2e2e",
         11493 => x"00000000",
         11494 => x"2530386c",
         11495 => x"78282530",
         11496 => x"3878292d",
         11497 => x"3e253038",
         11498 => x"6c782825",
         11499 => x"30387829",
         11500 => x"0a000000",
         11501 => x"44756d70",
         11502 => x"204d656d",
         11503 => x"6f72790a",
         11504 => x"00000000",
         11505 => x"0a436f6d",
         11506 => x"706c6574",
         11507 => x"652e0a00",
         11508 => x"25303858",
         11509 => x"20253032",
         11510 => x"582d0000",
         11511 => x"3f3f3f0a",
         11512 => x"00000000",
         11513 => x"25303858",
         11514 => x"20253034",
         11515 => x"582d0000",
         11516 => x"25303858",
         11517 => x"20253038",
         11518 => x"582d0000",
         11519 => x"44697361",
         11520 => x"626c696e",
         11521 => x"6720696e",
         11522 => x"74657272",
         11523 => x"75707473",
         11524 => x"0a000000",
         11525 => x"456e6162",
         11526 => x"6c696e67",
         11527 => x"20696e74",
         11528 => x"65727275",
         11529 => x"7074730a",
         11530 => x"00000000",
         11531 => x"44697361",
         11532 => x"626c6564",
         11533 => x"20756172",
         11534 => x"74206669",
         11535 => x"666f0a00",
         11536 => x"456e6162",
         11537 => x"6c696e67",
         11538 => x"20756172",
         11539 => x"74206669",
         11540 => x"666f0a00",
         11541 => x"45786563",
         11542 => x"7574696e",
         11543 => x"6720636f",
         11544 => x"64652040",
         11545 => x"20253038",
         11546 => x"78202e2e",
         11547 => x"2e0a0000",
         11548 => x"43616c6c",
         11549 => x"696e6720",
         11550 => x"636f6465",
         11551 => x"20402025",
         11552 => x"30387820",
         11553 => x"2e2e2e0a",
         11554 => x"00000000",
         11555 => x"43616c6c",
         11556 => x"20726574",
         11557 => x"75726e65",
         11558 => x"6420636f",
         11559 => x"64652028",
         11560 => x"2564292e",
         11561 => x"0a000000",
         11562 => x"52657374",
         11563 => x"61727469",
         11564 => x"6e672061",
         11565 => x"70706c69",
         11566 => x"63617469",
         11567 => x"6f6e2e2e",
         11568 => x"2e0a0000",
         11569 => x"436f6c64",
         11570 => x"20726562",
         11571 => x"6f6f7469",
         11572 => x"6e672e2e",
         11573 => x"2e0a0000",
         11574 => x"5a505500",
         11575 => x"62696e00",
         11576 => x"25643a5c",
         11577 => x"25735c25",
         11578 => x"732e2573",
         11579 => x"00000000",
         11580 => x"25643a5c",
         11581 => x"25735c25",
         11582 => x"73000000",
         11583 => x"25643a5c",
         11584 => x"25730000",
         11585 => x"42616420",
         11586 => x"636f6d6d",
         11587 => x"616e642e",
         11588 => x"00000000",
         11589 => x"52756e6e",
         11590 => x"696e672e",
         11591 => x"2e2e0a00",
         11592 => x"456e6162",
         11593 => x"6c696e67",
         11594 => x"20696e74",
         11595 => x"65727275",
         11596 => x"7074732e",
         11597 => x"2e2e0a00",
         11598 => x"25642f25",
         11599 => x"642f2564",
         11600 => x"2025643a",
         11601 => x"25643a25",
         11602 => x"642e2564",
         11603 => x"25640a00",
         11604 => x"536f4320",
         11605 => x"436f6e66",
         11606 => x"69677572",
         11607 => x"6174696f",
         11608 => x"6e000000",
         11609 => x"20286672",
         11610 => x"6f6d2053",
         11611 => x"6f432063",
         11612 => x"6f6e6669",
         11613 => x"67290000",
         11614 => x"3a0a4465",
         11615 => x"76696365",
         11616 => x"7320696d",
         11617 => x"706c656d",
         11618 => x"656e7465",
         11619 => x"643a0a00",
         11620 => x"20202020",
         11621 => x"57422053",
         11622 => x"4452414d",
         11623 => x"20202825",
         11624 => x"3038583a",
         11625 => x"25303858",
         11626 => x"292e0a00",
         11627 => x"20202020",
         11628 => x"53445241",
         11629 => x"4d202020",
         11630 => x"20202825",
         11631 => x"3038583a",
         11632 => x"25303858",
         11633 => x"292e0a00",
         11634 => x"20202020",
         11635 => x"494e534e",
         11636 => x"20425241",
         11637 => x"4d202825",
         11638 => x"3038583a",
         11639 => x"25303858",
         11640 => x"292e0a00",
         11641 => x"20202020",
         11642 => x"4252414d",
         11643 => x"20202020",
         11644 => x"20202825",
         11645 => x"3038583a",
         11646 => x"25303858",
         11647 => x"292e0a00",
         11648 => x"20202020",
         11649 => x"52414d20",
         11650 => x"20202020",
         11651 => x"20202825",
         11652 => x"3038583a",
         11653 => x"25303858",
         11654 => x"292e0a00",
         11655 => x"20202020",
         11656 => x"53442043",
         11657 => x"41524420",
         11658 => x"20202844",
         11659 => x"65766963",
         11660 => x"6573203d",
         11661 => x"25303264",
         11662 => x"292e0a00",
         11663 => x"20202020",
         11664 => x"54494d45",
         11665 => x"52312020",
         11666 => x"20202854",
         11667 => x"696d6572",
         11668 => x"7320203d",
         11669 => x"25303264",
         11670 => x"292e0a00",
         11671 => x"20202020",
         11672 => x"494e5452",
         11673 => x"20435452",
         11674 => x"4c202843",
         11675 => x"68616e6e",
         11676 => x"656c733d",
         11677 => x"25303264",
         11678 => x"292e0a00",
         11679 => x"20202020",
         11680 => x"57495348",
         11681 => x"424f4e45",
         11682 => x"20425553",
         11683 => x"0a000000",
         11684 => x"20202020",
         11685 => x"57422049",
         11686 => x"32430a00",
         11687 => x"20202020",
         11688 => x"494f4354",
         11689 => x"4c0a0000",
         11690 => x"20202020",
         11691 => x"5053320a",
         11692 => x"00000000",
         11693 => x"20202020",
         11694 => x"5350490a",
         11695 => x"00000000",
         11696 => x"41646472",
         11697 => x"65737365",
         11698 => x"733a0a00",
         11699 => x"20202020",
         11700 => x"43505520",
         11701 => x"52657365",
         11702 => x"74205665",
         11703 => x"63746f72",
         11704 => x"20416464",
         11705 => x"72657373",
         11706 => x"203d2025",
         11707 => x"3038580a",
         11708 => x"00000000",
         11709 => x"20202020",
         11710 => x"43505520",
         11711 => x"4d656d6f",
         11712 => x"72792053",
         11713 => x"74617274",
         11714 => x"20416464",
         11715 => x"72657373",
         11716 => x"203d2025",
         11717 => x"3038580a",
         11718 => x"00000000",
         11719 => x"20202020",
         11720 => x"53746163",
         11721 => x"6b205374",
         11722 => x"61727420",
         11723 => x"41646472",
         11724 => x"65737320",
         11725 => x"20202020",
         11726 => x"203d2025",
         11727 => x"3038580a",
         11728 => x"00000000",
         11729 => x"4d697363",
         11730 => x"3a0a0000",
         11731 => x"20202020",
         11732 => x"5a505520",
         11733 => x"49642020",
         11734 => x"20202020",
         11735 => x"20202020",
         11736 => x"20202020",
         11737 => x"20202020",
         11738 => x"203d2025",
         11739 => x"3034580a",
         11740 => x"00000000",
         11741 => x"20202020",
         11742 => x"53797374",
         11743 => x"656d2043",
         11744 => x"6c6f636b",
         11745 => x"20467265",
         11746 => x"71202020",
         11747 => x"20202020",
         11748 => x"203d2025",
         11749 => x"642e2530",
         11750 => x"34644d48",
         11751 => x"7a0a0000",
         11752 => x"20202020",
         11753 => x"53445241",
         11754 => x"4d20436c",
         11755 => x"6f636b20",
         11756 => x"46726571",
         11757 => x"20202020",
         11758 => x"20202020",
         11759 => x"203d2025",
         11760 => x"642e2530",
         11761 => x"34644d48",
         11762 => x"7a0a0000",
         11763 => x"20202020",
         11764 => x"57697368",
         11765 => x"626f6e65",
         11766 => x"20534452",
         11767 => x"414d2043",
         11768 => x"6c6f636b",
         11769 => x"20467265",
         11770 => x"713d2025",
         11771 => x"642e2530",
         11772 => x"34644d48",
         11773 => x"7a0a0000",
         11774 => x"536d616c",
         11775 => x"6c000000",
         11776 => x"4d656469",
         11777 => x"756d0000",
         11778 => x"466c6578",
         11779 => x"00000000",
         11780 => x"45564f00",
         11781 => x"45564f6d",
         11782 => x"696e0000",
         11783 => x"556e6b6e",
         11784 => x"6f776e00",
         11785 => x"00009980",
         11786 => x"01000000",
         11787 => x"00000002",
         11788 => x"0000997c",
         11789 => x"01000000",
         11790 => x"00000003",
         11791 => x"00009978",
         11792 => x"01000000",
         11793 => x"00000004",
         11794 => x"00009974",
         11795 => x"01000000",
         11796 => x"00000005",
         11797 => x"00009970",
         11798 => x"01000000",
         11799 => x"00000006",
         11800 => x"0000996c",
         11801 => x"01000000",
         11802 => x"00000007",
         11803 => x"00009968",
         11804 => x"01000000",
         11805 => x"00000001",
         11806 => x"00009964",
         11807 => x"01000000",
         11808 => x"00000008",
         11809 => x"00009960",
         11810 => x"01000000",
         11811 => x"0000000b",
         11812 => x"0000995c",
         11813 => x"01000000",
         11814 => x"00000009",
         11815 => x"00009958",
         11816 => x"01000000",
         11817 => x"0000000a",
         11818 => x"00009954",
         11819 => x"04000000",
         11820 => x"0000000d",
         11821 => x"00009950",
         11822 => x"04000000",
         11823 => x"0000000c",
         11824 => x"0000994c",
         11825 => x"04000000",
         11826 => x"0000000e",
         11827 => x"00009948",
         11828 => x"03000000",
         11829 => x"0000000f",
         11830 => x"00009944",
         11831 => x"04000000",
         11832 => x"0000000f",
         11833 => x"00009940",
         11834 => x"04000000",
         11835 => x"00000010",
         11836 => x"0000993c",
         11837 => x"04000000",
         11838 => x"00000011",
         11839 => x"00009938",
         11840 => x"03000000",
         11841 => x"00000012",
         11842 => x"00009934",
         11843 => x"03000000",
         11844 => x"00000013",
         11845 => x"00009930",
         11846 => x"03000000",
         11847 => x"00000014",
         11848 => x"0000992c",
         11849 => x"03000000",
         11850 => x"00000015",
         11851 => x"1b5b4400",
         11852 => x"1b5b4300",
         11853 => x"1b5b4200",
         11854 => x"1b5b4100",
         11855 => x"1b5b367e",
         11856 => x"1b5b357e",
         11857 => x"1b5b347e",
         11858 => x"1b304600",
         11859 => x"1b5b337e",
         11860 => x"1b5b327e",
         11861 => x"1b5b317e",
         11862 => x"10000000",
         11863 => x"0e000000",
         11864 => x"0d000000",
         11865 => x"0b000000",
         11866 => x"08000000",
         11867 => x"06000000",
         11868 => x"05000000",
         11869 => x"04000000",
         11870 => x"03000000",
         11871 => x"02000000",
         11872 => x"01000000",
         11873 => x"68697374",
         11874 => x"6f727900",
         11875 => x"68697374",
         11876 => x"00000000",
         11877 => x"21000000",
         11878 => x"25303464",
         11879 => x"20202573",
         11880 => x"0a000000",
         11881 => x"4661696c",
         11882 => x"65642074",
         11883 => x"6f207265",
         11884 => x"73657420",
         11885 => x"74686520",
         11886 => x"68697374",
         11887 => x"6f727920",
         11888 => x"66696c65",
         11889 => x"20746f20",
         11890 => x"454f462e",
         11891 => x"0a000000",
         11892 => x"43616e6e",
         11893 => x"6f74206f",
         11894 => x"70656e2f",
         11895 => x"63726561",
         11896 => x"74652068",
         11897 => x"6973746f",
         11898 => x"72792066",
         11899 => x"696c652c",
         11900 => x"20646973",
         11901 => x"61626c69",
         11902 => x"6e672e00",
         11903 => x"53440000",
         11904 => x"222a2b2c",
         11905 => x"3a3b3c3d",
         11906 => x"3e3f5b5d",
         11907 => x"7c7f0000",
         11908 => x"46415400",
         11909 => x"46415433",
         11910 => x"32000000",
         11911 => x"ebfe904d",
         11912 => x"53444f53",
         11913 => x"352e3000",
         11914 => x"4e4f204e",
         11915 => x"414d4520",
         11916 => x"20202046",
         11917 => x"41543332",
         11918 => x"20202000",
         11919 => x"4e4f204e",
         11920 => x"414d4520",
         11921 => x"20202046",
         11922 => x"41542020",
         11923 => x"20202000",
         11924 => x"000099fc",
         11925 => x"00000000",
         11926 => x"00000000",
         11927 => x"00000000",
         11928 => x"809a4541",
         11929 => x"8e418f80",
         11930 => x"45454549",
         11931 => x"49498e8f",
         11932 => x"9092924f",
         11933 => x"994f5555",
         11934 => x"59999a9b",
         11935 => x"9c9d9e9f",
         11936 => x"41494f55",
         11937 => x"a5a5a6a7",
         11938 => x"a8a9aaab",
         11939 => x"acadaeaf",
         11940 => x"b0b1b2b3",
         11941 => x"b4b5b6b7",
         11942 => x"b8b9babb",
         11943 => x"bcbdbebf",
         11944 => x"c0c1c2c3",
         11945 => x"c4c5c6c7",
         11946 => x"c8c9cacb",
         11947 => x"cccdcecf",
         11948 => x"d0d1d2d3",
         11949 => x"d4d5d6d7",
         11950 => x"d8d9dadb",
         11951 => x"dcdddedf",
         11952 => x"e0e1e2e3",
         11953 => x"e4e5e6e7",
         11954 => x"e8e9eaeb",
         11955 => x"ecedeeef",
         11956 => x"f0f1f2f3",
         11957 => x"f4f5f6f7",
         11958 => x"f8f9fafb",
         11959 => x"fcfdfeff",
         11960 => x"2b2e2c3b",
         11961 => x"3d5b5d2f",
         11962 => x"5c222a3a",
         11963 => x"3c3e3f7c",
         11964 => x"7f000000",
         11965 => x"00010004",
         11966 => x"00100040",
         11967 => x"01000200",
         11968 => x"00000000",
         11969 => x"00010002",
         11970 => x"00040008",
         11971 => x"00100020",
         11972 => x"00000000",
         11973 => x"00000000",
         11974 => x"00008ed0",
         11975 => x"01020100",
         11976 => x"00000000",
         11977 => x"00000000",
         11978 => x"00008ed8",
         11979 => x"01040100",
         11980 => x"00000000",
         11981 => x"00000000",
         11982 => x"00008ee0",
         11983 => x"01140300",
         11984 => x"00000000",
         11985 => x"00000000",
         11986 => x"00008ee8",
         11987 => x"012b0300",
         11988 => x"00000000",
         11989 => x"00000000",
         11990 => x"00008ef0",
         11991 => x"01300300",
         11992 => x"00000000",
         11993 => x"00000000",
         11994 => x"00008ef8",
         11995 => x"013c0400",
         11996 => x"00000000",
         11997 => x"00000000",
         11998 => x"00008f00",
         11999 => x"013d0400",
         12000 => x"00000000",
         12001 => x"00000000",
         12002 => x"00008f08",
         12003 => x"013f0400",
         12004 => x"00000000",
         12005 => x"00000000",
         12006 => x"00008f10",
         12007 => x"01400400",
         12008 => x"00000000",
         12009 => x"00000000",
         12010 => x"00008f18",
         12011 => x"01410400",
         12012 => x"00000000",
         12013 => x"00000000",
         12014 => x"00008f1c",
         12015 => x"01420400",
         12016 => x"00000000",
         12017 => x"00000000",
         12018 => x"00008f20",
         12019 => x"01430400",
         12020 => x"00000000",
         12021 => x"00000000",
         12022 => x"00008f24",
         12023 => x"01500500",
         12024 => x"00000000",
         12025 => x"00000000",
         12026 => x"00008f28",
         12027 => x"01510500",
         12028 => x"00000000",
         12029 => x"00000000",
         12030 => x"00008f2c",
         12031 => x"01540500",
         12032 => x"00000000",
         12033 => x"00000000",
         12034 => x"00008f30",
         12035 => x"01550500",
         12036 => x"00000000",
         12037 => x"00000000",
         12038 => x"00008f34",
         12039 => x"01790700",
         12040 => x"00000000",
         12041 => x"00000000",
         12042 => x"00008f3c",
         12043 => x"01780700",
         12044 => x"00000000",
         12045 => x"00000000",
         12046 => x"00008f40",
         12047 => x"01820800",
         12048 => x"00000000",
         12049 => x"00000000",
         12050 => x"00008f48",
         12051 => x"01830800",
         12052 => x"00000000",
         12053 => x"00000000",
         12054 => x"00008f50",
         12055 => x"01850800",
         12056 => x"00000000",
         12057 => x"00000000",
         12058 => x"00008f58",
         12059 => x"01870800",
         12060 => x"00000000",
         12061 => x"00000000",
         12062 => x"00008f60",
         12063 => x"018c0900",
         12064 => x"00000000",
         12065 => x"00000000",
         12066 => x"00008f68",
         12067 => x"018d0900",
         12068 => x"00000000",
         12069 => x"00000000",
         12070 => x"00008f70",
         12071 => x"018e0900",
         12072 => x"00000000",
         12073 => x"00000000",
         12074 => x"00008f78",
         12075 => x"018f0900",
         12076 => x"00000000",
         12077 => x"00000000",
         12078 => x"00000000",
         12079 => x"00000000",
         12080 => x"00007fff",
         12081 => x"00000000",
         12082 => x"00007fff",
         12083 => x"00010000",
         12084 => x"00007fff",
         12085 => x"00010000",
         12086 => x"00810000",
         12087 => x"01000000",
         12088 => x"017fffff",
         12089 => x"00000000",
         12090 => x"00000000",
         12091 => x"00007800",
         12092 => x"00000000",
         12093 => x"05f5e100",
         12094 => x"05f5e100",
         12095 => x"05f5e100",
         12096 => x"00000000",
         12097 => x"01010101",
         12098 => x"01010101",
         12099 => x"01011001",
         12100 => x"01000000",
         12101 => x"00000000",
         12102 => x"00000000",
         12103 => x"00000000",
         12104 => x"00000000",
         12105 => x"00000000",
         12106 => x"00000000",
         12107 => x"00000000",
         12108 => x"00000000",
         12109 => x"00000000",
         12110 => x"00000000",
         12111 => x"00000000",
         12112 => x"00000000",
         12113 => x"00000000",
         12114 => x"00000000",
         12115 => x"00000000",
         12116 => x"00000000",
         12117 => x"00000000",
         12118 => x"00000000",
         12119 => x"00000000",
         12120 => x"00000000",
         12121 => x"00000000",
         12122 => x"00000000",
         12123 => x"00000000",
         12124 => x"00000000",
         12125 => x"00009984",
         12126 => x"01000000",
         12127 => x"0000998c",
         12128 => x"01000000",
         12129 => x"00009994",
         12130 => x"02000000",
         12131 => x"00000000",
         12132 => x"00000000",
         12133 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

