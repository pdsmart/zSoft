-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0ba4",
             1 => x"800b0b0b",
             2 => x"0baabb04",
             3 => x"ffffffff",
             4 => x"ffffffff",
             5 => x"ffffffff",
             6 => x"ffffffff",
             7 => x"ffffffff",
             8 => x"0b0b0ba4",
             9 => x"80040b0b",
            10 => x"0ba48404",
            11 => x"0b0b0ba4",
            12 => x"93040b0b",
            13 => x"0ba4a304",
            14 => x"0b0b0ba4",
            15 => x"b3040b0b",
            16 => x"0ba4c304",
            17 => x"0b0b0ba4",
            18 => x"d3040b0b",
            19 => x"0ba4e304",
            20 => x"0b0b0ba4",
            21 => x"f3040b0b",
            22 => x"0ba58304",
            23 => x"0b0b0ba5",
            24 => x"93040b0b",
            25 => x"0ba5a304",
            26 => x"0b0b0ba5",
            27 => x"b3040b0b",
            28 => x"0ba5c304",
            29 => x"0b0b0ba5",
            30 => x"d3040b0b",
            31 => x"0ba5e204",
            32 => x"0b0b0ba5",
            33 => x"f1040b0b",
            34 => x"0ba68004",
            35 => x"0b0b0ba6",
            36 => x"8f040b0b",
            37 => x"0ba69e04",
            38 => x"0b0b0ba6",
            39 => x"ae040b0b",
            40 => x"0ba6be04",
            41 => x"0b0b0ba6",
            42 => x"ce040b0b",
            43 => x"0ba6de04",
            44 => x"0b0b0ba6",
            45 => x"ee040b0b",
            46 => x"0ba6fe04",
            47 => x"0b0b0ba7",
            48 => x"8e040b0b",
            49 => x"0ba79e04",
            50 => x"0b0b0ba7",
            51 => x"ae040b0b",
            52 => x"0ba7be04",
            53 => x"0b0b0ba7",
            54 => x"ce040b0b",
            55 => x"0ba7de04",
            56 => x"0b0b0ba7",
            57 => x"ee040b0b",
            58 => x"0ba7fe04",
            59 => x"0b0b0ba8",
            60 => x"8e040b0b",
            61 => x"0ba89e04",
            62 => x"0b0b0ba8",
            63 => x"ae040b0b",
            64 => x"0ba8be04",
            65 => x"0b0b0ba8",
            66 => x"ce040b0b",
            67 => x"0ba8de04",
            68 => x"0b0b0ba8",
            69 => x"ee040b0b",
            70 => x"0ba8fe04",
            71 => x"0b0b0ba9",
            72 => x"8e040b0b",
            73 => x"0ba99e04",
            74 => x"0b0b0ba9",
            75 => x"ae040b0b",
            76 => x"0ba9be04",
            77 => x"0b0b0ba9",
            78 => x"ce040b0b",
            79 => x"0ba9de04",
            80 => x"0b0b0ba9",
            81 => x"ee040b0b",
            82 => x"0ba9fe04",
            83 => x"0b0b0baa",
            84 => x"8d040b0b",
            85 => x"0baa9c04",
            86 => x"0b0b0baa",
            87 => x"ab040000",
            88 => x"00000000",
            89 => x"00000000",
            90 => x"00000000",
            91 => x"00000000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"00000000",
            97 => x"00000000",
            98 => x"00000000",
            99 => x"00000000",
           100 => x"00000000",
           101 => x"00000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"00000000",
           105 => x"00000000",
           106 => x"00000000",
           107 => x"00000000",
           108 => x"00000000",
           109 => x"00000000",
           110 => x"00000000",
           111 => x"00000000",
           112 => x"00000000",
           113 => x"00000000",
           114 => x"00000000",
           115 => x"00000000",
           116 => x"00000000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"00000000",
           121 => x"00000000",
           122 => x"00000000",
           123 => x"00000000",
           124 => x"00000000",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"00a48004",
           129 => x"828ce80c",
           130 => x"b8a02d82",
           131 => x"8ce80883",
           132 => x"80900482",
           133 => x"8ce80c80",
           134 => x"c9aa2d82",
           135 => x"8ce80883",
           136 => x"80900482",
           137 => x"8ce80c80",
           138 => x"c9e92d82",
           139 => x"8ce80883",
           140 => x"80900482",
           141 => x"8ce80c80",
           142 => x"ca872d82",
           143 => x"8ce80883",
           144 => x"80900482",
           145 => x"8ce80c80",
           146 => x"d0c52d82",
           147 => x"8ce80883",
           148 => x"80900482",
           149 => x"8ce80c80",
           150 => x"d1c32d82",
           151 => x"8ce80883",
           152 => x"80900482",
           153 => x"8ce80c80",
           154 => x"caaa2d82",
           155 => x"8ce80883",
           156 => x"80900482",
           157 => x"8ce80c80",
           158 => x"d1e02d82",
           159 => x"8ce80883",
           160 => x"80900482",
           161 => x"8ce80c80",
           162 => x"d3d22d82",
           163 => x"8ce80883",
           164 => x"80900482",
           165 => x"8ce80c80",
           166 => x"cfeb2d82",
           167 => x"8ce80883",
           168 => x"80900482",
           169 => x"8ce80c80",
           170 => x"cadc2d82",
           171 => x"8ce80883",
           172 => x"80900482",
           173 => x"8ce80c80",
           174 => x"d0812d82",
           175 => x"8ce80883",
           176 => x"80900482",
           177 => x"8ce80c80",
           178 => x"d0a52d82",
           179 => x"8ce80883",
           180 => x"80900482",
           181 => x"8ce80cba",
           182 => x"ad2d828c",
           183 => x"e8088380",
           184 => x"9004828c",
           185 => x"e80cbafe",
           186 => x"2d828ce8",
           187 => x"08838090",
           188 => x"04828ce8",
           189 => x"0cb39a2d",
           190 => x"828ce808",
           191 => x"83809004",
           192 => x"828ce80c",
           193 => x"b4cf2d82",
           194 => x"8ce80883",
           195 => x"80900482",
           196 => x"8ce80cb6",
           197 => x"822d828c",
           198 => x"e8088380",
           199 => x"9004828c",
           200 => x"e80c8198",
           201 => x"a52d828c",
           202 => x"e8088380",
           203 => x"9004828c",
           204 => x"e80c81a5",
           205 => x"962d828c",
           206 => x"e8088380",
           207 => x"9004828c",
           208 => x"e80c819d",
           209 => x"8a2d828c",
           210 => x"e8088380",
           211 => x"9004828c",
           212 => x"e80c81a0",
           213 => x"872d828c",
           214 => x"e8088380",
           215 => x"9004828c",
           216 => x"e80c81aa",
           217 => x"a52d828c",
           218 => x"e8088380",
           219 => x"9004828c",
           220 => x"e80c81b3",
           221 => x"852d828c",
           222 => x"e8088380",
           223 => x"9004828c",
           224 => x"e80c81a3",
           225 => x"f82d828c",
           226 => x"e8088380",
           227 => x"9004828c",
           228 => x"e80c81ad",
           229 => x"c42d828c",
           230 => x"e8088380",
           231 => x"9004828c",
           232 => x"e80c81ae",
           233 => x"e32d828c",
           234 => x"e8088380",
           235 => x"9004828c",
           236 => x"e80c81af",
           237 => x"822d828c",
           238 => x"e8088380",
           239 => x"9004828c",
           240 => x"e80c81b6",
           241 => x"ec2d828c",
           242 => x"e8088380",
           243 => x"9004828c",
           244 => x"e80c81b4",
           245 => x"d22d828c",
           246 => x"e8088380",
           247 => x"9004828c",
           248 => x"e80c81b9",
           249 => x"c02d828c",
           250 => x"e8088380",
           251 => x"9004828c",
           252 => x"e80c81b0",
           253 => x"862d828c",
           254 => x"e8088380",
           255 => x"9004828c",
           256 => x"e80c81bc",
           257 => x"c02d828c",
           258 => x"e8088380",
           259 => x"9004828c",
           260 => x"e80c81bd",
           261 => x"c12d828c",
           262 => x"e8088380",
           263 => x"9004828c",
           264 => x"e80c81a5",
           265 => x"f62d828c",
           266 => x"e8088380",
           267 => x"9004828c",
           268 => x"e80c81a5",
           269 => x"cf2d828c",
           270 => x"e8088380",
           271 => x"9004828c",
           272 => x"e80c81a6",
           273 => x"fa2d828c",
           274 => x"e8088380",
           275 => x"9004828c",
           276 => x"e80c81b0",
           277 => x"dd2d828c",
           278 => x"e8088380",
           279 => x"9004828c",
           280 => x"e80c81be",
           281 => x"b22d828c",
           282 => x"e8088380",
           283 => x"9004828c",
           284 => x"e80c81c0",
           285 => x"bc2d828c",
           286 => x"e8088380",
           287 => x"9004828c",
           288 => x"e80c81c3",
           289 => x"fe2d828c",
           290 => x"e8088380",
           291 => x"9004828c",
           292 => x"e80c8197",
           293 => x"c42d828c",
           294 => x"e8088380",
           295 => x"9004828c",
           296 => x"e80c81c6",
           297 => x"ea2d828c",
           298 => x"e8088380",
           299 => x"9004828c",
           300 => x"e80c81d5",
           301 => x"9f2d828c",
           302 => x"e8088380",
           303 => x"9004828c",
           304 => x"e80c81d3",
           305 => x"8b2d828c",
           306 => x"e8088380",
           307 => x"9004828c",
           308 => x"e80c80e8",
           309 => x"ff2d828c",
           310 => x"e8088380",
           311 => x"9004828c",
           312 => x"e80c80ea",
           313 => x"e92d828c",
           314 => x"e8088380",
           315 => x"9004828c",
           316 => x"e80c80ec",
           317 => x"cd2d828c",
           318 => x"e8088380",
           319 => x"9004828c",
           320 => x"e80cb3c3",
           321 => x"2d828ce8",
           322 => x"08838090",
           323 => x"04828ce8",
           324 => x"0cb4a52d",
           325 => x"828ce808",
           326 => x"83809004",
           327 => x"828ce80c",
           328 => x"b7922d82",
           329 => x"8ce80883",
           330 => x"80900482",
           331 => x"8ce80c81",
           332 => x"d6ba2d82",
           333 => x"8ce80883",
           334 => x"80900482",
           335 => x"8cdc7082",
           336 => x"a49c278e",
           337 => x"38807170",
           338 => x"8405530c",
           339 => x"0b0b0baa",
           340 => x"be04a480",
           341 => x"5181efa0",
           342 => x"043c0482",
           343 => x"8ce80802",
           344 => x"828ce80c",
           345 => x"fd3d0d80",
           346 => x"53828ce8",
           347 => x"088c0508",
           348 => x"52828ce8",
           349 => x"08880508",
           350 => x"5180c53f",
           351 => x"828cdc08",
           352 => x"70828cdc",
           353 => x"0c54853d",
           354 => x"0d828ce8",
           355 => x"0c04828c",
           356 => x"e8080282",
           357 => x"8ce80cfd",
           358 => x"3d0d8153",
           359 => x"828ce808",
           360 => x"8c050852",
           361 => x"828ce808",
           362 => x"88050851",
           363 => x"933f828c",
           364 => x"dc087082",
           365 => x"8cdc0c54",
           366 => x"853d0d82",
           367 => x"8ce80c04",
           368 => x"828ce808",
           369 => x"02828ce8",
           370 => x"0cfd3d0d",
           371 => x"810b828c",
           372 => x"e808fc05",
           373 => x"0c800b82",
           374 => x"8ce808f8",
           375 => x"050c828c",
           376 => x"e8088c05",
           377 => x"08828ce8",
           378 => x"08880508",
           379 => x"27b93882",
           380 => x"8ce808fc",
           381 => x"0508802e",
           382 => x"ae38800b",
           383 => x"828ce808",
           384 => x"8c050824",
           385 => x"a238828c",
           386 => x"e8088c05",
           387 => x"0810828c",
           388 => x"e8088c05",
           389 => x"0c828ce8",
           390 => x"08fc0508",
           391 => x"10828ce8",
           392 => x"08fc050c",
           393 => x"ffb83982",
           394 => x"8ce808fc",
           395 => x"0508802e",
           396 => x"80e13882",
           397 => x"8ce8088c",
           398 => x"0508828c",
           399 => x"e8088805",
           400 => x"0826ad38",
           401 => x"828ce808",
           402 => x"88050882",
           403 => x"8ce8088c",
           404 => x"05083182",
           405 => x"8ce80888",
           406 => x"050c828c",
           407 => x"e808f805",
           408 => x"08828ce8",
           409 => x"08fc0508",
           410 => x"07828ce8",
           411 => x"08f8050c",
           412 => x"828ce808",
           413 => x"fc050881",
           414 => x"2a828ce8",
           415 => x"08fc050c",
           416 => x"828ce808",
           417 => x"8c050881",
           418 => x"2a828ce8",
           419 => x"088c050c",
           420 => x"ff953982",
           421 => x"8ce80890",
           422 => x"0508802e",
           423 => x"9338828c",
           424 => x"e8088805",
           425 => x"0870828c",
           426 => x"e808f405",
           427 => x"0c519139",
           428 => x"828ce808",
           429 => x"f8050870",
           430 => x"828ce808",
           431 => x"f4050c51",
           432 => x"828ce808",
           433 => x"f4050882",
           434 => x"8cdc0c85",
           435 => x"3d0d828c",
           436 => x"e80c04fc",
           437 => x"3d0d7670",
           438 => x"797b5555",
           439 => x"55558f72",
           440 => x"278c3872",
           441 => x"75078306",
           442 => x"5170802e",
           443 => x"a938ff12",
           444 => x"5271ff2e",
           445 => x"98387270",
           446 => x"81055433",
           447 => x"74708105",
           448 => x"5634ff12",
           449 => x"5271ff2e",
           450 => x"098106ea",
           451 => x"3874828c",
           452 => x"dc0c863d",
           453 => x"0d047451",
           454 => x"72708405",
           455 => x"54087170",
           456 => x"8405530c",
           457 => x"72708405",
           458 => x"54087170",
           459 => x"8405530c",
           460 => x"72708405",
           461 => x"54087170",
           462 => x"8405530c",
           463 => x"72708405",
           464 => x"54087170",
           465 => x"8405530c",
           466 => x"f0125271",
           467 => x"8f26c938",
           468 => x"83722795",
           469 => x"38727084",
           470 => x"05540871",
           471 => x"70840553",
           472 => x"0cfc1252",
           473 => x"718326ed",
           474 => x"387054ff",
           475 => x"8139fc3d",
           476 => x"0d767971",
           477 => x"028c059f",
           478 => x"05335755",
           479 => x"53558372",
           480 => x"278a3874",
           481 => x"83065170",
           482 => x"802ea438",
           483 => x"ff125271",
           484 => x"ff2e9338",
           485 => x"73737081",
           486 => x"055534ff",
           487 => x"125271ff",
           488 => x"2e098106",
           489 => x"ef387482",
           490 => x"8cdc0c86",
           491 => x"3d0d0474",
           492 => x"74882b75",
           493 => x"07707190",
           494 => x"2b075154",
           495 => x"518f7227",
           496 => x"a5387271",
           497 => x"70840553",
           498 => x"0c727170",
           499 => x"8405530c",
           500 => x"72717084",
           501 => x"05530c72",
           502 => x"71708405",
           503 => x"530cf012",
           504 => x"52718f26",
           505 => x"dd388372",
           506 => x"27903872",
           507 => x"71708405",
           508 => x"530cfc12",
           509 => x"52718326",
           510 => x"f2387053",
           511 => x"ff8e39fc",
           512 => x"3d0d7670",
           513 => x"79707307",
           514 => x"83065454",
           515 => x"54557080",
           516 => x"c3387170",
           517 => x"08700970",
           518 => x"f7fbfdff",
           519 => x"130670f8",
           520 => x"84828180",
           521 => x"06515153",
           522 => x"535470a6",
           523 => x"38841472",
           524 => x"74708405",
           525 => x"560c7008",
           526 => x"700970f7",
           527 => x"fbfdff13",
           528 => x"0670f884",
           529 => x"82818006",
           530 => x"51515353",
           531 => x"5470802e",
           532 => x"dc387352",
           533 => x"71708105",
           534 => x"53335170",
           535 => x"73708105",
           536 => x"553470f0",
           537 => x"3874828c",
           538 => x"dc0c863d",
           539 => x"0d04fd3d",
           540 => x"0d757071",
           541 => x"83065355",
           542 => x"5270b838",
           543 => x"71700870",
           544 => x"09f7fbfd",
           545 => x"ff120670",
           546 => x"f8848281",
           547 => x"80065151",
           548 => x"5253709d",
           549 => x"38841370",
           550 => x"087009f7",
           551 => x"fbfdff12",
           552 => x"0670f884",
           553 => x"82818006",
           554 => x"51515253",
           555 => x"70802ee5",
           556 => x"38725271",
           557 => x"33517080",
           558 => x"2e8a3881",
           559 => x"12703352",
           560 => x"5270f838",
           561 => x"71743182",
           562 => x"8cdc0c85",
           563 => x"3d0d04fa",
           564 => x"3d0d787a",
           565 => x"7c705455",
           566 => x"55527280",
           567 => x"2e80d938",
           568 => x"71740783",
           569 => x"06517080",
           570 => x"2e80d638",
           571 => x"ff135372",
           572 => x"ff2eb138",
           573 => x"71337433",
           574 => x"56517471",
           575 => x"2e098106",
           576 => x"a9387280",
           577 => x"2e818938",
           578 => x"7081ff06",
           579 => x"5170802e",
           580 => x"80fe3881",
           581 => x"128115ff",
           582 => x"15555552",
           583 => x"72ff2e09",
           584 => x"8106d138",
           585 => x"71337433",
           586 => x"56517081",
           587 => x"ff067581",
           588 => x"ff067171",
           589 => x"31515252",
           590 => x"70828cdc",
           591 => x"0c883d0d",
           592 => x"04717457",
           593 => x"55837327",
           594 => x"88387108",
           595 => x"74082e88",
           596 => x"38747655",
           597 => x"52ff9539",
           598 => x"fc135372",
           599 => x"802eb138",
           600 => x"74087009",
           601 => x"f7fbfdff",
           602 => x"120670f8",
           603 => x"84828180",
           604 => x"06515151",
           605 => x"709a3884",
           606 => x"15841757",
           607 => x"55837327",
           608 => x"d0387408",
           609 => x"76082ed0",
           610 => x"38747655",
           611 => x"52fedd39",
           612 => x"800b828c",
           613 => x"dc0c883d",
           614 => x"0d04fe3d",
           615 => x"0d805283",
           616 => x"5371882b",
           617 => x"5287863f",
           618 => x"828cdc08",
           619 => x"81ff0672",
           620 => x"07ff1454",
           621 => x"52728025",
           622 => x"e8387182",
           623 => x"8cdc0c84",
           624 => x"3d0d04fb",
           625 => x"3d0d7770",
           626 => x"08705353",
           627 => x"5671802e",
           628 => x"80ca3871",
           629 => x"335170a0",
           630 => x"2e098106",
           631 => x"86388112",
           632 => x"52f13971",
           633 => x"53843981",
           634 => x"13538073",
           635 => x"337081ff",
           636 => x"06535555",
           637 => x"70a02e83",
           638 => x"38815570",
           639 => x"802e8438",
           640 => x"74e53873",
           641 => x"81ff0651",
           642 => x"70a02e09",
           643 => x"81068838",
           644 => x"80737081",
           645 => x"05553472",
           646 => x"760c7151",
           647 => x"70828cdc",
           648 => x"0c873d0d",
           649 => x"04fc3d0d",
           650 => x"76537208",
           651 => x"802e9138",
           652 => x"863dfc05",
           653 => x"5272519f",
           654 => x"993f828c",
           655 => x"dc088538",
           656 => x"80538339",
           657 => x"74537282",
           658 => x"8cdc0c86",
           659 => x"3d0d04fc",
           660 => x"3d0d7682",
           661 => x"1133ff05",
           662 => x"52538152",
           663 => x"708b2681",
           664 => x"98388313",
           665 => x"33ff0551",
           666 => x"8252709e",
           667 => x"26818a38",
           668 => x"84133351",
           669 => x"83527097",
           670 => x"2680fe38",
           671 => x"85133351",
           672 => x"845270bb",
           673 => x"2680f238",
           674 => x"86133351",
           675 => x"855270bb",
           676 => x"2680e638",
           677 => x"88132255",
           678 => x"86527487",
           679 => x"e72680d9",
           680 => x"388a1322",
           681 => x"54875273",
           682 => x"87e72680",
           683 => x"cc38810b",
           684 => x"87c0989c",
           685 => x"0c722287",
           686 => x"c098bc0c",
           687 => x"82133387",
           688 => x"c098b80c",
           689 => x"83133387",
           690 => x"c098b40c",
           691 => x"84133387",
           692 => x"c098b00c",
           693 => x"85133387",
           694 => x"c098ac0c",
           695 => x"86133387",
           696 => x"c098a80c",
           697 => x"7487c098",
           698 => x"a40c7387",
           699 => x"c098a00c",
           700 => x"800b87c0",
           701 => x"989c0c80",
           702 => x"5271828c",
           703 => x"dc0c863d",
           704 => x"0d04f33d",
           705 => x"0d7f5b87",
           706 => x"c0989c5d",
           707 => x"817d0c87",
           708 => x"c098bc08",
           709 => x"5e7d7b23",
           710 => x"87c098b8",
           711 => x"085a7982",
           712 => x"1c3487c0",
           713 => x"98b4085a",
           714 => x"79831c34",
           715 => x"87c098b0",
           716 => x"085a7984",
           717 => x"1c3487c0",
           718 => x"98ac085a",
           719 => x"79851c34",
           720 => x"87c098a8",
           721 => x"085a7986",
           722 => x"1c3487c0",
           723 => x"98a4085c",
           724 => x"7b881c23",
           725 => x"87c098a0",
           726 => x"085a798a",
           727 => x"1c23807d",
           728 => x"0c7983ff",
           729 => x"ff06597b",
           730 => x"83ffff06",
           731 => x"58861b33",
           732 => x"57851b33",
           733 => x"56841b33",
           734 => x"55831b33",
           735 => x"54821b33",
           736 => x"537d83ff",
           737 => x"ff065281",
           738 => x"f1e45198",
           739 => x"de3f8f3d",
           740 => x"0d04ff3d",
           741 => x"0d028f05",
           742 => x"33703070",
           743 => x"9f2a5152",
           744 => x"52700b0b",
           745 => x"8287d434",
           746 => x"833d0d04",
           747 => x"fb3d0d77",
           748 => x"0b0b8287",
           749 => x"d4337081",
           750 => x"ff065755",
           751 => x"5687c094",
           752 => x"84517480",
           753 => x"2e863887",
           754 => x"c0949451",
           755 => x"70087096",
           756 => x"2a708106",
           757 => x"53545270",
           758 => x"802e8c38",
           759 => x"71912a70",
           760 => x"81065151",
           761 => x"70d73872",
           762 => x"81327081",
           763 => x"06515170",
           764 => x"802e8d38",
           765 => x"71932a70",
           766 => x"81065151",
           767 => x"70ffbe38",
           768 => x"7381ff06",
           769 => x"5187c094",
           770 => x"80527080",
           771 => x"2e863887",
           772 => x"c0949052",
           773 => x"75720c75",
           774 => x"828cdc0c",
           775 => x"873d0d04",
           776 => x"fb3d0d02",
           777 => x"9f05330b",
           778 => x"0b8287d4",
           779 => x"337081ff",
           780 => x"06575556",
           781 => x"87c09484",
           782 => x"5174802e",
           783 => x"863887c0",
           784 => x"94945170",
           785 => x"0870962a",
           786 => x"70810653",
           787 => x"54527080",
           788 => x"2e8c3871",
           789 => x"912a7081",
           790 => x"06515170",
           791 => x"d7387281",
           792 => x"32708106",
           793 => x"51517080",
           794 => x"2e8d3871",
           795 => x"932a7081",
           796 => x"06515170",
           797 => x"ffbe3873",
           798 => x"81ff0651",
           799 => x"87c09480",
           800 => x"5270802e",
           801 => x"863887c0",
           802 => x"94905275",
           803 => x"720c873d",
           804 => x"0d04f93d",
           805 => x"0d795480",
           806 => x"74337081",
           807 => x"ff065353",
           808 => x"5770772e",
           809 => x"80fe3871",
           810 => x"81ff0681",
           811 => x"150b0b82",
           812 => x"87d43370",
           813 => x"81ff0659",
           814 => x"57555887",
           815 => x"c0948451",
           816 => x"75802e86",
           817 => x"3887c094",
           818 => x"94517008",
           819 => x"70962a70",
           820 => x"81065354",
           821 => x"5270802e",
           822 => x"8c387191",
           823 => x"2a708106",
           824 => x"515170d7",
           825 => x"38728132",
           826 => x"70810651",
           827 => x"5170802e",
           828 => x"8d387193",
           829 => x"2a708106",
           830 => x"515170ff",
           831 => x"be387481",
           832 => x"ff065187",
           833 => x"c0948052",
           834 => x"70802e86",
           835 => x"3887c094",
           836 => x"90527772",
           837 => x"0c811774",
           838 => x"337081ff",
           839 => x"06535357",
           840 => x"70ff8438",
           841 => x"76828cdc",
           842 => x"0c893d0d",
           843 => x"04fe3d0d",
           844 => x"0b0b8287",
           845 => x"d4337081",
           846 => x"ff065452",
           847 => x"87c09484",
           848 => x"5172802e",
           849 => x"863887c0",
           850 => x"94945170",
           851 => x"0870822a",
           852 => x"70810651",
           853 => x"51517080",
           854 => x"2ee23871",
           855 => x"81ff0651",
           856 => x"87c09480",
           857 => x"5270802e",
           858 => x"863887c0",
           859 => x"94905271",
           860 => x"087081ff",
           861 => x"06828cdc",
           862 => x"0c51843d",
           863 => x"0d04fe3d",
           864 => x"0d0b0b82",
           865 => x"87d43370",
           866 => x"81ff0652",
           867 => x"5387c094",
           868 => x"84527080",
           869 => x"2e863887",
           870 => x"c0949452",
           871 => x"71087082",
           872 => x"2a708106",
           873 => x"515151ff",
           874 => x"5270802e",
           875 => x"a0387281",
           876 => x"ff065187",
           877 => x"c0948052",
           878 => x"70802e86",
           879 => x"3887c094",
           880 => x"90527108",
           881 => x"70982b70",
           882 => x"982c5153",
           883 => x"5171828c",
           884 => x"dc0c843d",
           885 => x"0d04ff3d",
           886 => x"0d87c09e",
           887 => x"8008709c",
           888 => x"2a8a0651",
           889 => x"5170802e",
           890 => x"84b43887",
           891 => x"c09ea408",
           892 => x"8287d80c",
           893 => x"87c09ea8",
           894 => x"088287dc",
           895 => x"0c87c09e",
           896 => x"94088287",
           897 => x"e00c87c0",
           898 => x"9e980882",
           899 => x"87e40c87",
           900 => x"c09e9c08",
           901 => x"8287e80c",
           902 => x"87c09ea0",
           903 => x"088287ec",
           904 => x"0c87c09e",
           905 => x"ac088287",
           906 => x"f00c87c0",
           907 => x"9eb00882",
           908 => x"87f40c87",
           909 => x"c09eb408",
           910 => x"8287f80c",
           911 => x"87c09eb8",
           912 => x"088287fc",
           913 => x"0c87c09e",
           914 => x"bc088288",
           915 => x"800c87c0",
           916 => x"9ec00882",
           917 => x"88840c87",
           918 => x"c09ec408",
           919 => x"8288880c",
           920 => x"87c09e80",
           921 => x"08517082",
           922 => x"888c2387",
           923 => x"c09e8408",
           924 => x"8288900c",
           925 => x"87c09e88",
           926 => x"08828894",
           927 => x"0c87c09e",
           928 => x"8c088288",
           929 => x"980c810b",
           930 => x"82889c34",
           931 => x"800b87c0",
           932 => x"9e900870",
           933 => x"84800a06",
           934 => x"51525270",
           935 => x"802e8338",
           936 => x"81527182",
           937 => x"889d3480",
           938 => x"0b87c09e",
           939 => x"90087088",
           940 => x"800a0651",
           941 => x"52527080",
           942 => x"2e833881",
           943 => x"52718288",
           944 => x"9e34800b",
           945 => x"87c09e90",
           946 => x"08709080",
           947 => x"0a065152",
           948 => x"5270802e",
           949 => x"83388152",
           950 => x"7182889f",
           951 => x"34800b87",
           952 => x"c09e9008",
           953 => x"70888080",
           954 => x"06515252",
           955 => x"70802e83",
           956 => x"38815271",
           957 => x"8288a034",
           958 => x"800b87c0",
           959 => x"9e900870",
           960 => x"a0808006",
           961 => x"51525270",
           962 => x"802e8338",
           963 => x"81527182",
           964 => x"88a13480",
           965 => x"0b87c09e",
           966 => x"90087090",
           967 => x"80800651",
           968 => x"52527080",
           969 => x"2e833881",
           970 => x"52718288",
           971 => x"a234800b",
           972 => x"87c09e90",
           973 => x"08708480",
           974 => x"80065152",
           975 => x"5270802e",
           976 => x"83388152",
           977 => x"718288a3",
           978 => x"34800b87",
           979 => x"c09e9008",
           980 => x"70828080",
           981 => x"06515252",
           982 => x"70802e83",
           983 => x"38815271",
           984 => x"8288a434",
           985 => x"800b87c0",
           986 => x"9e900870",
           987 => x"81808006",
           988 => x"51525270",
           989 => x"802e8338",
           990 => x"81527182",
           991 => x"88a53480",
           992 => x"0b87c09e",
           993 => x"90087080",
           994 => x"c0800651",
           995 => x"52527080",
           996 => x"2e833881",
           997 => x"52718288",
           998 => x"a634800b",
           999 => x"87c09e90",
          1000 => x"0870a080",
          1001 => x"06515252",
          1002 => x"70802e83",
          1003 => x"38815271",
          1004 => x"8288a734",
          1005 => x"87c09e90",
          1006 => x"08709880",
          1007 => x"06708a2a",
          1008 => x"51515170",
          1009 => x"8288a834",
          1010 => x"800b87c0",
          1011 => x"9e900870",
          1012 => x"84800651",
          1013 => x"52527080",
          1014 => x"2e833881",
          1015 => x"52718288",
          1016 => x"a93487c0",
          1017 => x"9e900870",
          1018 => x"83f00670",
          1019 => x"842a5151",
          1020 => x"51708288",
          1021 => x"aa34800b",
          1022 => x"87c09e90",
          1023 => x"08708806",
          1024 => x"51525270",
          1025 => x"802e8338",
          1026 => x"81527182",
          1027 => x"88ab3487",
          1028 => x"c09e9008",
          1029 => x"70870651",
          1030 => x"51708288",
          1031 => x"ac34833d",
          1032 => x"0d04fb3d",
          1033 => x"0d81f1fc",
          1034 => x"5189dc3f",
          1035 => x"82889c33",
          1036 => x"5473802e",
          1037 => x"883881f2",
          1038 => x"905189cb",
          1039 => x"3f81f2a4",
          1040 => x"5189c43f",
          1041 => x"82889e33",
          1042 => x"5473802e",
          1043 => x"93388287",
          1044 => x"f8088287",
          1045 => x"fc081154",
          1046 => x"5281f2bc",
          1047 => x"518f8c3f",
          1048 => x"8288a333",
          1049 => x"5473802e",
          1050 => x"93388287",
          1051 => x"f0088287",
          1052 => x"f4081154",
          1053 => x"5281f2d8",
          1054 => x"518ef03f",
          1055 => x"8288a033",
          1056 => x"5473802e",
          1057 => x"93388287",
          1058 => x"d8088287",
          1059 => x"dc081154",
          1060 => x"5281f2f4",
          1061 => x"518ed43f",
          1062 => x"8288a133",
          1063 => x"5473802e",
          1064 => x"93388287",
          1065 => x"e0088287",
          1066 => x"e4081154",
          1067 => x"5281f390",
          1068 => x"518eb83f",
          1069 => x"8288a233",
          1070 => x"5473802e",
          1071 => x"93388287",
          1072 => x"e8088287",
          1073 => x"ec081154",
          1074 => x"5281f3ac",
          1075 => x"518e9c3f",
          1076 => x"8288a733",
          1077 => x"5473802e",
          1078 => x"8d388288",
          1079 => x"a8335281",
          1080 => x"f3c8518e",
          1081 => x"863f8288",
          1082 => x"ab335473",
          1083 => x"802e8d38",
          1084 => x"8288ac33",
          1085 => x"5281f3e8",
          1086 => x"518df03f",
          1087 => x"8288a933",
          1088 => x"5473802e",
          1089 => x"8d388288",
          1090 => x"aa335281",
          1091 => x"f488518d",
          1092 => x"da3f8288",
          1093 => x"9d335473",
          1094 => x"802e8838",
          1095 => x"81f4a851",
          1096 => x"87e53f82",
          1097 => x"889f3354",
          1098 => x"73802e88",
          1099 => x"3881f4bc",
          1100 => x"5187d43f",
          1101 => x"8288a433",
          1102 => x"5473802e",
          1103 => x"883881f4",
          1104 => x"c85187c3",
          1105 => x"3f8288a5",
          1106 => x"33547380",
          1107 => x"2e883881",
          1108 => x"f4d45187",
          1109 => x"b23f8288",
          1110 => x"a6335473",
          1111 => x"802e8838",
          1112 => x"81f4e051",
          1113 => x"87a13f81",
          1114 => x"f4ec5187",
          1115 => x"9a3f8288",
          1116 => x"80085281",
          1117 => x"f4f8518c",
          1118 => x"f23f8288",
          1119 => x"84085281",
          1120 => x"f5a0518c",
          1121 => x"e63f8288",
          1122 => x"88085281",
          1123 => x"f5c8518c",
          1124 => x"da3f81f5",
          1125 => x"f05186ef",
          1126 => x"3f82888c",
          1127 => x"225281f5",
          1128 => x"f8518cc7",
          1129 => x"3f828890",
          1130 => x"0856bd84",
          1131 => x"c0527551",
          1132 => x"e7a93f82",
          1133 => x"8cdc08bd",
          1134 => x"84c02976",
          1135 => x"71315454",
          1136 => x"828cdc08",
          1137 => x"5281f6a0",
          1138 => x"518ca03f",
          1139 => x"8288a333",
          1140 => x"5473802e",
          1141 => x"a8388288",
          1142 => x"940856bd",
          1143 => x"84c05275",
          1144 => x"51e6f83f",
          1145 => x"828cdc08",
          1146 => x"bd84c029",
          1147 => x"76713154",
          1148 => x"54828cdc",
          1149 => x"085281f6",
          1150 => x"cc518bef",
          1151 => x"3f82889e",
          1152 => x"33547380",
          1153 => x"2ea83882",
          1154 => x"88980856",
          1155 => x"bd84c052",
          1156 => x"7551e6c7",
          1157 => x"3f828cdc",
          1158 => x"08bd84c0",
          1159 => x"29767131",
          1160 => x"5454828c",
          1161 => x"dc085281",
          1162 => x"f6f8518b",
          1163 => x"be3f8285",
          1164 => x"a45185d3",
          1165 => x"3f873d0d",
          1166 => x"04fe3d0d",
          1167 => x"02920533",
          1168 => x"ff055271",
          1169 => x"8426ac38",
          1170 => x"7184290b",
          1171 => x"0b81f0d0",
          1172 => x"05527108",
          1173 => x"0481f7a4",
          1174 => x"519d3981",
          1175 => x"f7ac5197",
          1176 => x"3981f7b4",
          1177 => x"51913981",
          1178 => x"f7bc518b",
          1179 => x"3981f7c0",
          1180 => x"51853981",
          1181 => x"f7c85185",
          1182 => x"8e3f843d",
          1183 => x"0d047188",
          1184 => x"800c0480",
          1185 => x"0b87c096",
          1186 => x"840c0482",
          1187 => x"88b00887",
          1188 => x"c096840c",
          1189 => x"04fe3d0d",
          1190 => x"828cec08",
          1191 => x"893882a4",
          1192 => x"9c0b828c",
          1193 => x"ec0c828c",
          1194 => x"ec087511",
          1195 => x"5252ff53",
          1196 => x"7083b7f8",
          1197 => x"26883870",
          1198 => x"828cec0c",
          1199 => x"71537282",
          1200 => x"8cdc0c84",
          1201 => x"3d0d04f9",
          1202 => x"3d0d797b",
          1203 => x"841208a0",
          1204 => x"12901408",
          1205 => x"94150890",
          1206 => x"165e5a58",
          1207 => x"54595753",
          1208 => x"707726ba",
          1209 => x"38751388",
          1210 => x"14085351",
          1211 => x"81710c76",
          1212 => x"76318412",
          1213 => x"0c80730c",
          1214 => x"7584140c",
          1215 => x"728c120c",
          1216 => x"7188120c",
          1217 => x"708c130c",
          1218 => x"7088140c",
          1219 => x"7390120c",
          1220 => x"7494120c",
          1221 => x"7094150c",
          1222 => x"7090160c",
          1223 => x"8c398073",
          1224 => x"0c739016",
          1225 => x"0c749415",
          1226 => x"0c77828c",
          1227 => x"dc0c893d",
          1228 => x"0d04fc3d",
          1229 => x"0d768c11",
          1230 => x"08881208",
          1231 => x"56535371",
          1232 => x"08812e09",
          1233 => x"8106a338",
          1234 => x"84120870",
          1235 => x"13525570",
          1236 => x"732e0981",
          1237 => x"06943884",
          1238 => x"13081584",
          1239 => x"130c7388",
          1240 => x"130c718c",
          1241 => x"150c7153",
          1242 => x"9f398173",
          1243 => x"0c8288c4",
          1244 => x"0890140c",
          1245 => x"8288b40b",
          1246 => x"94140c72",
          1247 => x"8288c40c",
          1248 => x"90130873",
          1249 => x"94120c51",
          1250 => x"7308812e",
          1251 => x"098106b3",
          1252 => x"38841308",
          1253 => x"70145252",
          1254 => x"70742e09",
          1255 => x"8106a438",
          1256 => x"84140812",
          1257 => x"84140c94",
          1258 => x"14089015",
          1259 => x"08709013",
          1260 => x"0c529412",
          1261 => x"0c8c1408",
          1262 => x"88150870",
          1263 => x"88130c52",
          1264 => x"8c120c72",
          1265 => x"828cdc0c",
          1266 => x"863d0d04",
          1267 => x"f93d0d79",
          1268 => x"70555776",
          1269 => x"802e81b5",
          1270 => x"389f17f0",
          1271 => x"068288c4",
          1272 => x"08575775",
          1273 => x"08822e8f",
          1274 => x"38841608",
          1275 => x"772780c7",
          1276 => x"38901608",
          1277 => x"56ed3983",
          1278 => x"ffff17fc",
          1279 => x"80800670",
          1280 => x"5258fd91",
          1281 => x"3f828cdc",
          1282 => x"08828cdc",
          1283 => x"08307082",
          1284 => x"8cdc0807",
          1285 => x"8025828c",
          1286 => x"dc080970",
          1287 => x"30707207",
          1288 => x"80257307",
          1289 => x"53585851",
          1290 => x"54568054",
          1291 => x"72742e09",
          1292 => x"810680d9",
          1293 => x"38883976",
          1294 => x"52755180",
          1295 => x"c839810b",
          1296 => x"828cdc08",
          1297 => x"0c77828c",
          1298 => x"dc088405",
          1299 => x"0c8288c0",
          1300 => x"08537208",
          1301 => x"822e8c38",
          1302 => x"75732687",
          1303 => x"388c1308",
          1304 => x"53f03988",
          1305 => x"13088817",
          1306 => x"0c728c17",
          1307 => x"0c758814",
          1308 => x"0c881608",
          1309 => x"768c120c",
          1310 => x"537551fd",
          1311 => x"b53f7652",
          1312 => x"828cdc08",
          1313 => x"51fcc03f",
          1314 => x"828cdc08",
          1315 => x"5473828c",
          1316 => x"dc0c893d",
          1317 => x"0d04ff3d",
          1318 => x"0d735271",
          1319 => x"802e8738",
          1320 => x"f01251fd",
          1321 => x"8d3f833d",
          1322 => x"0d04fe3d",
          1323 => x"0d029305",
          1324 => x"3353728a",
          1325 => x"2e098106",
          1326 => x"85388d51",
          1327 => x"ed3f828c",
          1328 => x"f8085271",
          1329 => x"802e9038",
          1330 => x"72723482",
          1331 => x"8cf80881",
          1332 => x"05828cf8",
          1333 => x"0c8f3982",
          1334 => x"8cf00852",
          1335 => x"71802e85",
          1336 => x"38725171",
          1337 => x"2d843d0d",
          1338 => x"04fe3d0d",
          1339 => x"02970533",
          1340 => x"828cf008",
          1341 => x"76828cf0",
          1342 => x"0c5451ff",
          1343 => x"ad3f7282",
          1344 => x"8cf00c84",
          1345 => x"3d0d04fd",
          1346 => x"3d0d7554",
          1347 => x"73337081",
          1348 => x"ff065353",
          1349 => x"71802e8e",
          1350 => x"387281ff",
          1351 => x"06518114",
          1352 => x"54ff873f",
          1353 => x"e739853d",
          1354 => x"0d04fc3d",
          1355 => x"0d77828c",
          1356 => x"f0087882",
          1357 => x"8cf00c56",
          1358 => x"54733370",
          1359 => x"81ff0653",
          1360 => x"5371802e",
          1361 => x"8e387281",
          1362 => x"ff065181",
          1363 => x"1454feda",
          1364 => x"3fe73974",
          1365 => x"828cf00c",
          1366 => x"863d0d04",
          1367 => x"ec3d0d66",
          1368 => x"68595978",
          1369 => x"7081055a",
          1370 => x"33567580",
          1371 => x"2e84f838",
          1372 => x"75a52e09",
          1373 => x"810682de",
          1374 => x"3880707a",
          1375 => x"7081055c",
          1376 => x"33585b5b",
          1377 => x"75b02e09",
          1378 => x"81068538",
          1379 => x"815a8b39",
          1380 => x"75ad2e09",
          1381 => x"81068a38",
          1382 => x"825a7870",
          1383 => x"81055a33",
          1384 => x"5675aa2e",
          1385 => x"09810692",
          1386 => x"38778419",
          1387 => x"71087b70",
          1388 => x"81055d33",
          1389 => x"595d5953",
          1390 => x"9d39d016",
          1391 => x"53728926",
          1392 => x"95387a88",
          1393 => x"297b1005",
          1394 => x"7605d005",
          1395 => x"79708105",
          1396 => x"5b33575b",
          1397 => x"e5397580",
          1398 => x"ec327030",
          1399 => x"70720780",
          1400 => x"257880cc",
          1401 => x"32703070",
          1402 => x"72078025",
          1403 => x"73075354",
          1404 => x"58515553",
          1405 => x"73802e8c",
          1406 => x"38798407",
          1407 => x"79708105",
          1408 => x"5b33575a",
          1409 => x"75802e83",
          1410 => x"de387554",
          1411 => x"80e07627",
          1412 => x"8938e016",
          1413 => x"7081ff06",
          1414 => x"55537380",
          1415 => x"cf2e81aa",
          1416 => x"387380cf",
          1417 => x"24a23873",
          1418 => x"80c32e81",
          1419 => x"8e387380",
          1420 => x"c3248b38",
          1421 => x"7380c22e",
          1422 => x"818c3881",
          1423 => x"99397380",
          1424 => x"c42e818a",
          1425 => x"38818f39",
          1426 => x"7380d52e",
          1427 => x"81803873",
          1428 => x"80d5248a",
          1429 => x"387380d3",
          1430 => x"2e8e3880",
          1431 => x"f9397380",
          1432 => x"d82e80ee",
          1433 => x"3880ef39",
          1434 => x"77841971",
          1435 => x"08565953",
          1436 => x"80743354",
          1437 => x"5572752e",
          1438 => x"8d388115",
          1439 => x"70157033",
          1440 => x"51545572",
          1441 => x"f5387981",
          1442 => x"2a569039",
          1443 => x"74811656",
          1444 => x"53727b27",
          1445 => x"8f38a051",
          1446 => x"fc903f75",
          1447 => x"81065372",
          1448 => x"802ee938",
          1449 => x"7351fcdf",
          1450 => x"3f748116",
          1451 => x"5653727b",
          1452 => x"27fdb038",
          1453 => x"a051fbf2",
          1454 => x"3fef3977",
          1455 => x"84198312",
          1456 => x"33535953",
          1457 => x"9339825c",
          1458 => x"9539885c",
          1459 => x"91398a5c",
          1460 => x"8d39905c",
          1461 => x"89397551",
          1462 => x"fbd03ffd",
          1463 => x"86397982",
          1464 => x"2a708106",
          1465 => x"51537280",
          1466 => x"2e883877",
          1467 => x"84195953",
          1468 => x"86398418",
          1469 => x"78545872",
          1470 => x"087480c4",
          1471 => x"32703070",
          1472 => x"72078025",
          1473 => x"51555555",
          1474 => x"7480258d",
          1475 => x"3872802e",
          1476 => x"88387430",
          1477 => x"7a90075b",
          1478 => x"55800b8f",
          1479 => x"3d5e577b",
          1480 => x"527451dc",
          1481 => x"e93f828c",
          1482 => x"dc0881ff",
          1483 => x"067c5375",
          1484 => x"5254dca7",
          1485 => x"3f828cdc",
          1486 => x"08558974",
          1487 => x"279238a7",
          1488 => x"14537580",
          1489 => x"f82e8438",
          1490 => x"87145372",
          1491 => x"81ff0654",
          1492 => x"b0145372",
          1493 => x"7d708105",
          1494 => x"5f348117",
          1495 => x"75307077",
          1496 => x"079f2a51",
          1497 => x"5457769f",
          1498 => x"26853872",
          1499 => x"ffb13879",
          1500 => x"842a7081",
          1501 => x"06515372",
          1502 => x"802e8e38",
          1503 => x"963d7705",
          1504 => x"e00553ad",
          1505 => x"73348117",
          1506 => x"57767a81",
          1507 => x"065455b0",
          1508 => x"54728338",
          1509 => x"a0547981",
          1510 => x"2a708106",
          1511 => x"5456729f",
          1512 => x"38811755",
          1513 => x"767b2797",
          1514 => x"387351f9",
          1515 => x"fd3f7581",
          1516 => x"0653728b",
          1517 => x"38748116",
          1518 => x"56537a73",
          1519 => x"26eb3896",
          1520 => x"3d7705e0",
          1521 => x"0553ff17",
          1522 => x"ff147033",
          1523 => x"535457f9",
          1524 => x"d93f76f2",
          1525 => x"38748116",
          1526 => x"5653727b",
          1527 => x"27fb8438",
          1528 => x"a051f9c6",
          1529 => x"3fef3996",
          1530 => x"3d0d04fd",
          1531 => x"3d0d863d",
          1532 => x"70708405",
          1533 => x"52085552",
          1534 => x"7351fae0",
          1535 => x"3f853d0d",
          1536 => x"04fe3d0d",
          1537 => x"74828cf8",
          1538 => x"0c853d88",
          1539 => x"05527551",
          1540 => x"faca3f82",
          1541 => x"8cf80853",
          1542 => x"80733480",
          1543 => x"0b828cf8",
          1544 => x"0c843d0d",
          1545 => x"04fd3d0d",
          1546 => x"828cf008",
          1547 => x"76828cf0",
          1548 => x"0c873d88",
          1549 => x"05537752",
          1550 => x"53faa13f",
          1551 => x"72828cf0",
          1552 => x"0c853d0d",
          1553 => x"04fb3d0d",
          1554 => x"7779828c",
          1555 => x"f4087056",
          1556 => x"54575580",
          1557 => x"5471802e",
          1558 => x"80e03882",
          1559 => x"8cf40852",
          1560 => x"712d828c",
          1561 => x"dc0881ff",
          1562 => x"06537280",
          1563 => x"2e80cb38",
          1564 => x"728d2eb9",
          1565 => x"38728832",
          1566 => x"70307080",
          1567 => x"25515152",
          1568 => x"73802e8b",
          1569 => x"3871802e",
          1570 => x"8638ff14",
          1571 => x"5497399f",
          1572 => x"7325c838",
          1573 => x"ff165273",
          1574 => x"7225c038",
          1575 => x"74145272",
          1576 => x"72348114",
          1577 => x"547251f8",
          1578 => x"813fffaf",
          1579 => x"39731552",
          1580 => x"8072348a",
          1581 => x"51f7f33f",
          1582 => x"81537282",
          1583 => x"8cdc0c87",
          1584 => x"3d0d04fe",
          1585 => x"3d0d828c",
          1586 => x"f4087582",
          1587 => x"8cf40c77",
          1588 => x"53765253",
          1589 => x"feef3f72",
          1590 => x"828cf40c",
          1591 => x"843d0d04",
          1592 => x"f83d0d7a",
          1593 => x"7c5a5680",
          1594 => x"707a0c58",
          1595 => x"75087033",
          1596 => x"555373a0",
          1597 => x"2e098106",
          1598 => x"87388113",
          1599 => x"760ced39",
          1600 => x"73ad2e09",
          1601 => x"81068e38",
          1602 => x"81760811",
          1603 => x"770c7608",
          1604 => x"70335654",
          1605 => x"5873b02e",
          1606 => x"09810680",
          1607 => x"c2387508",
          1608 => x"8105760c",
          1609 => x"75087033",
          1610 => x"55537380",
          1611 => x"e22e8b38",
          1612 => x"90577380",
          1613 => x"f82e8538",
          1614 => x"8f398257",
          1615 => x"8113760c",
          1616 => x"75087033",
          1617 => x"5553ac39",
          1618 => x"8155a074",
          1619 => x"2780fa38",
          1620 => x"d0145380",
          1621 => x"55885789",
          1622 => x"73279838",
          1623 => x"80eb39d0",
          1624 => x"14538055",
          1625 => x"72892680",
          1626 => x"e0388639",
          1627 => x"805580d9",
          1628 => x"398a5780",
          1629 => x"55a07427",
          1630 => x"80c23880",
          1631 => x"e0742789",
          1632 => x"38e01470",
          1633 => x"81ff0655",
          1634 => x"53d01470",
          1635 => x"81ff0655",
          1636 => x"53907427",
          1637 => x"8e38f914",
          1638 => x"7081ff06",
          1639 => x"55538974",
          1640 => x"27ca3873",
          1641 => x"7727c538",
          1642 => x"74772914",
          1643 => x"76088105",
          1644 => x"770c7608",
          1645 => x"70335654",
          1646 => x"55ffba39",
          1647 => x"77802e84",
          1648 => x"38743055",
          1649 => x"74790c81",
          1650 => x"5574828c",
          1651 => x"dc0c8a3d",
          1652 => x"0d04f83d",
          1653 => x"0d7a7c5a",
          1654 => x"5680707a",
          1655 => x"0c587508",
          1656 => x"70335553",
          1657 => x"73a02e09",
          1658 => x"81068738",
          1659 => x"8113760c",
          1660 => x"ed3973ad",
          1661 => x"2e098106",
          1662 => x"8e388176",
          1663 => x"0811770c",
          1664 => x"76087033",
          1665 => x"56545873",
          1666 => x"b02e0981",
          1667 => x"0680c238",
          1668 => x"75088105",
          1669 => x"760c7508",
          1670 => x"70335553",
          1671 => x"7380e22e",
          1672 => x"8b389057",
          1673 => x"7380f82e",
          1674 => x"85388f39",
          1675 => x"82578113",
          1676 => x"760c7508",
          1677 => x"70335553",
          1678 => x"ac398155",
          1679 => x"a0742780",
          1680 => x"fa38d014",
          1681 => x"53805588",
          1682 => x"57897327",
          1683 => x"983880eb",
          1684 => x"39d01453",
          1685 => x"80557289",
          1686 => x"2680e038",
          1687 => x"86398055",
          1688 => x"80d9398a",
          1689 => x"578055a0",
          1690 => x"742780c2",
          1691 => x"3880e074",
          1692 => x"278938e0",
          1693 => x"147081ff",
          1694 => x"065553d0",
          1695 => x"147081ff",
          1696 => x"06555390",
          1697 => x"74278e38",
          1698 => x"f9147081",
          1699 => x"ff065553",
          1700 => x"897427ca",
          1701 => x"38737727",
          1702 => x"c5387477",
          1703 => x"29147608",
          1704 => x"8105770c",
          1705 => x"76087033",
          1706 => x"565455ff",
          1707 => x"ba397780",
          1708 => x"2e843874",
          1709 => x"30557479",
          1710 => x"0c815574",
          1711 => x"828cdc0c",
          1712 => x"8a3d0d04",
          1713 => x"fd3d0d76",
          1714 => x"982b7098",
          1715 => x"2c79982b",
          1716 => x"70982c72",
          1717 => x"10137082",
          1718 => x"2b515351",
          1719 => x"54515180",
          1720 => x"0b81f8dc",
          1721 => x"12335553",
          1722 => x"7174259c",
          1723 => x"3881f8d8",
          1724 => x"11081202",
          1725 => x"84059705",
          1726 => x"33713352",
          1727 => x"52527072",
          1728 => x"2e098106",
          1729 => x"83388153",
          1730 => x"72828cdc",
          1731 => x"0c853d0d",
          1732 => x"04fc3d0d",
          1733 => x"78028405",
          1734 => x"9f053371",
          1735 => x"33545553",
          1736 => x"71802e9f",
          1737 => x"388851f3",
          1738 => x"813fa051",
          1739 => x"f2fc3f88",
          1740 => x"51f2f73f",
          1741 => x"7233ff05",
          1742 => x"52717334",
          1743 => x"7181ff06",
          1744 => x"52de3976",
          1745 => x"51f3c03f",
          1746 => x"73733486",
          1747 => x"3d0d04f6",
          1748 => x"3d0d7c02",
          1749 => x"8405b705",
          1750 => x"33028805",
          1751 => x"bb053382",
          1752 => x"89a83370",
          1753 => x"84298288",
          1754 => x"d0057008",
          1755 => x"5159595a",
          1756 => x"58597480",
          1757 => x"2e863874",
          1758 => x"51f29b3f",
          1759 => x"8289a833",
          1760 => x"70842982",
          1761 => x"88d00581",
          1762 => x"19705458",
          1763 => x"565af0bc",
          1764 => x"3f828cdc",
          1765 => x"08750c82",
          1766 => x"89a83370",
          1767 => x"84298288",
          1768 => x"d0057008",
          1769 => x"51565a74",
          1770 => x"802ea638",
          1771 => x"75537852",
          1772 => x"7451d69f",
          1773 => x"3f8289a8",
          1774 => x"33810555",
          1775 => x"748289a8",
          1776 => x"347481ff",
          1777 => x"06559375",
          1778 => x"27873880",
          1779 => x"0b8289a8",
          1780 => x"3477802e",
          1781 => x"b6388289",
          1782 => x"a4085675",
          1783 => x"802eac38",
          1784 => x"8289a033",
          1785 => x"5574a438",
          1786 => x"8c3dfc05",
          1787 => x"54765378",
          1788 => x"52755180",
          1789 => x"c8913f82",
          1790 => x"89a40852",
          1791 => x"8a5180fd",
          1792 => x"9e3f8289",
          1793 => x"a4085180",
          1794 => x"cbee3f8c",
          1795 => x"3d0d04dc",
          1796 => x"3d0d8157",
          1797 => x"80528289",
          1798 => x"a4085180",
          1799 => x"d2873f82",
          1800 => x"8cdc0880",
          1801 => x"d1388289",
          1802 => x"a4085380",
          1803 => x"f852883d",
          1804 => x"70525680",
          1805 => x"fad53f82",
          1806 => x"8cdc0880",
          1807 => x"2eb83875",
          1808 => x"51d8ab3f",
          1809 => x"828cdc08",
          1810 => x"55800b82",
          1811 => x"8cdc0825",
          1812 => x"9c38828c",
          1813 => x"dc08ff05",
          1814 => x"70175555",
          1815 => x"80743475",
          1816 => x"53765281",
          1817 => x"1781f7f0",
          1818 => x"5257f6ff",
          1819 => x"3f74ff2e",
          1820 => x"098106ff",
          1821 => x"b138a63d",
          1822 => x"0d04d93d",
          1823 => x"0daa3d08",
          1824 => x"ad3d085a",
          1825 => x"5a817058",
          1826 => x"58805282",
          1827 => x"89a40851",
          1828 => x"80d1923f",
          1829 => x"828cdc08",
          1830 => x"819138ff",
          1831 => x"0b8289a4",
          1832 => x"08545580",
          1833 => x"f8528b3d",
          1834 => x"70525680",
          1835 => x"f9dd3f82",
          1836 => x"8cdc0880",
          1837 => x"2ea43875",
          1838 => x"51d7b33f",
          1839 => x"828cdc08",
          1840 => x"81185855",
          1841 => x"800b828c",
          1842 => x"dc08258e",
          1843 => x"38828cdc",
          1844 => x"08ff0570",
          1845 => x"17555580",
          1846 => x"74347409",
          1847 => x"70307072",
          1848 => x"079f2a51",
          1849 => x"55557877",
          1850 => x"2e853873",
          1851 => x"ffad3882",
          1852 => x"89a4088c",
          1853 => x"11085351",
          1854 => x"80d0aa3f",
          1855 => x"828cdc08",
          1856 => x"802e8838",
          1857 => x"81f7fc51",
          1858 => x"effd3f78",
          1859 => x"772e0981",
          1860 => x"06993875",
          1861 => x"527951d5",
          1862 => x"e63f7951",
          1863 => x"d6d03fab",
          1864 => x"3d085482",
          1865 => x"8cdc0874",
          1866 => x"34805877",
          1867 => x"828cdc0c",
          1868 => x"a93d0d04",
          1869 => x"f63d0d7c",
          1870 => x"7e715c71",
          1871 => x"72335759",
          1872 => x"5a5873a0",
          1873 => x"2e098106",
          1874 => x"a2387833",
          1875 => x"78055677",
          1876 => x"76279838",
          1877 => x"8117705b",
          1878 => x"70713356",
          1879 => x"585573a0",
          1880 => x"2e098106",
          1881 => x"86387575",
          1882 => x"26ea3880",
          1883 => x"54738829",
          1884 => x"8289ac05",
          1885 => x"70085255",
          1886 => x"d5f43f82",
          1887 => x"8cdc0853",
          1888 => x"79527408",
          1889 => x"51d6c83f",
          1890 => x"828cdc08",
          1891 => x"80c43884",
          1892 => x"15335574",
          1893 => x"812e8838",
          1894 => x"74822e88",
          1895 => x"38b439fc",
          1896 => x"ee3fab39",
          1897 => x"811a5a8c",
          1898 => x"3dfc1153",
          1899 => x"f80551f6",
          1900 => x"af3f828c",
          1901 => x"dc08802e",
          1902 => x"99387a53",
          1903 => x"78527751",
          1904 => x"fdb83f82",
          1905 => x"8cdc0881",
          1906 => x"ff065574",
          1907 => x"85387454",
          1908 => x"91398114",
          1909 => x"7081ff06",
          1910 => x"51548274",
          1911 => x"27ff8e38",
          1912 => x"80547382",
          1913 => x"8cdc0c8c",
          1914 => x"3d0d04d3",
          1915 => x"3d0db03d",
          1916 => x"08028405",
          1917 => x"81c30533",
          1918 => x"5f5a800b",
          1919 => x"af3d3482",
          1920 => x"89a8335b",
          1921 => x"8289a408",
          1922 => x"81a33882",
          1923 => x"89a03354",
          1924 => x"73819a38",
          1925 => x"a851ebb4",
          1926 => x"3f828cdc",
          1927 => x"088289a4",
          1928 => x"0c828cdc",
          1929 => x"08802e80",
          1930 => x"fe389353",
          1931 => x"8288cc08",
          1932 => x"52828cdc",
          1933 => x"0851bbed",
          1934 => x"3f828cdc",
          1935 => x"08802e8b",
          1936 => x"3881f8a8",
          1937 => x"51f3a43f",
          1938 => x"80e33982",
          1939 => x"89a40853",
          1940 => x"80f85290",
          1941 => x"3d705254",
          1942 => x"80f6b03f",
          1943 => x"828cdc08",
          1944 => x"56828cdc",
          1945 => x"08742e09",
          1946 => x"810680c1",
          1947 => x"38828cdc",
          1948 => x"0851d3fa",
          1949 => x"3f828cdc",
          1950 => x"0855800b",
          1951 => x"828cdc08",
          1952 => x"259a3882",
          1953 => x"8cdc08ff",
          1954 => x"05701755",
          1955 => x"55807434",
          1956 => x"80537481",
          1957 => x"ff065275",
          1958 => x"51f9b43f",
          1959 => x"74ff2e09",
          1960 => x"8106ffa7",
          1961 => x"38873981",
          1962 => x"0b8289a0",
          1963 => x"348f3d5d",
          1964 => x"ddcc3f82",
          1965 => x"8cdc0898",
          1966 => x"2b70982c",
          1967 => x"515978ff",
          1968 => x"2eee3878",
          1969 => x"81ff0682",
          1970 => x"8d803370",
          1971 => x"982b7098",
          1972 => x"2c828cfc",
          1973 => x"3370982b",
          1974 => x"70972c71",
          1975 => x"982c0570",
          1976 => x"842981f8",
          1977 => x"d8057008",
          1978 => x"15703351",
          1979 => x"51515159",
          1980 => x"5951595d",
          1981 => x"58815673",
          1982 => x"782e80e9",
          1983 => x"38777427",
          1984 => x"b4387481",
          1985 => x"800a2981",
          1986 => x"ff0a0570",
          1987 => x"982c5155",
          1988 => x"80752480",
          1989 => x"ce387653",
          1990 => x"74527751",
          1991 => x"f7a63f82",
          1992 => x"8cdc0881",
          1993 => x"ff065473",
          1994 => x"802ed738",
          1995 => x"74828cfc",
          1996 => x"348156b1",
          1997 => x"39748180",
          1998 => x"0a298180",
          1999 => x"0a057098",
          2000 => x"2c7081ff",
          2001 => x"06565155",
          2002 => x"738a2697",
          2003 => x"38765374",
          2004 => x"527751f6",
          2005 => x"ef3f828c",
          2006 => x"dc0881ff",
          2007 => x"065473cc",
          2008 => x"38d33980",
          2009 => x"5675802e",
          2010 => x"80ca3881",
          2011 => x"1c557482",
          2012 => x"8d803474",
          2013 => x"982b7098",
          2014 => x"2c828cfc",
          2015 => x"3370982b",
          2016 => x"70982c70",
          2017 => x"10117082",
          2018 => x"2b81f8dc",
          2019 => x"11335e51",
          2020 => x"51515758",
          2021 => x"51557477",
          2022 => x"2e098106",
          2023 => x"fe923881",
          2024 => x"f8e01408",
          2025 => x"7d0c800b",
          2026 => x"828d8034",
          2027 => x"800b828c",
          2028 => x"fc349239",
          2029 => x"75828d80",
          2030 => x"3475828c",
          2031 => x"fc3478af",
          2032 => x"3d34757d",
          2033 => x"0c7e5473",
          2034 => x"8b26fde1",
          2035 => x"38738429",
          2036 => x"81f0e405",
          2037 => x"54730804",
          2038 => x"828d8833",
          2039 => x"54737e2e",
          2040 => x"fdcb3882",
          2041 => x"8d843355",
          2042 => x"737527ab",
          2043 => x"3874982b",
          2044 => x"70982c51",
          2045 => x"55737524",
          2046 => x"9e38741a",
          2047 => x"54733381",
          2048 => x"15347481",
          2049 => x"800a2981",
          2050 => x"ff0a0570",
          2051 => x"982c828d",
          2052 => x"88335651",
          2053 => x"55df3982",
          2054 => x"8d883381",
          2055 => x"11565474",
          2056 => x"828d8834",
          2057 => x"731a54ae",
          2058 => x"3d337434",
          2059 => x"828d8433",
          2060 => x"54737e27",
          2061 => x"89388114",
          2062 => x"5473828d",
          2063 => x"8434828d",
          2064 => x"88337081",
          2065 => x"800a2981",
          2066 => x"ff0a0570",
          2067 => x"982c828d",
          2068 => x"84335a51",
          2069 => x"56567477",
          2070 => x"25a23874",
          2071 => x"1a703352",
          2072 => x"54e8c73f",
          2073 => x"7481800a",
          2074 => x"2981800a",
          2075 => x"0570982c",
          2076 => x"828d8433",
          2077 => x"56515573",
          2078 => x"7524e038",
          2079 => x"828d8833",
          2080 => x"70982b70",
          2081 => x"982c828d",
          2082 => x"84335a51",
          2083 => x"56567477",
          2084 => x"25fc9a38",
          2085 => x"8851e892",
          2086 => x"3f748180",
          2087 => x"0a298180",
          2088 => x"0a057098",
          2089 => x"2c828d84",
          2090 => x"33565155",
          2091 => x"737524e4",
          2092 => x"38fbfa39",
          2093 => x"828d8833",
          2094 => x"7081ff06",
          2095 => x"55557380",
          2096 => x"2efbea38",
          2097 => x"828d8433",
          2098 => x"ff055473",
          2099 => x"828d8434",
          2100 => x"ff155473",
          2101 => x"828d8834",
          2102 => x"8851e7ce",
          2103 => x"3f828d88",
          2104 => x"3370982b",
          2105 => x"70982c82",
          2106 => x"8d843357",
          2107 => x"51565774",
          2108 => x"7425a738",
          2109 => x"741a5481",
          2110 => x"14337434",
          2111 => x"733351e7",
          2112 => x"a93f7481",
          2113 => x"800a2981",
          2114 => x"800a0570",
          2115 => x"982c828d",
          2116 => x"84335851",
          2117 => x"55757524",
          2118 => x"db38a051",
          2119 => x"e78c3f82",
          2120 => x"8d883370",
          2121 => x"982b7098",
          2122 => x"2c828d84",
          2123 => x"33575156",
          2124 => x"57747424",
          2125 => x"faf73888",
          2126 => x"51e6ef3f",
          2127 => x"7481800a",
          2128 => x"2981800a",
          2129 => x"0570982c",
          2130 => x"828d8433",
          2131 => x"58515575",
          2132 => x"7525e438",
          2133 => x"fad73982",
          2134 => x"8d84337a",
          2135 => x"05548074",
          2136 => x"348a51e6",
          2137 => x"c53f828d",
          2138 => x"84527951",
          2139 => x"f7c63f82",
          2140 => x"8cdc0881",
          2141 => x"ff065473",
          2142 => x"9838828d",
          2143 => x"84335473",
          2144 => x"802e84c9",
          2145 => x"38815373",
          2146 => x"527951f3",
          2147 => x"c23f84bd",
          2148 => x"39807a34",
          2149 => x"84b73982",
          2150 => x"8d883354",
          2151 => x"73802efa",
          2152 => x"8c388851",
          2153 => x"e6843f82",
          2154 => x"8d8833ff",
          2155 => x"05547382",
          2156 => x"8d883473",
          2157 => x"81ff0654",
          2158 => x"e339828d",
          2159 => x"8833828d",
          2160 => x"84335555",
          2161 => x"73752ef9",
          2162 => x"e438ff14",
          2163 => x"5473828d",
          2164 => x"84347498",
          2165 => x"2b70982c",
          2166 => x"7581ff06",
          2167 => x"56515574",
          2168 => x"7425a738",
          2169 => x"741a5481",
          2170 => x"14337434",
          2171 => x"733351e5",
          2172 => x"b93f7481",
          2173 => x"800a2981",
          2174 => x"800a0570",
          2175 => x"982c828d",
          2176 => x"84335851",
          2177 => x"55757524",
          2178 => x"db38a051",
          2179 => x"e59c3f82",
          2180 => x"8d883370",
          2181 => x"982b7098",
          2182 => x"2c828d84",
          2183 => x"33575156",
          2184 => x"57747424",
          2185 => x"f9873888",
          2186 => x"51e4ff3f",
          2187 => x"7481800a",
          2188 => x"2981800a",
          2189 => x"0570982c",
          2190 => x"828d8433",
          2191 => x"58515575",
          2192 => x"7525e438",
          2193 => x"f8e73982",
          2194 => x"8d883370",
          2195 => x"81ff0682",
          2196 => x"8d843359",
          2197 => x"56547477",
          2198 => x"27f8d238",
          2199 => x"81145473",
          2200 => x"828d8834",
          2201 => x"741a7033",
          2202 => x"5254e4be",
          2203 => x"3f828d88",
          2204 => x"337081ff",
          2205 => x"06828d84",
          2206 => x"33585654",
          2207 => x"757526dc",
          2208 => x"38f8aa39",
          2209 => x"7aae3882",
          2210 => x"899c0855",
          2211 => x"74802ea4",
          2212 => x"387451cb",
          2213 => x"d93f828c",
          2214 => x"dc08828d",
          2215 => x"8434828c",
          2216 => x"dc0881ff",
          2217 => x"06810553",
          2218 => x"74527951",
          2219 => x"c8a53f93",
          2220 => x"5b81c139",
          2221 => x"7a842982",
          2222 => x"88d005fc",
          2223 => x"11085654",
          2224 => x"74802ea5",
          2225 => x"387451cb",
          2226 => x"a53f828c",
          2227 => x"dc08828d",
          2228 => x"8434828c",
          2229 => x"dc0881ff",
          2230 => x"06810553",
          2231 => x"74527951",
          2232 => x"c7f13fff",
          2233 => x"1b5480de",
          2234 => x"39730855",
          2235 => x"74802ef7",
          2236 => x"bc387451",
          2237 => x"caf83f80",
          2238 => x"e2397a93",
          2239 => x"2e098106",
          2240 => x"93388288",
          2241 => x"d0085574",
          2242 => x"802e8938",
          2243 => x"7451cade",
          2244 => x"3f80c839",
          2245 => x"7a842982",
          2246 => x"88d00584",
          2247 => x"11085654",
          2248 => x"74802ea9",
          2249 => x"387451ca",
          2250 => x"c53f828c",
          2251 => x"dc08828d",
          2252 => x"8434828c",
          2253 => x"dc0881ff",
          2254 => x"06810553",
          2255 => x"74527951",
          2256 => x"c7913f81",
          2257 => x"1b547381",
          2258 => x"ff065ba8",
          2259 => x"39730855",
          2260 => x"74802ef6",
          2261 => x"d8387451",
          2262 => x"ca943f82",
          2263 => x"8cdc0882",
          2264 => x"8d843482",
          2265 => x"8cdc0881",
          2266 => x"ff068105",
          2267 => x"53745279",
          2268 => x"51c6e03f",
          2269 => x"828d8853",
          2270 => x"828d8433",
          2271 => x"527951ef",
          2272 => x"903ff6a9",
          2273 => x"39828d88",
          2274 => x"337081ff",
          2275 => x"06828d84",
          2276 => x"33595654",
          2277 => x"747727f6",
          2278 => x"94388114",
          2279 => x"5473828d",
          2280 => x"8834741a",
          2281 => x"70335254",
          2282 => x"e2803ff6",
          2283 => x"8039828d",
          2284 => x"88335473",
          2285 => x"802ef5f5",
          2286 => x"388851e1",
          2287 => x"ed3f828d",
          2288 => x"8833ff05",
          2289 => x"5473828d",
          2290 => x"8834f5e1",
          2291 => x"39800b82",
          2292 => x"8d883480",
          2293 => x"0b828d84",
          2294 => x"3479828c",
          2295 => x"dc0caf3d",
          2296 => x"0d04ff3d",
          2297 => x"0d028f05",
          2298 => x"33518152",
          2299 => x"70722687",
          2300 => x"388289c4",
          2301 => x"11335271",
          2302 => x"828cdc0c",
          2303 => x"833d0d04",
          2304 => x"fc3d0d02",
          2305 => x"9b053302",
          2306 => x"84059f05",
          2307 => x"33565383",
          2308 => x"51728126",
          2309 => x"80e03872",
          2310 => x"842b87c0",
          2311 => x"928c1153",
          2312 => x"51885474",
          2313 => x"802e8438",
          2314 => x"81885473",
          2315 => x"720c87c0",
          2316 => x"928c1151",
          2317 => x"81710c85",
          2318 => x"0b87c098",
          2319 => x"8c0c7052",
          2320 => x"71087082",
          2321 => x"06515170",
          2322 => x"802e8a38",
          2323 => x"87c0988c",
          2324 => x"085170ec",
          2325 => x"387108fc",
          2326 => x"80800652",
          2327 => x"71923887",
          2328 => x"c0988c08",
          2329 => x"5170802e",
          2330 => x"87387182",
          2331 => x"89c41434",
          2332 => x"8289c413",
          2333 => x"33517082",
          2334 => x"8cdc0c86",
          2335 => x"3d0d04f3",
          2336 => x"3d0d6062",
          2337 => x"64028c05",
          2338 => x"bf053357",
          2339 => x"40585b83",
          2340 => x"74525afe",
          2341 => x"cd3f828c",
          2342 => x"dc088106",
          2343 => x"7a545271",
          2344 => x"81be3871",
          2345 => x"7275842b",
          2346 => x"87c09280",
          2347 => x"1187c092",
          2348 => x"8c1287c0",
          2349 => x"92841341",
          2350 => x"5a40575a",
          2351 => x"58850b87",
          2352 => x"c0988c0c",
          2353 => x"767d0c84",
          2354 => x"760c7508",
          2355 => x"70852a70",
          2356 => x"81065153",
          2357 => x"5471802e",
          2358 => x"8e387b08",
          2359 => x"52717b70",
          2360 => x"81055d34",
          2361 => x"81195980",
          2362 => x"74a20653",
          2363 => x"5371732e",
          2364 => x"83388153",
          2365 => x"7883ff26",
          2366 => x"8f387280",
          2367 => x"2e8a3887",
          2368 => x"c0988c08",
          2369 => x"5271c338",
          2370 => x"87c0988c",
          2371 => x"08527180",
          2372 => x"2e873878",
          2373 => x"84802e99",
          2374 => x"3881760c",
          2375 => x"87c0928c",
          2376 => x"15537208",
          2377 => x"70820651",
          2378 => x"5271f738",
          2379 => x"ff1a5a8d",
          2380 => x"39848017",
          2381 => x"81197081",
          2382 => x"ff065a53",
          2383 => x"5779802e",
          2384 => x"903873fc",
          2385 => x"80800652",
          2386 => x"7187387d",
          2387 => x"7826feed",
          2388 => x"3873fc80",
          2389 => x"80065271",
          2390 => x"802e8338",
          2391 => x"81527153",
          2392 => x"72828cdc",
          2393 => x"0c8f3d0d",
          2394 => x"04f33d0d",
          2395 => x"60626402",
          2396 => x"8c05bf05",
          2397 => x"33574058",
          2398 => x"5b835980",
          2399 => x"745258fc",
          2400 => x"e13f828c",
          2401 => x"dc088106",
          2402 => x"79545271",
          2403 => x"782e0981",
          2404 => x"0681b138",
          2405 => x"7774842b",
          2406 => x"87c09280",
          2407 => x"1187c092",
          2408 => x"8c1287c0",
          2409 => x"92841340",
          2410 => x"595f565a",
          2411 => x"850b87c0",
          2412 => x"988c0c76",
          2413 => x"7d0c8276",
          2414 => x"0c805875",
          2415 => x"0870842a",
          2416 => x"70810651",
          2417 => x"53547180",
          2418 => x"2e8c387a",
          2419 => x"7081055c",
          2420 => x"337c0c81",
          2421 => x"18587381",
          2422 => x"2a708106",
          2423 => x"51527180",
          2424 => x"2e8a3887",
          2425 => x"c0988c08",
          2426 => x"5271d038",
          2427 => x"87c0988c",
          2428 => x"08527180",
          2429 => x"2e873877",
          2430 => x"84802e99",
          2431 => x"3881760c",
          2432 => x"87c0928c",
          2433 => x"15537208",
          2434 => x"70820651",
          2435 => x"5271f738",
          2436 => x"ff19598d",
          2437 => x"39811a70",
          2438 => x"81ff0684",
          2439 => x"8019595b",
          2440 => x"5278802e",
          2441 => x"903873fc",
          2442 => x"80800652",
          2443 => x"7187387d",
          2444 => x"7a26fef8",
          2445 => x"3873fc80",
          2446 => x"80065271",
          2447 => x"802e8338",
          2448 => x"81527153",
          2449 => x"72828cdc",
          2450 => x"0c8f3d0d",
          2451 => x"04fa3d0d",
          2452 => x"7a028405",
          2453 => x"a3053302",
          2454 => x"8805a705",
          2455 => x"33715454",
          2456 => x"5657fafe",
          2457 => x"3f828cdc",
          2458 => x"08810653",
          2459 => x"83547280",
          2460 => x"fe38850b",
          2461 => x"87c0988c",
          2462 => x"0c815671",
          2463 => x"762e80dc",
          2464 => x"38717624",
          2465 => x"93387484",
          2466 => x"2b87c092",
          2467 => x"8c115454",
          2468 => x"71802e8d",
          2469 => x"3880d439",
          2470 => x"71832e80",
          2471 => x"c63880cb",
          2472 => x"39720870",
          2473 => x"812a7081",
          2474 => x"06515152",
          2475 => x"71802e8a",
          2476 => x"3887c098",
          2477 => x"8c085271",
          2478 => x"e83887c0",
          2479 => x"988c0852",
          2480 => x"71963881",
          2481 => x"730c87c0",
          2482 => x"928c1453",
          2483 => x"72087082",
          2484 => x"06515271",
          2485 => x"f7389639",
          2486 => x"80569239",
          2487 => x"88800a77",
          2488 => x"0c853981",
          2489 => x"80770c72",
          2490 => x"56833984",
          2491 => x"56755473",
          2492 => x"828cdc0c",
          2493 => x"883d0d04",
          2494 => x"fe3d0d74",
          2495 => x"81113371",
          2496 => x"3371882b",
          2497 => x"07828cdc",
          2498 => x"0c535184",
          2499 => x"3d0d04fd",
          2500 => x"3d0d7583",
          2501 => x"11338212",
          2502 => x"3371902b",
          2503 => x"71882b07",
          2504 => x"81143370",
          2505 => x"7207882b",
          2506 => x"75337107",
          2507 => x"828cdc0c",
          2508 => x"52535456",
          2509 => x"5452853d",
          2510 => x"0d04ff3d",
          2511 => x"0d730284",
          2512 => x"05920522",
          2513 => x"52527072",
          2514 => x"70810554",
          2515 => x"3470882a",
          2516 => x"51707234",
          2517 => x"833d0d04",
          2518 => x"ff3d0d73",
          2519 => x"75525270",
          2520 => x"72708105",
          2521 => x"54347088",
          2522 => x"2a517072",
          2523 => x"70810554",
          2524 => x"3470882a",
          2525 => x"51707270",
          2526 => x"81055434",
          2527 => x"70882a51",
          2528 => x"70723483",
          2529 => x"3d0d04fe",
          2530 => x"3d0d7675",
          2531 => x"77545451",
          2532 => x"70802e92",
          2533 => x"38717081",
          2534 => x"05533373",
          2535 => x"70810555",
          2536 => x"34ff1151",
          2537 => x"eb39843d",
          2538 => x"0d04fe3d",
          2539 => x"0d757776",
          2540 => x"54525372",
          2541 => x"72708105",
          2542 => x"5434ff11",
          2543 => x"5170f438",
          2544 => x"843d0d04",
          2545 => x"fc3d0d78",
          2546 => x"77795656",
          2547 => x"53747081",
          2548 => x"05563374",
          2549 => x"70810556",
          2550 => x"33717131",
          2551 => x"ff165652",
          2552 => x"52527280",
          2553 => x"2e863871",
          2554 => x"802ee238",
          2555 => x"71828cdc",
          2556 => x"0c863d0d",
          2557 => x"04fe3d0d",
          2558 => x"74765451",
          2559 => x"89397173",
          2560 => x"2e8a3881",
          2561 => x"11517033",
          2562 => x"5271f338",
          2563 => x"7033828c",
          2564 => x"dc0c843d",
          2565 => x"0d04800b",
          2566 => x"828cdc0c",
          2567 => x"04800b82",
          2568 => x"8cdc0c04",
          2569 => x"f73d0d7b",
          2570 => x"56800b83",
          2571 => x"1733565a",
          2572 => x"747a2e80",
          2573 => x"d6388154",
          2574 => x"b0160853",
          2575 => x"b4167053",
          2576 => x"81173352",
          2577 => x"59faa23f",
          2578 => x"828cdc08",
          2579 => x"7a2e0981",
          2580 => x"06b73882",
          2581 => x"8cdc0883",
          2582 => x"1734b016",
          2583 => x"0870a418",
          2584 => x"08319c18",
          2585 => x"08595658",
          2586 => x"7477279f",
          2587 => x"38821633",
          2588 => x"5574822e",
          2589 => x"09810693",
          2590 => x"38815476",
          2591 => x"18537852",
          2592 => x"81163351",
          2593 => x"f9e33f83",
          2594 => x"39815a79",
          2595 => x"828cdc0c",
          2596 => x"8b3d0d04",
          2597 => x"fa3d0d78",
          2598 => x"7a565680",
          2599 => x"5774b017",
          2600 => x"082eaf38",
          2601 => x"7551fefc",
          2602 => x"3f828cdc",
          2603 => x"0857828c",
          2604 => x"dc089f38",
          2605 => x"81547453",
          2606 => x"b4165281",
          2607 => x"163351f7",
          2608 => x"be3f828c",
          2609 => x"dc08802e",
          2610 => x"8538ff55",
          2611 => x"815774b0",
          2612 => x"170c7682",
          2613 => x"8cdc0c88",
          2614 => x"3d0d04f8",
          2615 => x"3d0d7a70",
          2616 => x"5257fec0",
          2617 => x"3f828cdc",
          2618 => x"0858828c",
          2619 => x"dc088191",
          2620 => x"38763355",
          2621 => x"74832e09",
          2622 => x"810680f0",
          2623 => x"38841733",
          2624 => x"5978812e",
          2625 => x"09810680",
          2626 => x"e3388480",
          2627 => x"53828cdc",
          2628 => x"0852b417",
          2629 => x"705256fd",
          2630 => x"913f82d4",
          2631 => x"d55284b2",
          2632 => x"1751fc96",
          2633 => x"3f848b85",
          2634 => x"a4d25275",
          2635 => x"51fca93f",
          2636 => x"868a85e4",
          2637 => x"f2528498",
          2638 => x"1751fc9c",
          2639 => x"3f901708",
          2640 => x"52849c17",
          2641 => x"51fc913f",
          2642 => x"8c170852",
          2643 => x"84a01751",
          2644 => x"fc863fa0",
          2645 => x"17088105",
          2646 => x"70b0190c",
          2647 => x"79555375",
          2648 => x"52811733",
          2649 => x"51f8823f",
          2650 => x"77841834",
          2651 => x"80538052",
          2652 => x"81173351",
          2653 => x"f9d73f82",
          2654 => x"8cdc0880",
          2655 => x"2e833881",
          2656 => x"5877828c",
          2657 => x"dc0c8a3d",
          2658 => x"0d04fb3d",
          2659 => x"0d77fe1a",
          2660 => x"981208fe",
          2661 => x"05555654",
          2662 => x"80567473",
          2663 => x"278d388a",
          2664 => x"14227571",
          2665 => x"29ac1608",
          2666 => x"05575375",
          2667 => x"828cdc0c",
          2668 => x"873d0d04",
          2669 => x"f93d0d7a",
          2670 => x"7a700856",
          2671 => x"54578177",
          2672 => x"2781df38",
          2673 => x"76981508",
          2674 => x"2781d738",
          2675 => x"ff743354",
          2676 => x"5872822e",
          2677 => x"80f53872",
          2678 => x"82248938",
          2679 => x"72812e8d",
          2680 => x"3881bf39",
          2681 => x"72832e81",
          2682 => x"8e3881b6",
          2683 => x"3976812a",
          2684 => x"1770892a",
          2685 => x"a4160805",
          2686 => x"53745255",
          2687 => x"fd963f82",
          2688 => x"8cdc0881",
          2689 => x"9f387483",
          2690 => x"ff0614b4",
          2691 => x"11338117",
          2692 => x"70892aa4",
          2693 => x"18080555",
          2694 => x"76545757",
          2695 => x"53fcf53f",
          2696 => x"828cdc08",
          2697 => x"80fe3874",
          2698 => x"83ff0614",
          2699 => x"b4113370",
          2700 => x"882b7807",
          2701 => x"79810671",
          2702 => x"842a5c52",
          2703 => x"58515372",
          2704 => x"80e23875",
          2705 => x"9fff0658",
          2706 => x"80da3976",
          2707 => x"882aa415",
          2708 => x"08055273",
          2709 => x"51fcbd3f",
          2710 => x"828cdc08",
          2711 => x"80c63876",
          2712 => x"1083fe06",
          2713 => x"7405b405",
          2714 => x"51f98d3f",
          2715 => x"828cdc08",
          2716 => x"83ffff06",
          2717 => x"58ae3976",
          2718 => x"872aa415",
          2719 => x"08055273",
          2720 => x"51fc913f",
          2721 => x"828cdc08",
          2722 => x"9b387682",
          2723 => x"2b83fc06",
          2724 => x"7405b405",
          2725 => x"51f8f83f",
          2726 => x"828cdc08",
          2727 => x"f00a0658",
          2728 => x"83398158",
          2729 => x"77828cdc",
          2730 => x"0c893d0d",
          2731 => x"04f83d0d",
          2732 => x"7a7c7e5a",
          2733 => x"58568259",
          2734 => x"81772782",
          2735 => x"9e387698",
          2736 => x"17082782",
          2737 => x"96387533",
          2738 => x"5372792e",
          2739 => x"819d3872",
          2740 => x"79248938",
          2741 => x"72812e8d",
          2742 => x"38828039",
          2743 => x"72832e81",
          2744 => x"b83881f7",
          2745 => x"3976812a",
          2746 => x"1770892a",
          2747 => x"a4180805",
          2748 => x"53765255",
          2749 => x"fb9e3f82",
          2750 => x"8cdc0859",
          2751 => x"828cdc08",
          2752 => x"81d93874",
          2753 => x"83ff0616",
          2754 => x"b4058116",
          2755 => x"78810659",
          2756 => x"56547753",
          2757 => x"76802e8f",
          2758 => x"3877842b",
          2759 => x"9ff00674",
          2760 => x"338f0671",
          2761 => x"07515372",
          2762 => x"7434810b",
          2763 => x"83173474",
          2764 => x"892aa417",
          2765 => x"08055275",
          2766 => x"51fad93f",
          2767 => x"828cdc08",
          2768 => x"59828cdc",
          2769 => x"08819438",
          2770 => x"7483ff06",
          2771 => x"16b40578",
          2772 => x"842a5454",
          2773 => x"768f3877",
          2774 => x"882a7433",
          2775 => x"81f00671",
          2776 => x"8f060751",
          2777 => x"53727434",
          2778 => x"80ec3976",
          2779 => x"882aa417",
          2780 => x"08055275",
          2781 => x"51fa9d3f",
          2782 => x"828cdc08",
          2783 => x"59828cdc",
          2784 => x"0880d838",
          2785 => x"7783ffff",
          2786 => x"06527610",
          2787 => x"83fe0676",
          2788 => x"05b40551",
          2789 => x"f7a43fbe",
          2790 => x"3976872a",
          2791 => x"a4170805",
          2792 => x"527551f9",
          2793 => x"ef3f828c",
          2794 => x"dc085982",
          2795 => x"8cdc08ab",
          2796 => x"3877f00a",
          2797 => x"0677822b",
          2798 => x"83fc0670",
          2799 => x"18b40570",
          2800 => x"54515454",
          2801 => x"f6c93f82",
          2802 => x"8cdc088f",
          2803 => x"0a067407",
          2804 => x"527251f7",
          2805 => x"833f810b",
          2806 => x"83173478",
          2807 => x"828cdc0c",
          2808 => x"8a3d0d04",
          2809 => x"f83d0d7a",
          2810 => x"7c7e7208",
          2811 => x"59565659",
          2812 => x"817527a4",
          2813 => x"38749817",
          2814 => x"08279d38",
          2815 => x"73802eaa",
          2816 => x"38ff5373",
          2817 => x"527551fd",
          2818 => x"a43f828c",
          2819 => x"dc085482",
          2820 => x"8cdc0880",
          2821 => x"f2389339",
          2822 => x"825480eb",
          2823 => x"39815480",
          2824 => x"e639828c",
          2825 => x"dc085480",
          2826 => x"de397452",
          2827 => x"7851fb84",
          2828 => x"3f828cdc",
          2829 => x"0858828c",
          2830 => x"dc08802e",
          2831 => x"80c73882",
          2832 => x"8cdc0881",
          2833 => x"2ed23882",
          2834 => x"8cdc08ff",
          2835 => x"2ecf3880",
          2836 => x"53745275",
          2837 => x"51fcd63f",
          2838 => x"828cdc08",
          2839 => x"c5389816",
          2840 => x"08fe1190",
          2841 => x"18085755",
          2842 => x"57747427",
          2843 => x"90388115",
          2844 => x"90170c84",
          2845 => x"16338107",
          2846 => x"54738417",
          2847 => x"34775576",
          2848 => x"7826ffa6",
          2849 => x"38805473",
          2850 => x"828cdc0c",
          2851 => x"8a3d0d04",
          2852 => x"f63d0d7c",
          2853 => x"7e710859",
          2854 => x"5b5b7995",
          2855 => x"388c1708",
          2856 => x"5877802e",
          2857 => x"88389817",
          2858 => x"087826b2",
          2859 => x"388158ae",
          2860 => x"3979527a",
          2861 => x"51f9fd3f",
          2862 => x"81557482",
          2863 => x"8cdc0827",
          2864 => x"82e03882",
          2865 => x"8cdc0855",
          2866 => x"828cdc08",
          2867 => x"ff2e82d2",
          2868 => x"38981708",
          2869 => x"828cdc08",
          2870 => x"2682c738",
          2871 => x"79589017",
          2872 => x"08705654",
          2873 => x"73802e82",
          2874 => x"b938777a",
          2875 => x"2e098106",
          2876 => x"80e23881",
          2877 => x"1a569817",
          2878 => x"08762683",
          2879 => x"38825675",
          2880 => x"527a51f9",
          2881 => x"af3f8059",
          2882 => x"828cdc08",
          2883 => x"812e0981",
          2884 => x"06863882",
          2885 => x"8cdc0859",
          2886 => x"828cdc08",
          2887 => x"09703070",
          2888 => x"72078025",
          2889 => x"707c0782",
          2890 => x"8cdc0854",
          2891 => x"51515555",
          2892 => x"7381ef38",
          2893 => x"828cdc08",
          2894 => x"802e9538",
          2895 => x"8c170854",
          2896 => x"81742790",
          2897 => x"38739818",
          2898 => x"08278938",
          2899 => x"73588539",
          2900 => x"7580db38",
          2901 => x"77568116",
          2902 => x"56981708",
          2903 => x"76268938",
          2904 => x"82567578",
          2905 => x"2681ac38",
          2906 => x"75527a51",
          2907 => x"f8c63f82",
          2908 => x"8cdc0880",
          2909 => x"2eb83880",
          2910 => x"59828cdc",
          2911 => x"08812e09",
          2912 => x"81068638",
          2913 => x"828cdc08",
          2914 => x"59828cdc",
          2915 => x"08097030",
          2916 => x"70720780",
          2917 => x"25707c07",
          2918 => x"51515555",
          2919 => x"7380f838",
          2920 => x"75782e09",
          2921 => x"8106ffae",
          2922 => x"38735580",
          2923 => x"f539ff53",
          2924 => x"75527651",
          2925 => x"f9f73f82",
          2926 => x"8cdc0882",
          2927 => x"8cdc0830",
          2928 => x"70828cdc",
          2929 => x"08078025",
          2930 => x"51555579",
          2931 => x"802e9438",
          2932 => x"73802e8f",
          2933 => x"38755379",
          2934 => x"527651f9",
          2935 => x"d03f828c",
          2936 => x"dc085574",
          2937 => x"a538758c",
          2938 => x"180c9817",
          2939 => x"08fe0590",
          2940 => x"18085654",
          2941 => x"74742686",
          2942 => x"38ff1590",
          2943 => x"180c8417",
          2944 => x"33810754",
          2945 => x"73841834",
          2946 => x"9739ff56",
          2947 => x"74812e90",
          2948 => x"388c3980",
          2949 => x"558c3982",
          2950 => x"8cdc0855",
          2951 => x"85398156",
          2952 => x"75557482",
          2953 => x"8cdc0c8c",
          2954 => x"3d0d04f8",
          2955 => x"3d0d7a70",
          2956 => x"5255f3f0",
          2957 => x"3f828cdc",
          2958 => x"08588156",
          2959 => x"828cdc08",
          2960 => x"80d8387b",
          2961 => x"527451f6",
          2962 => x"c13f828c",
          2963 => x"dc08828c",
          2964 => x"dc08b017",
          2965 => x"0c598480",
          2966 => x"537752b4",
          2967 => x"15705257",
          2968 => x"f2c83f77",
          2969 => x"56843981",
          2970 => x"16568a15",
          2971 => x"22587578",
          2972 => x"27973881",
          2973 => x"54751953",
          2974 => x"76528115",
          2975 => x"3351ede9",
          2976 => x"3f828cdc",
          2977 => x"08802edf",
          2978 => x"388a1522",
          2979 => x"76327030",
          2980 => x"70720770",
          2981 => x"9f2a5351",
          2982 => x"56567582",
          2983 => x"8cdc0c8a",
          2984 => x"3d0d04f8",
          2985 => x"3d0d7a7c",
          2986 => x"71085856",
          2987 => x"5774f080",
          2988 => x"0a2680f1",
          2989 => x"38749f06",
          2990 => x"537280e9",
          2991 => x"38749018",
          2992 => x"0c881708",
          2993 => x"5473aa38",
          2994 => x"75335382",
          2995 => x"73278838",
          2996 => x"a8160854",
          2997 => x"739b3874",
          2998 => x"852a5382",
          2999 => x"0b881722",
          3000 => x"5a587279",
          3001 => x"2780fe38",
          3002 => x"a8160898",
          3003 => x"180c80cd",
          3004 => x"398a1622",
          3005 => x"70892b54",
          3006 => x"58727526",
          3007 => x"b2387352",
          3008 => x"7651f5b0",
          3009 => x"3f828cdc",
          3010 => x"0854828c",
          3011 => x"dc08ff2e",
          3012 => x"bd38810b",
          3013 => x"828cdc08",
          3014 => x"278b3898",
          3015 => x"1608828c",
          3016 => x"dc082685",
          3017 => x"388258bd",
          3018 => x"39747331",
          3019 => x"55cb3973",
          3020 => x"527551f4",
          3021 => x"d53f828c",
          3022 => x"dc089818",
          3023 => x"0c739418",
          3024 => x"0c981708",
          3025 => x"53825872",
          3026 => x"802e9a38",
          3027 => x"85398158",
          3028 => x"94397489",
          3029 => x"2a139818",
          3030 => x"0c7483ff",
          3031 => x"0616b405",
          3032 => x"9c180c80",
          3033 => x"5877828c",
          3034 => x"dc0c8a3d",
          3035 => x"0d04f83d",
          3036 => x"0d7a7008",
          3037 => x"901208a0",
          3038 => x"05595754",
          3039 => x"f0800a77",
          3040 => x"27863880",
          3041 => x"0b98150c",
          3042 => x"98140853",
          3043 => x"84557280",
          3044 => x"2e81cb38",
          3045 => x"7683ff06",
          3046 => x"587781b5",
          3047 => x"38811398",
          3048 => x"150c9414",
          3049 => x"08557492",
          3050 => x"3876852a",
          3051 => x"88172256",
          3052 => x"53747326",
          3053 => x"819b3880",
          3054 => x"c0398a16",
          3055 => x"22ff0577",
          3056 => x"892a0653",
          3057 => x"72818a38",
          3058 => x"74527351",
          3059 => x"f3e63f82",
          3060 => x"8cdc0853",
          3061 => x"8255810b",
          3062 => x"828cdc08",
          3063 => x"2780ff38",
          3064 => x"8155828c",
          3065 => x"dc08ff2e",
          3066 => x"80f43898",
          3067 => x"1608828c",
          3068 => x"dc082680",
          3069 => x"ca387b8a",
          3070 => x"38779815",
          3071 => x"0c845580",
          3072 => x"dd399414",
          3073 => x"08527351",
          3074 => x"f9863f82",
          3075 => x"8cdc0853",
          3076 => x"8755828c",
          3077 => x"dc08802e",
          3078 => x"80c43882",
          3079 => x"55828cdc",
          3080 => x"08812eba",
          3081 => x"38815582",
          3082 => x"8cdc08ff",
          3083 => x"2eb03882",
          3084 => x"8cdc0852",
          3085 => x"7551fbf3",
          3086 => x"3f828cdc",
          3087 => x"08a03872",
          3088 => x"94150c72",
          3089 => x"527551f2",
          3090 => x"c13f828c",
          3091 => x"dc089815",
          3092 => x"0c769015",
          3093 => x"0c7716b4",
          3094 => x"059c150c",
          3095 => x"80557482",
          3096 => x"8cdc0c8a",
          3097 => x"3d0d04f7",
          3098 => x"3d0d7b7d",
          3099 => x"71085b5b",
          3100 => x"57805276",
          3101 => x"51fcac3f",
          3102 => x"828cdc08",
          3103 => x"54828cdc",
          3104 => x"0880ec38",
          3105 => x"828cdc08",
          3106 => x"56981708",
          3107 => x"527851f0",
          3108 => x"833f828c",
          3109 => x"dc085482",
          3110 => x"8cdc0880",
          3111 => x"d238828c",
          3112 => x"dc089c18",
          3113 => x"08703351",
          3114 => x"54587281",
          3115 => x"e52e0981",
          3116 => x"06833881",
          3117 => x"58828cdc",
          3118 => x"08557283",
          3119 => x"38815577",
          3120 => x"75075372",
          3121 => x"802e8e38",
          3122 => x"81165675",
          3123 => x"7a2e0981",
          3124 => x"068838a5",
          3125 => x"39828cdc",
          3126 => x"08568152",
          3127 => x"7651fd8e",
          3128 => x"3f828cdc",
          3129 => x"0854828c",
          3130 => x"dc08802e",
          3131 => x"ff9b3873",
          3132 => x"842e0981",
          3133 => x"06833887",
          3134 => x"5473828c",
          3135 => x"dc0c8b3d",
          3136 => x"0d04fd3d",
          3137 => x"0d769a11",
          3138 => x"5254ebec",
          3139 => x"3f828cdc",
          3140 => x"0883ffff",
          3141 => x"06767033",
          3142 => x"51535371",
          3143 => x"832e0981",
          3144 => x"06903894",
          3145 => x"1451ebd0",
          3146 => x"3f828cdc",
          3147 => x"08902b73",
          3148 => x"07537282",
          3149 => x"8cdc0c85",
          3150 => x"3d0d04fc",
          3151 => x"3d0d7779",
          3152 => x"7083ffff",
          3153 => x"06549a12",
          3154 => x"535555eb",
          3155 => x"ed3f7670",
          3156 => x"33515372",
          3157 => x"832e0981",
          3158 => x"068b3873",
          3159 => x"902a5294",
          3160 => x"1551ebd6",
          3161 => x"3f863d0d",
          3162 => x"04f73d0d",
          3163 => x"7b7d5b55",
          3164 => x"8475085a",
          3165 => x"58981508",
          3166 => x"802e818a",
          3167 => x"38981508",
          3168 => x"527851ee",
          3169 => x"8f3f828c",
          3170 => x"dc085882",
          3171 => x"8cdc0880",
          3172 => x"f5389c15",
          3173 => x"08703355",
          3174 => x"53738638",
          3175 => x"845880e6",
          3176 => x"398b1333",
          3177 => x"70bf0670",
          3178 => x"81ff0658",
          3179 => x"51537286",
          3180 => x"1634828c",
          3181 => x"dc085373",
          3182 => x"81e52e83",
          3183 => x"38815373",
          3184 => x"ae2ea938",
          3185 => x"81707406",
          3186 => x"54577280",
          3187 => x"2e9e3875",
          3188 => x"8f2e9938",
          3189 => x"828cdc08",
          3190 => x"76df0654",
          3191 => x"5472882e",
          3192 => x"09810683",
          3193 => x"38765473",
          3194 => x"7a2ea038",
          3195 => x"80527451",
          3196 => x"fafc3f82",
          3197 => x"8cdc0858",
          3198 => x"828cdc08",
          3199 => x"89389815",
          3200 => x"08fefa38",
          3201 => x"8639800b",
          3202 => x"98160c77",
          3203 => x"828cdc0c",
          3204 => x"8b3d0d04",
          3205 => x"fb3d0d77",
          3206 => x"70085754",
          3207 => x"81527351",
          3208 => x"fcc53f82",
          3209 => x"8cdc0855",
          3210 => x"828cdc08",
          3211 => x"b4389814",
          3212 => x"08527551",
          3213 => x"ecde3f82",
          3214 => x"8cdc0855",
          3215 => x"828cdc08",
          3216 => x"a038a053",
          3217 => x"828cdc08",
          3218 => x"529c1408",
          3219 => x"51eadb3f",
          3220 => x"8b53a014",
          3221 => x"529c1408",
          3222 => x"51eaac3f",
          3223 => x"810b8317",
          3224 => x"3474828c",
          3225 => x"dc0c873d",
          3226 => x"0d04fd3d",
          3227 => x"0d757008",
          3228 => x"98120854",
          3229 => x"70535553",
          3230 => x"ec9a3f82",
          3231 => x"8cdc088d",
          3232 => x"389c1308",
          3233 => x"53e57334",
          3234 => x"810b8315",
          3235 => x"34853d0d",
          3236 => x"04fa3d0d",
          3237 => x"787a5757",
          3238 => x"800b8917",
          3239 => x"34981708",
          3240 => x"802e8182",
          3241 => x"38807089",
          3242 => x"18555555",
          3243 => x"9c170814",
          3244 => x"70338116",
          3245 => x"56515271",
          3246 => x"a02ea838",
          3247 => x"71852e09",
          3248 => x"81068438",
          3249 => x"81e55273",
          3250 => x"892e0981",
          3251 => x"068b38ae",
          3252 => x"73708105",
          3253 => x"55348115",
          3254 => x"55717370",
          3255 => x"81055534",
          3256 => x"8115558a",
          3257 => x"7427c538",
          3258 => x"75158805",
          3259 => x"52800b81",
          3260 => x"13349c17",
          3261 => x"08528b12",
          3262 => x"33881734",
          3263 => x"9c17089c",
          3264 => x"115252e8",
          3265 => x"8a3f828c",
          3266 => x"dc08760c",
          3267 => x"961251e7",
          3268 => x"e73f828c",
          3269 => x"dc088617",
          3270 => x"23981251",
          3271 => x"e7da3f82",
          3272 => x"8cdc0884",
          3273 => x"1723883d",
          3274 => x"0d04f33d",
          3275 => x"0d7f7008",
          3276 => x"5e5b8061",
          3277 => x"70335155",
          3278 => x"5573af2e",
          3279 => x"83388155",
          3280 => x"7380dc2e",
          3281 => x"91387480",
          3282 => x"2e8c3894",
          3283 => x"1d08881c",
          3284 => x"0caa3981",
          3285 => x"15418061",
          3286 => x"70335656",
          3287 => x"5673af2e",
          3288 => x"09810683",
          3289 => x"38815673",
          3290 => x"80dc3270",
          3291 => x"30708025",
          3292 => x"78075151",
          3293 => x"5473dc38",
          3294 => x"73881c0c",
          3295 => x"60703351",
          3296 => x"54739f26",
          3297 => x"9638ff80",
          3298 => x"0bab1c34",
          3299 => x"80527a51",
          3300 => x"f6913f82",
          3301 => x"8cdc0855",
          3302 => x"85983991",
          3303 => x"3d61a01d",
          3304 => x"5c5a5e8b",
          3305 => x"53a05279",
          3306 => x"51e7ff3f",
          3307 => x"80705957",
          3308 => x"88793355",
          3309 => x"5c73ae2e",
          3310 => x"09810680",
          3311 => x"d4387818",
          3312 => x"7033811a",
          3313 => x"71ae3270",
          3314 => x"30709f2a",
          3315 => x"73822607",
          3316 => x"5151535a",
          3317 => x"5754738c",
          3318 => x"38791754",
          3319 => x"75743481",
          3320 => x"1757db39",
          3321 => x"75af3270",
          3322 => x"30709f2a",
          3323 => x"51515475",
          3324 => x"80dc2e8c",
          3325 => x"3873802e",
          3326 => x"873875a0",
          3327 => x"2682bd38",
          3328 => x"77197e0c",
          3329 => x"a454a076",
          3330 => x"2782bd38",
          3331 => x"a05482b8",
          3332 => x"39781870",
          3333 => x"33811a5a",
          3334 => x"5754a076",
          3335 => x"2781fc38",
          3336 => x"75af3270",
          3337 => x"307780dc",
          3338 => x"32703072",
          3339 => x"80257180",
          3340 => x"25075151",
          3341 => x"56515573",
          3342 => x"802eac38",
          3343 => x"84398118",
          3344 => x"5880781a",
          3345 => x"70335155",
          3346 => x"5573af2e",
          3347 => x"09810683",
          3348 => x"38815573",
          3349 => x"80dc3270",
          3350 => x"30708025",
          3351 => x"77075151",
          3352 => x"5473db38",
          3353 => x"81b53975",
          3354 => x"ae2e0981",
          3355 => x"06833881",
          3356 => x"54767c27",
          3357 => x"74075473",
          3358 => x"802ea238",
          3359 => x"7b8b3270",
          3360 => x"3077ae32",
          3361 => x"70307280",
          3362 => x"25719f2a",
          3363 => x"07535156",
          3364 => x"51557481",
          3365 => x"a7388857",
          3366 => x"8b5cfef5",
          3367 => x"3975982b",
          3368 => x"54738025",
          3369 => x"8c387580",
          3370 => x"ff0681fa",
          3371 => x"ec113357",
          3372 => x"547551e6",
          3373 => x"e13f828c",
          3374 => x"dc08802e",
          3375 => x"b2387818",
          3376 => x"7033811a",
          3377 => x"71545a56",
          3378 => x"54e6d23f",
          3379 => x"828cdc08",
          3380 => x"802e80e8",
          3381 => x"38ff1c54",
          3382 => x"76742780",
          3383 => x"df387917",
          3384 => x"54757434",
          3385 => x"81177a11",
          3386 => x"55577474",
          3387 => x"34a73975",
          3388 => x"5281fa8c",
          3389 => x"51e5fe3f",
          3390 => x"828cdc08",
          3391 => x"bf38ff9f",
          3392 => x"16547399",
          3393 => x"268938e0",
          3394 => x"167081ff",
          3395 => x"06575479",
          3396 => x"17547574",
          3397 => x"34811757",
          3398 => x"fdf73977",
          3399 => x"197e0c76",
          3400 => x"802e9938",
          3401 => x"79335473",
          3402 => x"81e52e09",
          3403 => x"81068438",
          3404 => x"857a3484",
          3405 => x"54a07627",
          3406 => x"8f388b39",
          3407 => x"865581f2",
          3408 => x"39845680",
          3409 => x"f3398054",
          3410 => x"738b1b34",
          3411 => x"807b0858",
          3412 => x"527a51f2",
          3413 => x"ce3f828c",
          3414 => x"dc085682",
          3415 => x"8cdc0880",
          3416 => x"d738981b",
          3417 => x"08527651",
          3418 => x"e6aa3f82",
          3419 => x"8cdc0856",
          3420 => x"828cdc08",
          3421 => x"80c2389c",
          3422 => x"1b087033",
          3423 => x"55557380",
          3424 => x"2effbe38",
          3425 => x"8b1533bf",
          3426 => x"06547386",
          3427 => x"1c348b15",
          3428 => x"3370832a",
          3429 => x"70810651",
          3430 => x"55587392",
          3431 => x"388b5379",
          3432 => x"527451e4",
          3433 => x"9f3f828c",
          3434 => x"dc08802e",
          3435 => x"8b387552",
          3436 => x"7a51f3ba",
          3437 => x"3fff9f39",
          3438 => x"75ab1c33",
          3439 => x"57557480",
          3440 => x"2ebb3874",
          3441 => x"842e0981",
          3442 => x"0680e738",
          3443 => x"75852a70",
          3444 => x"81067782",
          3445 => x"2a585154",
          3446 => x"73802e96",
          3447 => x"38758106",
          3448 => x"5473802e",
          3449 => x"fbb538ff",
          3450 => x"800bab1c",
          3451 => x"34805580",
          3452 => x"c1397581",
          3453 => x"065473ba",
          3454 => x"388555b6",
          3455 => x"3975822a",
          3456 => x"70810651",
          3457 => x"5473ab38",
          3458 => x"861b3370",
          3459 => x"842a7081",
          3460 => x"06515555",
          3461 => x"73802ee1",
          3462 => x"38901b08",
          3463 => x"83ff061d",
          3464 => x"b405527c",
          3465 => x"51f5db3f",
          3466 => x"828cdc08",
          3467 => x"881c0cfa",
          3468 => x"ea397482",
          3469 => x"8cdc0c8f",
          3470 => x"3d0d04f6",
          3471 => x"3d0d7c5b",
          3472 => x"ff7b0870",
          3473 => x"71735559",
          3474 => x"5c555973",
          3475 => x"802e81c6",
          3476 => x"38757081",
          3477 => x"05573370",
          3478 => x"a0265252",
          3479 => x"71ba2e8d",
          3480 => x"3870ee38",
          3481 => x"71ba2e09",
          3482 => x"810681a5",
          3483 => x"387333d0",
          3484 => x"117081ff",
          3485 => x"06515253",
          3486 => x"70892691",
          3487 => x"38821473",
          3488 => x"81ff06d0",
          3489 => x"05565271",
          3490 => x"762e80f7",
          3491 => x"38800b81",
          3492 => x"fadc5955",
          3493 => x"77087a55",
          3494 => x"57767081",
          3495 => x"05583374",
          3496 => x"70810556",
          3497 => x"33ff9f12",
          3498 => x"53535370",
          3499 => x"99268938",
          3500 => x"e0137081",
          3501 => x"ff065451",
          3502 => x"ff9f1251",
          3503 => x"70992689",
          3504 => x"38e01270",
          3505 => x"81ff0653",
          3506 => x"51723070",
          3507 => x"9f2a5151",
          3508 => x"72722e09",
          3509 => x"81068538",
          3510 => x"70ffbe38",
          3511 => x"72307477",
          3512 => x"32703070",
          3513 => x"72079f2a",
          3514 => x"739f2a07",
          3515 => x"53545451",
          3516 => x"70802e8f",
          3517 => x"38811584",
          3518 => x"19595583",
          3519 => x"7525ff94",
          3520 => x"388b3974",
          3521 => x"83248638",
          3522 => x"74767c0c",
          3523 => x"59785186",
          3524 => x"39828da0",
          3525 => x"33517082",
          3526 => x"8cdc0c8c",
          3527 => x"3d0d04fa",
          3528 => x"3d0d7856",
          3529 => x"800b8317",
          3530 => x"34ff0bb0",
          3531 => x"170c7952",
          3532 => x"7551e2e0",
          3533 => x"3f845582",
          3534 => x"8cdc0881",
          3535 => x"803884b2",
          3536 => x"1651dfb4",
          3537 => x"3f828cdc",
          3538 => x"0883ffff",
          3539 => x"06548355",
          3540 => x"7382d4d5",
          3541 => x"2e098106",
          3542 => x"80e33880",
          3543 => x"0bb41733",
          3544 => x"56577481",
          3545 => x"e92e0981",
          3546 => x"06833881",
          3547 => x"577481eb",
          3548 => x"32703070",
          3549 => x"80257907",
          3550 => x"51515473",
          3551 => x"8a387481",
          3552 => x"e82e0981",
          3553 => x"06b53883",
          3554 => x"5381fa9c",
          3555 => x"5280ea16",
          3556 => x"51e0b13f",
          3557 => x"828cdc08",
          3558 => x"55828cdc",
          3559 => x"08802e9d",
          3560 => x"38855381",
          3561 => x"faa05281",
          3562 => x"861651e0",
          3563 => x"973f828c",
          3564 => x"dc085582",
          3565 => x"8cdc0880",
          3566 => x"2e833882",
          3567 => x"5574828c",
          3568 => x"dc0c883d",
          3569 => x"0d04f23d",
          3570 => x"0d610284",
          3571 => x"0580cb05",
          3572 => x"33585580",
          3573 => x"750c6051",
          3574 => x"fce13f82",
          3575 => x"8cdc0858",
          3576 => x"8b56800b",
          3577 => x"828cdc08",
          3578 => x"2486fc38",
          3579 => x"828cdc08",
          3580 => x"8429828d",
          3581 => x"8c057008",
          3582 => x"55538c56",
          3583 => x"73802e86",
          3584 => x"e6387375",
          3585 => x"0c7681fe",
          3586 => x"06743354",
          3587 => x"5772802e",
          3588 => x"ae388114",
          3589 => x"3351d7ca",
          3590 => x"3f828cdc",
          3591 => x"0881ff06",
          3592 => x"70810654",
          3593 => x"55729838",
          3594 => x"76802e86",
          3595 => x"b8387482",
          3596 => x"2a708106",
          3597 => x"51538a56",
          3598 => x"7286ac38",
          3599 => x"86a73980",
          3600 => x"74347781",
          3601 => x"15348152",
          3602 => x"81143351",
          3603 => x"d7b23f82",
          3604 => x"8cdc0881",
          3605 => x"ff067081",
          3606 => x"06545583",
          3607 => x"56728687",
          3608 => x"3876802e",
          3609 => x"8f387482",
          3610 => x"2a708106",
          3611 => x"51538a56",
          3612 => x"7285f438",
          3613 => x"80705374",
          3614 => x"525bfda3",
          3615 => x"3f828cdc",
          3616 => x"0881ff06",
          3617 => x"5776822e",
          3618 => x"09810680",
          3619 => x"e2388c3d",
          3620 => x"74565883",
          3621 => x"5683f615",
          3622 => x"33705853",
          3623 => x"72802e8d",
          3624 => x"3883fa15",
          3625 => x"51dce83f",
          3626 => x"828cdc08",
          3627 => x"57767870",
          3628 => x"84055a0c",
          3629 => x"ff169016",
          3630 => x"56567580",
          3631 => x"25d73880",
          3632 => x"0b8d3d54",
          3633 => x"56727084",
          3634 => x"0554085b",
          3635 => x"83577a80",
          3636 => x"2e95387a",
          3637 => x"527351fc",
          3638 => x"c63f828c",
          3639 => x"dc0881ff",
          3640 => x"06578177",
          3641 => x"27893881",
          3642 => x"16568376",
          3643 => x"27d73881",
          3644 => x"5676842e",
          3645 => x"84f1388d",
          3646 => x"56768126",
          3647 => x"84e938bf",
          3648 => x"1451dbf4",
          3649 => x"3f828cdc",
          3650 => x"0883ffff",
          3651 => x"06537284",
          3652 => x"802e0981",
          3653 => x"0684d038",
          3654 => x"80ca1451",
          3655 => x"dbda3f82",
          3656 => x"8cdc0883",
          3657 => x"ffff0658",
          3658 => x"778d3880",
          3659 => x"d81451db",
          3660 => x"de3f828c",
          3661 => x"dc085877",
          3662 => x"9c150c80",
          3663 => x"c4143382",
          3664 => x"153480c4",
          3665 => x"1433ff11",
          3666 => x"7081ff06",
          3667 => x"5154558d",
          3668 => x"56728126",
          3669 => x"84913874",
          3670 => x"81ff0678",
          3671 => x"712980c1",
          3672 => x"16335259",
          3673 => x"53728a15",
          3674 => x"2372802e",
          3675 => x"8b38ff13",
          3676 => x"73065372",
          3677 => x"802e8638",
          3678 => x"8d5683eb",
          3679 => x"3980c514",
          3680 => x"51daf53f",
          3681 => x"828cdc08",
          3682 => x"53828cdc",
          3683 => x"08881523",
          3684 => x"728f0657",
          3685 => x"8d567683",
          3686 => x"ce3880c7",
          3687 => x"1451dad8",
          3688 => x"3f828cdc",
          3689 => x"0883ffff",
          3690 => x"0655748d",
          3691 => x"3880d414",
          3692 => x"51dadc3f",
          3693 => x"828cdc08",
          3694 => x"5580c214",
          3695 => x"51dab93f",
          3696 => x"828cdc08",
          3697 => x"83ffff06",
          3698 => x"538d5672",
          3699 => x"802e8397",
          3700 => x"38881422",
          3701 => x"78147184",
          3702 => x"2a055a5a",
          3703 => x"78752683",
          3704 => x"86388a14",
          3705 => x"22527479",
          3706 => x"3151ff96",
          3707 => x"ee3f828c",
          3708 => x"dc085582",
          3709 => x"8cdc0880",
          3710 => x"2e82ec38",
          3711 => x"828cdc08",
          3712 => x"80ffffff",
          3713 => x"f5268338",
          3714 => x"83577483",
          3715 => x"fff52683",
          3716 => x"38825774",
          3717 => x"9ff52685",
          3718 => x"38815789",
          3719 => x"398d5676",
          3720 => x"802e82c3",
          3721 => x"38821570",
          3722 => x"98160c7b",
          3723 => x"a0160c73",
          3724 => x"1c70a417",
          3725 => x"0c7a1dac",
          3726 => x"170c5455",
          3727 => x"76832e09",
          3728 => x"8106af38",
          3729 => x"80de1451",
          3730 => x"d9ae3f82",
          3731 => x"8cdc0883",
          3732 => x"ffff0653",
          3733 => x"8d567282",
          3734 => x"8e387982",
          3735 => x"8a3880e0",
          3736 => x"1451d9ab",
          3737 => x"3f828cdc",
          3738 => x"08a8150c",
          3739 => x"74822b53",
          3740 => x"a2398d56",
          3741 => x"79802e81",
          3742 => x"ee387713",
          3743 => x"a8150c74",
          3744 => x"15537682",
          3745 => x"2e8d3874",
          3746 => x"10157081",
          3747 => x"2a768106",
          3748 => x"05515383",
          3749 => x"ff13892a",
          3750 => x"538d5672",
          3751 => x"9c150826",
          3752 => x"81c538ff",
          3753 => x"0b90150c",
          3754 => x"ff0b8c15",
          3755 => x"0cff800b",
          3756 => x"84153476",
          3757 => x"832e0981",
          3758 => x"06819238",
          3759 => x"80e41451",
          3760 => x"d8b63f82",
          3761 => x"8cdc0883",
          3762 => x"ffff0653",
          3763 => x"72812e09",
          3764 => x"810680f9",
          3765 => x"38811b52",
          3766 => x"7351dbb8",
          3767 => x"3f828cdc",
          3768 => x"0880ea38",
          3769 => x"828cdc08",
          3770 => x"84153484",
          3771 => x"b21451d8",
          3772 => x"873f828c",
          3773 => x"dc0883ff",
          3774 => x"ff065372",
          3775 => x"82d4d52e",
          3776 => x"09810680",
          3777 => x"c838b414",
          3778 => x"51d8843f",
          3779 => x"828cdc08",
          3780 => x"848b85a4",
          3781 => x"d22e0981",
          3782 => x"06b33884",
          3783 => x"981451d7",
          3784 => x"ee3f828c",
          3785 => x"dc08868a",
          3786 => x"85e4f22e",
          3787 => x"0981069d",
          3788 => x"38849c14",
          3789 => x"51d7d83f",
          3790 => x"828cdc08",
          3791 => x"90150c84",
          3792 => x"a01451d7",
          3793 => x"ca3f828c",
          3794 => x"dc088c15",
          3795 => x"0c767434",
          3796 => x"828d9c22",
          3797 => x"81055372",
          3798 => x"828d9c23",
          3799 => x"72861523",
          3800 => x"800b9415",
          3801 => x"0c805675",
          3802 => x"828cdc0c",
          3803 => x"903d0d04",
          3804 => x"fb3d0d77",
          3805 => x"54895573",
          3806 => x"802eb938",
          3807 => x"73085372",
          3808 => x"802eb138",
          3809 => x"72335271",
          3810 => x"802ea938",
          3811 => x"86132284",
          3812 => x"15225752",
          3813 => x"71762e09",
          3814 => x"81069938",
          3815 => x"81133351",
          3816 => x"d0c03f82",
          3817 => x"8cdc0881",
          3818 => x"06527188",
          3819 => x"38717408",
          3820 => x"54558339",
          3821 => x"80537873",
          3822 => x"710c5274",
          3823 => x"828cdc0c",
          3824 => x"873d0d04",
          3825 => x"fa3d0d02",
          3826 => x"ab05337a",
          3827 => x"58893dfc",
          3828 => x"055256f4",
          3829 => x"e63f8b54",
          3830 => x"800b828c",
          3831 => x"dc0824bc",
          3832 => x"38828cdc",
          3833 => x"08842982",
          3834 => x"8d8c0570",
          3835 => x"08555573",
          3836 => x"802e8438",
          3837 => x"80743478",
          3838 => x"5473802e",
          3839 => x"84388074",
          3840 => x"3478750c",
          3841 => x"75547580",
          3842 => x"2e923880",
          3843 => x"53893d70",
          3844 => x"53840551",
          3845 => x"f7b03f82",
          3846 => x"8cdc0854",
          3847 => x"73828cdc",
          3848 => x"0c883d0d",
          3849 => x"04eb3d0d",
          3850 => x"67028405",
          3851 => x"80e70533",
          3852 => x"59598954",
          3853 => x"78802e84",
          3854 => x"c83877bf",
          3855 => x"06705498",
          3856 => x"3dd00553",
          3857 => x"993d8405",
          3858 => x"5258f6fa",
          3859 => x"3f828cdc",
          3860 => x"0855828c",
          3861 => x"dc0884a4",
          3862 => x"387a5c68",
          3863 => x"528c3d70",
          3864 => x"5256edc6",
          3865 => x"3f828cdc",
          3866 => x"0855828c",
          3867 => x"dc089238",
          3868 => x"0280d705",
          3869 => x"3370982b",
          3870 => x"55577380",
          3871 => x"25833886",
          3872 => x"55779c06",
          3873 => x"5473802e",
          3874 => x"81ab3874",
          3875 => x"802e9538",
          3876 => x"74842e09",
          3877 => x"8106aa38",
          3878 => x"7551eaf8",
          3879 => x"3f828cdc",
          3880 => x"08559e39",
          3881 => x"02b20533",
          3882 => x"91065473",
          3883 => x"81b83877",
          3884 => x"822a7081",
          3885 => x"06515473",
          3886 => x"802e8e38",
          3887 => x"885583bc",
          3888 => x"39778807",
          3889 => x"587483b4",
          3890 => x"3877832a",
          3891 => x"70810651",
          3892 => x"5473802e",
          3893 => x"81af3862",
          3894 => x"527a51e8",
          3895 => x"a53f828c",
          3896 => x"dc085682",
          3897 => x"88b20a52",
          3898 => x"628e0551",
          3899 => x"d4ea3f62",
          3900 => x"54a00b8b",
          3901 => x"15348053",
          3902 => x"62527a51",
          3903 => x"e8bd3f80",
          3904 => x"52629c05",
          3905 => x"51d4d13f",
          3906 => x"7a54810b",
          3907 => x"83153475",
          3908 => x"802e80f1",
          3909 => x"387ab011",
          3910 => x"08515480",
          3911 => x"53755297",
          3912 => x"3dd40551",
          3913 => x"ddbe3f82",
          3914 => x"8cdc0855",
          3915 => x"828cdc08",
          3916 => x"82ca38b7",
          3917 => x"397482c4",
          3918 => x"3802b205",
          3919 => x"3370842a",
          3920 => x"70810651",
          3921 => x"55567380",
          3922 => x"2e863884",
          3923 => x"5582ad39",
          3924 => x"77812a70",
          3925 => x"81065154",
          3926 => x"73802ea9",
          3927 => x"38758106",
          3928 => x"5473802e",
          3929 => x"a0388755",
          3930 => x"82923973",
          3931 => x"527a51d6",
          3932 => x"a33f828c",
          3933 => x"dc087bff",
          3934 => x"188c120c",
          3935 => x"5555828c",
          3936 => x"dc0881f8",
          3937 => x"3877832a",
          3938 => x"70810651",
          3939 => x"5473802e",
          3940 => x"86387780",
          3941 => x"c007587a",
          3942 => x"b01108a0",
          3943 => x"1b0c63a4",
          3944 => x"1b0c6353",
          3945 => x"705257e6",
          3946 => x"d93f828c",
          3947 => x"dc08828c",
          3948 => x"dc08881b",
          3949 => x"0c639c05",
          3950 => x"525ad2d3",
          3951 => x"3f828cdc",
          3952 => x"08828cdc",
          3953 => x"088c1b0c",
          3954 => x"777a0c56",
          3955 => x"86172284",
          3956 => x"1a237790",
          3957 => x"1a34800b",
          3958 => x"911a3480",
          3959 => x"0b9c1a0c",
          3960 => x"800b941a",
          3961 => x"0c77852a",
          3962 => x"70810651",
          3963 => x"5473802e",
          3964 => x"818d3882",
          3965 => x"8cdc0880",
          3966 => x"2e818438",
          3967 => x"828cdc08",
          3968 => x"941a0c8a",
          3969 => x"17227089",
          3970 => x"2b7b5259",
          3971 => x"57a83976",
          3972 => x"527851d7",
          3973 => x"9f3f828c",
          3974 => x"dc085782",
          3975 => x"8cdc0881",
          3976 => x"26833882",
          3977 => x"55828cdc",
          3978 => x"08ff2e09",
          3979 => x"81068338",
          3980 => x"79557578",
          3981 => x"31567430",
          3982 => x"70760780",
          3983 => x"25515477",
          3984 => x"76278a38",
          3985 => x"81707506",
          3986 => x"555a73c3",
          3987 => x"3876981a",
          3988 => x"0c74a938",
          3989 => x"7583ff06",
          3990 => x"5473802e",
          3991 => x"a2387652",
          3992 => x"7a51d6a6",
          3993 => x"3f828cdc",
          3994 => x"08853882",
          3995 => x"558e3975",
          3996 => x"892a828c",
          3997 => x"dc08059c",
          3998 => x"1a0c8439",
          3999 => x"80790c74",
          4000 => x"5473828c",
          4001 => x"dc0c973d",
          4002 => x"0d04f23d",
          4003 => x"0d606365",
          4004 => x"6440405d",
          4005 => x"59807e0c",
          4006 => x"903dfc05",
          4007 => x"527851f9",
          4008 => x"cf3f828c",
          4009 => x"dc085582",
          4010 => x"8cdc088a",
          4011 => x"38911933",
          4012 => x"5574802e",
          4013 => x"86387456",
          4014 => x"82c43990",
          4015 => x"19338106",
          4016 => x"55875674",
          4017 => x"802e82b6",
          4018 => x"38953982",
          4019 => x"0b911a34",
          4020 => x"825682aa",
          4021 => x"39810b91",
          4022 => x"1a348156",
          4023 => x"82a0398c",
          4024 => x"1908941a",
          4025 => x"08315574",
          4026 => x"7c278338",
          4027 => x"745c7b80",
          4028 => x"2e828938",
          4029 => x"94190870",
          4030 => x"83ff0656",
          4031 => x"567481b2",
          4032 => x"387e8a11",
          4033 => x"22ff0577",
          4034 => x"892a065b",
          4035 => x"5579a838",
          4036 => x"75873888",
          4037 => x"1908558f",
          4038 => x"39981908",
          4039 => x"527851d5",
          4040 => x"933f828c",
          4041 => x"dc085581",
          4042 => x"7527ff9f",
          4043 => x"3874ff2e",
          4044 => x"ffa33874",
          4045 => x"981a0c98",
          4046 => x"1908527e",
          4047 => x"51d4cb3f",
          4048 => x"828cdc08",
          4049 => x"802eff83",
          4050 => x"38828cdc",
          4051 => x"081a7c89",
          4052 => x"2a595777",
          4053 => x"802e80d6",
          4054 => x"38771a7f",
          4055 => x"8a112258",
          4056 => x"5c557575",
          4057 => x"27853875",
          4058 => x"7a315877",
          4059 => x"5476537c",
          4060 => x"52811b33",
          4061 => x"51ca883f",
          4062 => x"828cdc08",
          4063 => x"fed7387e",
          4064 => x"83113356",
          4065 => x"5674802e",
          4066 => x"9f38b016",
          4067 => x"08773155",
          4068 => x"74782794",
          4069 => x"38848053",
          4070 => x"b41652b0",
          4071 => x"16087731",
          4072 => x"892b7d05",
          4073 => x"51cfe03f",
          4074 => x"77892b56",
          4075 => x"b939769c",
          4076 => x"1a0c9419",
          4077 => x"0883ff06",
          4078 => x"84807131",
          4079 => x"57557b76",
          4080 => x"2783387b",
          4081 => x"569c1908",
          4082 => x"527e51d1",
          4083 => x"c73f828c",
          4084 => x"dc08fe81",
          4085 => x"38755394",
          4086 => x"190883ff",
          4087 => x"061fb405",
          4088 => x"527c51cf",
          4089 => x"a23f7b76",
          4090 => x"317e0817",
          4091 => x"7f0c761e",
          4092 => x"941b0818",
          4093 => x"941c0c5e",
          4094 => x"5cfdf339",
          4095 => x"80567582",
          4096 => x"8cdc0c90",
          4097 => x"3d0d04f2",
          4098 => x"3d0d6063",
          4099 => x"65644040",
          4100 => x"5d58807e",
          4101 => x"0c903dfc",
          4102 => x"05527751",
          4103 => x"f6d23f82",
          4104 => x"8cdc0855",
          4105 => x"828cdc08",
          4106 => x"8a389118",
          4107 => x"33557480",
          4108 => x"2e863874",
          4109 => x"5683b839",
          4110 => x"90183370",
          4111 => x"812a7081",
          4112 => x"06515656",
          4113 => x"87567480",
          4114 => x"2e83a438",
          4115 => x"9539820b",
          4116 => x"91193482",
          4117 => x"56839839",
          4118 => x"810b9119",
          4119 => x"34815683",
          4120 => x"8e399418",
          4121 => x"087c1156",
          4122 => x"56747627",
          4123 => x"84387509",
          4124 => x"5c7b802e",
          4125 => x"82ec3894",
          4126 => x"18087083",
          4127 => x"ff065656",
          4128 => x"7481fd38",
          4129 => x"7e8a1122",
          4130 => x"ff057789",
          4131 => x"2a065c55",
          4132 => x"7abf3875",
          4133 => x"8c388818",
          4134 => x"0855749c",
          4135 => x"387a5285",
          4136 => x"39981808",
          4137 => x"527751d7",
          4138 => x"e73f828c",
          4139 => x"dc085582",
          4140 => x"8cdc0880",
          4141 => x"2e82ab38",
          4142 => x"74812eff",
          4143 => x"913874ff",
          4144 => x"2eff9538",
          4145 => x"7498190c",
          4146 => x"88180885",
          4147 => x"38748819",
          4148 => x"0c7e55b0",
          4149 => x"15089c19",
          4150 => x"082e0981",
          4151 => x"068d3874",
          4152 => x"51cec13f",
          4153 => x"828cdc08",
          4154 => x"feee3898",
          4155 => x"1808527e",
          4156 => x"51d1973f",
          4157 => x"828cdc08",
          4158 => x"802efed2",
          4159 => x"38828cdc",
          4160 => x"081b7c89",
          4161 => x"2a5a5778",
          4162 => x"802e80d5",
          4163 => x"38781b7f",
          4164 => x"8a112258",
          4165 => x"5b557575",
          4166 => x"27853875",
          4167 => x"7b315978",
          4168 => x"5476537c",
          4169 => x"52811a33",
          4170 => x"51c8be3f",
          4171 => x"828cdc08",
          4172 => x"fea6387e",
          4173 => x"b0110878",
          4174 => x"31565674",
          4175 => x"79279b38",
          4176 => x"848053b0",
          4177 => x"16087731",
          4178 => x"892b7d05",
          4179 => x"52b41651",
          4180 => x"ccb53f7e",
          4181 => x"55800b83",
          4182 => x"16347889",
          4183 => x"2b5680db",
          4184 => x"398c1808",
          4185 => x"94190826",
          4186 => x"93387e51",
          4187 => x"cdb63f82",
          4188 => x"8cdc08fd",
          4189 => x"e3387e77",
          4190 => x"b0120c55",
          4191 => x"769c190c",
          4192 => x"94180883",
          4193 => x"ff068480",
          4194 => x"71315755",
          4195 => x"7b762783",
          4196 => x"387b569c",
          4197 => x"1808527e",
          4198 => x"51cdf93f",
          4199 => x"828cdc08",
          4200 => x"fdb63875",
          4201 => x"537c5294",
          4202 => x"180883ff",
          4203 => x"061fb405",
          4204 => x"51cbd43f",
          4205 => x"7e55810b",
          4206 => x"8316347b",
          4207 => x"76317e08",
          4208 => x"177f0c76",
          4209 => x"1e941a08",
          4210 => x"1870941c",
          4211 => x"0c8c1b08",
          4212 => x"58585e5c",
          4213 => x"74762783",
          4214 => x"38755574",
          4215 => x"8c190cfd",
          4216 => x"90399018",
          4217 => x"3380c007",
          4218 => x"55749019",
          4219 => x"34805675",
          4220 => x"828cdc0c",
          4221 => x"903d0d04",
          4222 => x"f83d0d7a",
          4223 => x"8b3dfc05",
          4224 => x"53705256",
          4225 => x"f2ea3f82",
          4226 => x"8cdc0857",
          4227 => x"828cdc08",
          4228 => x"80fb3890",
          4229 => x"16337086",
          4230 => x"2a708106",
          4231 => x"51555573",
          4232 => x"802e80e9",
          4233 => x"38a01608",
          4234 => x"527851cc",
          4235 => x"e73f828c",
          4236 => x"dc085782",
          4237 => x"8cdc0880",
          4238 => x"d438a416",
          4239 => x"088b1133",
          4240 => x"a0075555",
          4241 => x"738b1634",
          4242 => x"88160853",
          4243 => x"74527508",
          4244 => x"51dde83f",
          4245 => x"8c160852",
          4246 => x"9c1551c9",
          4247 => x"fb3f8288",
          4248 => x"b20a5296",
          4249 => x"1551c9f0",
          4250 => x"3f765292",
          4251 => x"1551c9ca",
          4252 => x"3f785481",
          4253 => x"0b831534",
          4254 => x"7851ccdf",
          4255 => x"3f828cdc",
          4256 => x"08901733",
          4257 => x"81bf0655",
          4258 => x"57739017",
          4259 => x"3476828c",
          4260 => x"dc0c8a3d",
          4261 => x"0d04fc3d",
          4262 => x"0d767052",
          4263 => x"54fed93f",
          4264 => x"828cdc08",
          4265 => x"53828cdc",
          4266 => x"089c3886",
          4267 => x"3dfc0552",
          4268 => x"7351f1bc",
          4269 => x"3f828cdc",
          4270 => x"0853828c",
          4271 => x"dc088738",
          4272 => x"828cdc08",
          4273 => x"740c7282",
          4274 => x"8cdc0c86",
          4275 => x"3d0d04ff",
          4276 => x"3d0d843d",
          4277 => x"51e6e43f",
          4278 => x"8b52800b",
          4279 => x"828cdc08",
          4280 => x"248b3882",
          4281 => x"8cdc0882",
          4282 => x"8da03480",
          4283 => x"5271828c",
          4284 => x"dc0c833d",
          4285 => x"0d04ef3d",
          4286 => x"0d805393",
          4287 => x"3dd00552",
          4288 => x"943d51e9",
          4289 => x"c13f828c",
          4290 => x"dc085582",
          4291 => x"8cdc0880",
          4292 => x"e0387658",
          4293 => x"6352933d",
          4294 => x"d40551e0",
          4295 => x"8d3f828c",
          4296 => x"dc085582",
          4297 => x"8cdc08bc",
          4298 => x"380280c7",
          4299 => x"05337098",
          4300 => x"2b555673",
          4301 => x"80258938",
          4302 => x"767a9412",
          4303 => x"0c54b239",
          4304 => x"02a20533",
          4305 => x"70842a70",
          4306 => x"81065155",
          4307 => x"5673802e",
          4308 => x"9e38767f",
          4309 => x"53705254",
          4310 => x"dba83f82",
          4311 => x"8cdc0894",
          4312 => x"150c8e39",
          4313 => x"828cdc08",
          4314 => x"842e0981",
          4315 => x"06833885",
          4316 => x"5574828c",
          4317 => x"dc0c933d",
          4318 => x"0d04e43d",
          4319 => x"0d6f6f5b",
          4320 => x"5b807a34",
          4321 => x"80539e3d",
          4322 => x"ffb80552",
          4323 => x"9f3d51e8",
          4324 => x"b53f828c",
          4325 => x"dc085782",
          4326 => x"8cdc0882",
          4327 => x"fc387b43",
          4328 => x"7a7c9411",
          4329 => x"08475558",
          4330 => x"64547380",
          4331 => x"2e81ed38",
          4332 => x"a052933d",
          4333 => x"705255d5",
          4334 => x"ea3f828c",
          4335 => x"dc085782",
          4336 => x"8cdc0882",
          4337 => x"d4386852",
          4338 => x"7b51c9c8",
          4339 => x"3f828cdc",
          4340 => x"0857828c",
          4341 => x"dc0882c1",
          4342 => x"3869527b",
          4343 => x"51daa33f",
          4344 => x"828cdc08",
          4345 => x"45765274",
          4346 => x"51d5b83f",
          4347 => x"828cdc08",
          4348 => x"57828cdc",
          4349 => x"0882a238",
          4350 => x"80527451",
          4351 => x"daeb3f82",
          4352 => x"8cdc0857",
          4353 => x"828cdc08",
          4354 => x"a4386952",
          4355 => x"7b51d9f2",
          4356 => x"3f73828c",
          4357 => x"dc082ea6",
          4358 => x"38765274",
          4359 => x"51d6cf3f",
          4360 => x"828cdc08",
          4361 => x"57828cdc",
          4362 => x"08802ecc",
          4363 => x"3876842e",
          4364 => x"09810686",
          4365 => x"38825781",
          4366 => x"e0397681",
          4367 => x"dc389e3d",
          4368 => x"ffbc0552",
          4369 => x"7451dcc9",
          4370 => x"3f76903d",
          4371 => x"78118111",
          4372 => x"3351565a",
          4373 => x"5673802e",
          4374 => x"913802b9",
          4375 => x"05558116",
          4376 => x"81167033",
          4377 => x"56565673",
          4378 => x"f5388116",
          4379 => x"54737826",
          4380 => x"81903875",
          4381 => x"802e9938",
          4382 => x"78168105",
          4383 => x"55ff186f",
          4384 => x"11ff18ff",
          4385 => x"18585855",
          4386 => x"58743374",
          4387 => x"3475ee38",
          4388 => x"ff186f11",
          4389 => x"5558af74",
          4390 => x"34fe8d39",
          4391 => x"777b2e09",
          4392 => x"81068a38",
          4393 => x"ff186f11",
          4394 => x"5558af74",
          4395 => x"34800b82",
          4396 => x"8da03370",
          4397 => x"842981fa",
          4398 => x"dc057008",
          4399 => x"7033525c",
          4400 => x"56565673",
          4401 => x"762e8d38",
          4402 => x"8116701a",
          4403 => x"70335155",
          4404 => x"5673f538",
          4405 => x"82165473",
          4406 => x"7826a738",
          4407 => x"80557476",
          4408 => x"27913874",
          4409 => x"19547333",
          4410 => x"7a708105",
          4411 => x"5c348115",
          4412 => x"55ec39ba",
          4413 => x"7a708105",
          4414 => x"5c3474ff",
          4415 => x"2e098106",
          4416 => x"85389157",
          4417 => x"94396e18",
          4418 => x"81195954",
          4419 => x"73337a70",
          4420 => x"81055c34",
          4421 => x"7a7826ee",
          4422 => x"38807a34",
          4423 => x"76828cdc",
          4424 => x"0c9e3d0d",
          4425 => x"04f73d0d",
          4426 => x"7b7d8d3d",
          4427 => x"fc055471",
          4428 => x"535755ec",
          4429 => x"bb3f828c",
          4430 => x"dc085382",
          4431 => x"8cdc0882",
          4432 => x"fa389115",
          4433 => x"33537282",
          4434 => x"f2388c15",
          4435 => x"08547376",
          4436 => x"27923890",
          4437 => x"15337081",
          4438 => x"2a708106",
          4439 => x"51545772",
          4440 => x"83387356",
          4441 => x"94150854",
          4442 => x"80709417",
          4443 => x"0c587578",
          4444 => x"2e829738",
          4445 => x"798a1122",
          4446 => x"70892b59",
          4447 => x"51537378",
          4448 => x"2eb73876",
          4449 => x"52ff1651",
          4450 => x"feffd03f",
          4451 => x"828cdc08",
          4452 => x"ff157854",
          4453 => x"70535553",
          4454 => x"feffc03f",
          4455 => x"828cdc08",
          4456 => x"73269638",
          4457 => x"76307075",
          4458 => x"06709418",
          4459 => x"0c777131",
          4460 => x"98180857",
          4461 => x"585153b1",
          4462 => x"39881508",
          4463 => x"5473a638",
          4464 => x"73527451",
          4465 => x"cdca3f82",
          4466 => x"8cdc0854",
          4467 => x"828cdc08",
          4468 => x"812e819a",
          4469 => x"38828cdc",
          4470 => x"08ff2e81",
          4471 => x"9b38828c",
          4472 => x"dc088816",
          4473 => x"0c739816",
          4474 => x"0c73802e",
          4475 => x"819c3876",
          4476 => x"762780dc",
          4477 => x"38757731",
          4478 => x"94160818",
          4479 => x"94170c90",
          4480 => x"16337081",
          4481 => x"2a708106",
          4482 => x"51555a56",
          4483 => x"72802e9a",
          4484 => x"38735274",
          4485 => x"51ccf93f",
          4486 => x"828cdc08",
          4487 => x"54828cdc",
          4488 => x"08943882",
          4489 => x"8cdc0856",
          4490 => x"a7397352",
          4491 => x"7451c784",
          4492 => x"3f828cdc",
          4493 => x"085473ff",
          4494 => x"2ebe3881",
          4495 => x"7427af38",
          4496 => x"79537398",
          4497 => x"140827a6",
          4498 => x"38739816",
          4499 => x"0cffa039",
          4500 => x"94150816",
          4501 => x"94160c75",
          4502 => x"83ff0653",
          4503 => x"72802eaa",
          4504 => x"38735279",
          4505 => x"51c6a33f",
          4506 => x"828cdc08",
          4507 => x"9438820b",
          4508 => x"91163482",
          4509 => x"5380c439",
          4510 => x"810b9116",
          4511 => x"348153bb",
          4512 => x"3975892a",
          4513 => x"828cdc08",
          4514 => x"05589415",
          4515 => x"08548c15",
          4516 => x"08742790",
          4517 => x"38738c16",
          4518 => x"0c901533",
          4519 => x"80c00753",
          4520 => x"72901634",
          4521 => x"7383ff06",
          4522 => x"5372802e",
          4523 => x"8c38779c",
          4524 => x"16082e85",
          4525 => x"38779c16",
          4526 => x"0c805372",
          4527 => x"828cdc0c",
          4528 => x"8b3d0d04",
          4529 => x"f93d0d79",
          4530 => x"56895475",
          4531 => x"802e818a",
          4532 => x"38805389",
          4533 => x"3dfc0552",
          4534 => x"8a3d8405",
          4535 => x"51e1e73f",
          4536 => x"828cdc08",
          4537 => x"55828cdc",
          4538 => x"0880ea38",
          4539 => x"77760c7a",
          4540 => x"527551d8",
          4541 => x"b53f828c",
          4542 => x"dc085582",
          4543 => x"8cdc0880",
          4544 => x"c338ab16",
          4545 => x"3370982b",
          4546 => x"55578074",
          4547 => x"24a23886",
          4548 => x"16337084",
          4549 => x"2a708106",
          4550 => x"51555773",
          4551 => x"802ead38",
          4552 => x"9c160852",
          4553 => x"7751d3da",
          4554 => x"3f828cdc",
          4555 => x"0888170c",
          4556 => x"77548614",
          4557 => x"22841723",
          4558 => x"74527551",
          4559 => x"cee53f82",
          4560 => x"8cdc0855",
          4561 => x"74842e09",
          4562 => x"81068538",
          4563 => x"85558639",
          4564 => x"74802e84",
          4565 => x"3880760c",
          4566 => x"74547382",
          4567 => x"8cdc0c89",
          4568 => x"3d0d04fc",
          4569 => x"3d0d7687",
          4570 => x"3dfc0553",
          4571 => x"705253e7",
          4572 => x"ff3f828c",
          4573 => x"dc088738",
          4574 => x"828cdc08",
          4575 => x"730c863d",
          4576 => x"0d04fb3d",
          4577 => x"0d777989",
          4578 => x"3dfc0554",
          4579 => x"71535654",
          4580 => x"e7de3f82",
          4581 => x"8cdc0853",
          4582 => x"828cdc08",
          4583 => x"80df3874",
          4584 => x"9338828c",
          4585 => x"dc085273",
          4586 => x"51cdf83f",
          4587 => x"828cdc08",
          4588 => x"5380ca39",
          4589 => x"828cdc08",
          4590 => x"527351d3",
          4591 => x"ac3f828c",
          4592 => x"dc085382",
          4593 => x"8cdc0884",
          4594 => x"2e098106",
          4595 => x"85388053",
          4596 => x"8739828c",
          4597 => x"dc08a638",
          4598 => x"74527351",
          4599 => x"d5b33f72",
          4600 => x"527351cf",
          4601 => x"893f828c",
          4602 => x"dc088432",
          4603 => x"70307072",
          4604 => x"079f2c70",
          4605 => x"828cdc08",
          4606 => x"06515154",
          4607 => x"5472828c",
          4608 => x"dc0c873d",
          4609 => x"0d04ee3d",
          4610 => x"0d655780",
          4611 => x"53893d70",
          4612 => x"53963d52",
          4613 => x"56dfaf3f",
          4614 => x"828cdc08",
          4615 => x"55828cdc",
          4616 => x"08b23864",
          4617 => x"527551d6",
          4618 => x"813f828c",
          4619 => x"dc085582",
          4620 => x"8cdc08a0",
          4621 => x"380280cb",
          4622 => x"05337098",
          4623 => x"2b555873",
          4624 => x"80258538",
          4625 => x"86558d39",
          4626 => x"76802e88",
          4627 => x"38765275",
          4628 => x"51d4be3f",
          4629 => x"74828cdc",
          4630 => x"0c943d0d",
          4631 => x"04f03d0d",
          4632 => x"6365555c",
          4633 => x"8053923d",
          4634 => x"ec055293",
          4635 => x"3d51ded6",
          4636 => x"3f828cdc",
          4637 => x"085b828c",
          4638 => x"dc088280",
          4639 => x"387c740c",
          4640 => x"73089811",
          4641 => x"08fe1190",
          4642 => x"13085956",
          4643 => x"58557574",
          4644 => x"26913875",
          4645 => x"7c0c81e4",
          4646 => x"39815b81",
          4647 => x"cc39825b",
          4648 => x"81c73982",
          4649 => x"8cdc0875",
          4650 => x"33555973",
          4651 => x"812e0981",
          4652 => x"06bf3882",
          4653 => x"755f5776",
          4654 => x"52923df0",
          4655 => x"0551c1f4",
          4656 => x"3f828cdc",
          4657 => x"08ff2ed1",
          4658 => x"38828cdc",
          4659 => x"08812ece",
          4660 => x"38828cdc",
          4661 => x"08307082",
          4662 => x"8cdc0807",
          4663 => x"80257a05",
          4664 => x"81197f53",
          4665 => x"595a5498",
          4666 => x"14087726",
          4667 => x"ca3880f9",
          4668 => x"39a41508",
          4669 => x"828cdc08",
          4670 => x"57587598",
          4671 => x"38775281",
          4672 => x"187d5258",
          4673 => x"ffbf8d3f",
          4674 => x"828cdc08",
          4675 => x"5b828cdc",
          4676 => x"0880d638",
          4677 => x"7c703377",
          4678 => x"12ff1a5d",
          4679 => x"52565474",
          4680 => x"822e0981",
          4681 => x"069e38b4",
          4682 => x"1451ffbb",
          4683 => x"cb3f828c",
          4684 => x"dc0883ff",
          4685 => x"ff067030",
          4686 => x"7080251b",
          4687 => x"8219595b",
          4688 => x"51549b39",
          4689 => x"b41451ff",
          4690 => x"bbc53f82",
          4691 => x"8cdc08f0",
          4692 => x"0a067030",
          4693 => x"7080251b",
          4694 => x"8419595b",
          4695 => x"51547583",
          4696 => x"ff067a58",
          4697 => x"5679ff92",
          4698 => x"38787c0c",
          4699 => x"7c799012",
          4700 => x"0c841133",
          4701 => x"81075654",
          4702 => x"74841534",
          4703 => x"7a828cdc",
          4704 => x"0c923d0d",
          4705 => x"04f93d0d",
          4706 => x"798a3dfc",
          4707 => x"05537052",
          4708 => x"57e3dd3f",
          4709 => x"828cdc08",
          4710 => x"56828cdc",
          4711 => x"0881a838",
          4712 => x"91173356",
          4713 => x"7581a038",
          4714 => x"90173370",
          4715 => x"812a7081",
          4716 => x"06515555",
          4717 => x"87557380",
          4718 => x"2e818e38",
          4719 => x"94170854",
          4720 => x"738c1808",
          4721 => x"27818038",
          4722 => x"739b3882",
          4723 => x"8cdc0853",
          4724 => x"88170852",
          4725 => x"7651c48c",
          4726 => x"3f828cdc",
          4727 => x"08748819",
          4728 => x"0c5680c9",
          4729 => x"39981708",
          4730 => x"527651ff",
          4731 => x"bfc63f82",
          4732 => x"8cdc08ff",
          4733 => x"2e098106",
          4734 => x"83388156",
          4735 => x"828cdc08",
          4736 => x"812e0981",
          4737 => x"06853882",
          4738 => x"56a33975",
          4739 => x"a0387754",
          4740 => x"828cdc08",
          4741 => x"98150827",
          4742 => x"94389817",
          4743 => x"0853828c",
          4744 => x"dc085276",
          4745 => x"51c3bd3f",
          4746 => x"828cdc08",
          4747 => x"56941708",
          4748 => x"8c180c90",
          4749 => x"173380c0",
          4750 => x"07547390",
          4751 => x"18347580",
          4752 => x"2e853875",
          4753 => x"91183475",
          4754 => x"5574828c",
          4755 => x"dc0c893d",
          4756 => x"0d04e23d",
          4757 => x"0d8253a0",
          4758 => x"3dffa405",
          4759 => x"52a13d51",
          4760 => x"dae43f82",
          4761 => x"8cdc0855",
          4762 => x"828cdc08",
          4763 => x"81f53878",
          4764 => x"45a13d08",
          4765 => x"52953d70",
          4766 => x"5258d1ae",
          4767 => x"3f828cdc",
          4768 => x"0855828c",
          4769 => x"dc0881db",
          4770 => x"380280fb",
          4771 => x"05337085",
          4772 => x"2a708106",
          4773 => x"51555686",
          4774 => x"557381c7",
          4775 => x"3875982b",
          4776 => x"54807424",
          4777 => x"81bd3802",
          4778 => x"80d60533",
          4779 => x"70810658",
          4780 => x"54875576",
          4781 => x"81ad386b",
          4782 => x"527851cc",
          4783 => x"c53f828c",
          4784 => x"dc087484",
          4785 => x"2a708106",
          4786 => x"51555673",
          4787 => x"802e80d4",
          4788 => x"38785482",
          4789 => x"8cdc0894",
          4790 => x"15082e81",
          4791 => x"8638735a",
          4792 => x"828cdc08",
          4793 => x"5c76528a",
          4794 => x"3d705254",
          4795 => x"c7b53f82",
          4796 => x"8cdc0855",
          4797 => x"828cdc08",
          4798 => x"80e93882",
          4799 => x"8cdc0852",
          4800 => x"7351cce5",
          4801 => x"3f828cdc",
          4802 => x"0855828c",
          4803 => x"dc088638",
          4804 => x"875580cf",
          4805 => x"39828cdc",
          4806 => x"08842e88",
          4807 => x"38828cdc",
          4808 => x"0880c038",
          4809 => x"7751cec2",
          4810 => x"3f828cdc",
          4811 => x"08828cdc",
          4812 => x"08307082",
          4813 => x"8cdc0807",
          4814 => x"80255155",
          4815 => x"5575802e",
          4816 => x"94387380",
          4817 => x"2e8f3880",
          4818 => x"53755277",
          4819 => x"51c1953f",
          4820 => x"828cdc08",
          4821 => x"55748c38",
          4822 => x"7851ffba",
          4823 => x"fe3f828c",
          4824 => x"dc085574",
          4825 => x"828cdc0c",
          4826 => x"a03d0d04",
          4827 => x"e93d0d82",
          4828 => x"53993dc0",
          4829 => x"05529a3d",
          4830 => x"51d8cb3f",
          4831 => x"828cdc08",
          4832 => x"54828cdc",
          4833 => x"0882b038",
          4834 => x"785e6952",
          4835 => x"8e3d7052",
          4836 => x"58cf973f",
          4837 => x"828cdc08",
          4838 => x"54828cdc",
          4839 => x"08863888",
          4840 => x"54829439",
          4841 => x"828cdc08",
          4842 => x"842e0981",
          4843 => x"06828838",
          4844 => x"0280df05",
          4845 => x"3370852a",
          4846 => x"81065155",
          4847 => x"86547481",
          4848 => x"f638785a",
          4849 => x"74528a3d",
          4850 => x"705257c1",
          4851 => x"c33f828c",
          4852 => x"dc087555",
          4853 => x"56828cdc",
          4854 => x"08833887",
          4855 => x"54828cdc",
          4856 => x"08812e09",
          4857 => x"81068338",
          4858 => x"8254828c",
          4859 => x"dc08ff2e",
          4860 => x"09810686",
          4861 => x"38815481",
          4862 => x"b4397381",
          4863 => x"b038828c",
          4864 => x"dc085278",
          4865 => x"51c4a43f",
          4866 => x"828cdc08",
          4867 => x"54828cdc",
          4868 => x"08819a38",
          4869 => x"8b53a052",
          4870 => x"b41951ff",
          4871 => x"b78c3f78",
          4872 => x"54ae0bb4",
          4873 => x"15347854",
          4874 => x"900bbf15",
          4875 => x"348288b2",
          4876 => x"0a5280ca",
          4877 => x"1951ffb6",
          4878 => x"9f3f7553",
          4879 => x"78b41153",
          4880 => x"51c9f83f",
          4881 => x"a05378b4",
          4882 => x"115380d4",
          4883 => x"0551ffb6",
          4884 => x"b63f7854",
          4885 => x"ae0b80d5",
          4886 => x"15347f53",
          4887 => x"7880d411",
          4888 => x"5351c9d7",
          4889 => x"3f785481",
          4890 => x"0b831534",
          4891 => x"7751cba4",
          4892 => x"3f828cdc",
          4893 => x"0854828c",
          4894 => x"dc08b238",
          4895 => x"8288b20a",
          4896 => x"52649605",
          4897 => x"51ffb5d0",
          4898 => x"3f755364",
          4899 => x"527851c9",
          4900 => x"aa3f6454",
          4901 => x"900b8b15",
          4902 => x"34785481",
          4903 => x"0b831534",
          4904 => x"7851ffb8",
          4905 => x"b63f828c",
          4906 => x"dc08548b",
          4907 => x"39805375",
          4908 => x"527651ff",
          4909 => x"beae3f73",
          4910 => x"828cdc0c",
          4911 => x"993d0d04",
          4912 => x"da3d0da9",
          4913 => x"3d840551",
          4914 => x"d2f13f82",
          4915 => x"53a83dff",
          4916 => x"840552a9",
          4917 => x"3d51d5ee",
          4918 => x"3f828cdc",
          4919 => x"0855828c",
          4920 => x"dc0882d3",
          4921 => x"38784da9",
          4922 => x"3d08529d",
          4923 => x"3d705258",
          4924 => x"ccb83f82",
          4925 => x"8cdc0855",
          4926 => x"828cdc08",
          4927 => x"82b93802",
          4928 => x"819b0533",
          4929 => x"81a00654",
          4930 => x"86557382",
          4931 => x"aa38a053",
          4932 => x"a43d0852",
          4933 => x"a83dff88",
          4934 => x"0551ffb4",
          4935 => x"ea3fac53",
          4936 => x"7752923d",
          4937 => x"705254ff",
          4938 => x"b4dd3faa",
          4939 => x"3d085273",
          4940 => x"51cbf73f",
          4941 => x"828cdc08",
          4942 => x"55828cdc",
          4943 => x"08953863",
          4944 => x"6f2e0981",
          4945 => x"06883865",
          4946 => x"a23d082e",
          4947 => x"92388855",
          4948 => x"81e53982",
          4949 => x"8cdc0884",
          4950 => x"2e098106",
          4951 => x"81b83873",
          4952 => x"51c9b13f",
          4953 => x"828cdc08",
          4954 => x"55828cdc",
          4955 => x"0881c838",
          4956 => x"68569353",
          4957 => x"a83dff95",
          4958 => x"05528d16",
          4959 => x"51ffb487",
          4960 => x"3f02af05",
          4961 => x"338b1734",
          4962 => x"8b163370",
          4963 => x"842a7081",
          4964 => x"06515555",
          4965 => x"73893874",
          4966 => x"a0075473",
          4967 => x"8b173478",
          4968 => x"54810b83",
          4969 => x"15348b16",
          4970 => x"3370842a",
          4971 => x"70810651",
          4972 => x"55557380",
          4973 => x"2e80e538",
          4974 => x"6e642e80",
          4975 => x"df387552",
          4976 => x"7851c6be",
          4977 => x"3f828cdc",
          4978 => x"08527851",
          4979 => x"ffb7bb3f",
          4980 => x"8255828c",
          4981 => x"dc08802e",
          4982 => x"80dd3882",
          4983 => x"8cdc0852",
          4984 => x"7851ffb5",
          4985 => x"af3f828c",
          4986 => x"dc087980",
          4987 => x"d4115858",
          4988 => x"55828cdc",
          4989 => x"0880c038",
          4990 => x"81163354",
          4991 => x"73ae2e09",
          4992 => x"81069938",
          4993 => x"63537552",
          4994 => x"7651c6af",
          4995 => x"3f785481",
          4996 => x"0b831534",
          4997 => x"8739828c",
          4998 => x"dc089c38",
          4999 => x"7751c8ca",
          5000 => x"3f828cdc",
          5001 => x"0855828c",
          5002 => x"dc088c38",
          5003 => x"7851ffb5",
          5004 => x"aa3f828c",
          5005 => x"dc085574",
          5006 => x"828cdc0c",
          5007 => x"a83d0d04",
          5008 => x"ed3d0d02",
          5009 => x"80db0533",
          5010 => x"02840580",
          5011 => x"df053357",
          5012 => x"57825395",
          5013 => x"3dd00552",
          5014 => x"963d51d2",
          5015 => x"e93f828c",
          5016 => x"dc085582",
          5017 => x"8cdc0880",
          5018 => x"cf38785a",
          5019 => x"6552953d",
          5020 => x"d40551c9",
          5021 => x"b53f828c",
          5022 => x"dc085582",
          5023 => x"8cdc08b8",
          5024 => x"380280cf",
          5025 => x"053381a0",
          5026 => x"06548655",
          5027 => x"73aa3875",
          5028 => x"a7066171",
          5029 => x"098b1233",
          5030 => x"71067a74",
          5031 => x"06075157",
          5032 => x"5556748b",
          5033 => x"15347854",
          5034 => x"810b8315",
          5035 => x"347851ff",
          5036 => x"b4a93f82",
          5037 => x"8cdc0855",
          5038 => x"74828cdc",
          5039 => x"0c953d0d",
          5040 => x"04ef3d0d",
          5041 => x"64568253",
          5042 => x"933dd005",
          5043 => x"52943d51",
          5044 => x"d1f43f82",
          5045 => x"8cdc0855",
          5046 => x"828cdc08",
          5047 => x"80cb3876",
          5048 => x"58635293",
          5049 => x"3dd40551",
          5050 => x"c8c03f82",
          5051 => x"8cdc0855",
          5052 => x"828cdc08",
          5053 => x"b4380280",
          5054 => x"c7053381",
          5055 => x"a0065486",
          5056 => x"5573a638",
          5057 => x"84162286",
          5058 => x"17227190",
          5059 => x"2b075354",
          5060 => x"961f51ff",
          5061 => x"b0c23f76",
          5062 => x"54810b83",
          5063 => x"15347651",
          5064 => x"ffb3b83f",
          5065 => x"828cdc08",
          5066 => x"5574828c",
          5067 => x"dc0c933d",
          5068 => x"0d04ea3d",
          5069 => x"0d696b5c",
          5070 => x"5a805398",
          5071 => x"3dd00552",
          5072 => x"993d51d1",
          5073 => x"813f828c",
          5074 => x"dc08828c",
          5075 => x"dc083070",
          5076 => x"828cdc08",
          5077 => x"07802551",
          5078 => x"55577980",
          5079 => x"2e818538",
          5080 => x"81707506",
          5081 => x"55557380",
          5082 => x"2e80f938",
          5083 => x"7b5d805f",
          5084 => x"80528d3d",
          5085 => x"705254ff",
          5086 => x"bea93f82",
          5087 => x"8cdc0857",
          5088 => x"828cdc08",
          5089 => x"80d13874",
          5090 => x"527351c3",
          5091 => x"dc3f828c",
          5092 => x"dc085782",
          5093 => x"8cdc08bf",
          5094 => x"38828cdc",
          5095 => x"08828cdc",
          5096 => x"08655b59",
          5097 => x"56781881",
          5098 => x"197b1856",
          5099 => x"59557433",
          5100 => x"74348116",
          5101 => x"568a7827",
          5102 => x"ec388b56",
          5103 => x"751a5480",
          5104 => x"74347580",
          5105 => x"2e9e38ff",
          5106 => x"16701b70",
          5107 => x"33515556",
          5108 => x"73a02ee8",
          5109 => x"388e3976",
          5110 => x"842e0981",
          5111 => x"06863880",
          5112 => x"7a348057",
          5113 => x"76307078",
          5114 => x"07802551",
          5115 => x"547a802e",
          5116 => x"80c13873",
          5117 => x"802ebc38",
          5118 => x"7ba01108",
          5119 => x"5351ffb1",
          5120 => x"933f828c",
          5121 => x"dc085782",
          5122 => x"8cdc08a7",
          5123 => x"387b7033",
          5124 => x"555580c3",
          5125 => x"5673832e",
          5126 => x"8b3880e4",
          5127 => x"5673842e",
          5128 => x"8338a756",
          5129 => x"7515b405",
          5130 => x"51ffade3",
          5131 => x"3f828cdc",
          5132 => x"087b0c76",
          5133 => x"828cdc0c",
          5134 => x"983d0d04",
          5135 => x"e63d0d82",
          5136 => x"539c3dff",
          5137 => x"b805529d",
          5138 => x"3d51cefa",
          5139 => x"3f828cdc",
          5140 => x"08828cdc",
          5141 => x"08565482",
          5142 => x"8cdc0883",
          5143 => x"98388b53",
          5144 => x"a0528b3d",
          5145 => x"705259ff",
          5146 => x"aec03f73",
          5147 => x"6d703370",
          5148 => x"81ff0652",
          5149 => x"5755579f",
          5150 => x"742781bc",
          5151 => x"38785874",
          5152 => x"81ff066d",
          5153 => x"81054e70",
          5154 => x"5255ffaf",
          5155 => x"893f828c",
          5156 => x"dc08802e",
          5157 => x"a5386c70",
          5158 => x"33705357",
          5159 => x"54ffaefd",
          5160 => x"3f828cdc",
          5161 => x"08802e8d",
          5162 => x"3874882b",
          5163 => x"76076d81",
          5164 => x"054e5586",
          5165 => x"39828cdc",
          5166 => x"0855ff9f",
          5167 => x"157083ff",
          5168 => x"ff065154",
          5169 => x"7399268a",
          5170 => x"38e01570",
          5171 => x"83ffff06",
          5172 => x"565480ff",
          5173 => x"75278738",
          5174 => x"81f9ec15",
          5175 => x"33557480",
          5176 => x"2ea33874",
          5177 => x"5281fbec",
          5178 => x"51ffae89",
          5179 => x"3f828cdc",
          5180 => x"08933881",
          5181 => x"ff752788",
          5182 => x"38768926",
          5183 => x"88388b39",
          5184 => x"8a772786",
          5185 => x"38865581",
          5186 => x"ec3981ff",
          5187 => x"75278f38",
          5188 => x"74882a54",
          5189 => x"73787081",
          5190 => x"055a3481",
          5191 => x"17577478",
          5192 => x"7081055a",
          5193 => x"3481176d",
          5194 => x"70337081",
          5195 => x"ff065257",
          5196 => x"5557739f",
          5197 => x"26fec838",
          5198 => x"8b3d3354",
          5199 => x"86557381",
          5200 => x"e52e81b1",
          5201 => x"3876802e",
          5202 => x"993802a7",
          5203 => x"05557615",
          5204 => x"70335154",
          5205 => x"73a02e09",
          5206 => x"81068738",
          5207 => x"ff175776",
          5208 => x"ed387941",
          5209 => x"80438052",
          5210 => x"913d7052",
          5211 => x"55ffbab3",
          5212 => x"3f828cdc",
          5213 => x"0854828c",
          5214 => x"dc0880f7",
          5215 => x"38815274",
          5216 => x"51ffbfe5",
          5217 => x"3f828cdc",
          5218 => x"0854828c",
          5219 => x"dc088d38",
          5220 => x"7680c438",
          5221 => x"6754e574",
          5222 => x"3480c639",
          5223 => x"828cdc08",
          5224 => x"842e0981",
          5225 => x"0680cc38",
          5226 => x"80547674",
          5227 => x"2e80c438",
          5228 => x"81527451",
          5229 => x"ffbdb03f",
          5230 => x"828cdc08",
          5231 => x"54828cdc",
          5232 => x"08b138a0",
          5233 => x"53828cdc",
          5234 => x"08526751",
          5235 => x"ffabdb3f",
          5236 => x"6754880b",
          5237 => x"8b15348b",
          5238 => x"53785267",
          5239 => x"51ffaba7",
          5240 => x"3f795481",
          5241 => x"0b831534",
          5242 => x"7951ffad",
          5243 => x"ee3f828c",
          5244 => x"dc085473",
          5245 => x"5574828c",
          5246 => x"dc0c9c3d",
          5247 => x"0d04f23d",
          5248 => x"0d606202",
          5249 => x"880580cb",
          5250 => x"0533933d",
          5251 => x"fc055572",
          5252 => x"54405e5a",
          5253 => x"d2da3f82",
          5254 => x"8cdc0858",
          5255 => x"828cdc08",
          5256 => x"82bd3891",
          5257 => x"1a335877",
          5258 => x"82b5387c",
          5259 => x"802e9738",
          5260 => x"8c1a0859",
          5261 => x"78903890",
          5262 => x"1a337081",
          5263 => x"2a708106",
          5264 => x"51555573",
          5265 => x"90388754",
          5266 => x"82973982",
          5267 => x"58829039",
          5268 => x"8158828b",
          5269 => x"397e8a11",
          5270 => x"2270892b",
          5271 => x"70557f54",
          5272 => x"565656fe",
          5273 => x"e5f53fff",
          5274 => x"147d0670",
          5275 => x"30707207",
          5276 => x"9f2a828c",
          5277 => x"dc08058c",
          5278 => x"19087c40",
          5279 => x"5a5d5555",
          5280 => x"81772788",
          5281 => x"38981608",
          5282 => x"77268338",
          5283 => x"82577677",
          5284 => x"56598056",
          5285 => x"74527951",
          5286 => x"ffae993f",
          5287 => x"81157f55",
          5288 => x"55981408",
          5289 => x"75268338",
          5290 => x"8255828c",
          5291 => x"dc08812e",
          5292 => x"ff993882",
          5293 => x"8cdc08ff",
          5294 => x"2eff9538",
          5295 => x"828cdc08",
          5296 => x"8e388116",
          5297 => x"56757b2e",
          5298 => x"09810687",
          5299 => x"38933974",
          5300 => x"59805674",
          5301 => x"772e0981",
          5302 => x"06ffb938",
          5303 => x"875880ff",
          5304 => x"397d802e",
          5305 => x"ba38787b",
          5306 => x"55557a80",
          5307 => x"2eb43881",
          5308 => x"15567381",
          5309 => x"2e098106",
          5310 => x"8338ff56",
          5311 => x"75537452",
          5312 => x"7e51ffaf",
          5313 => x"a83f828c",
          5314 => x"dc085882",
          5315 => x"8cdc0880",
          5316 => x"ce387481",
          5317 => x"16ff1656",
          5318 => x"565c73d3",
          5319 => x"388439ff",
          5320 => x"195c7e7c",
          5321 => x"8c120c55",
          5322 => x"7d802eb3",
          5323 => x"3878881b",
          5324 => x"0c7c8c1b",
          5325 => x"0c901a33",
          5326 => x"80c00754",
          5327 => x"73901b34",
          5328 => x"981508fe",
          5329 => x"05901608",
          5330 => x"57547574",
          5331 => x"26913875",
          5332 => x"7b319016",
          5333 => x"0c841533",
          5334 => x"81075473",
          5335 => x"84163477",
          5336 => x"5473828c",
          5337 => x"dc0c903d",
          5338 => x"0d04e93d",
          5339 => x"0d6b6d02",
          5340 => x"880580eb",
          5341 => x"05339d3d",
          5342 => x"545a5c59",
          5343 => x"c5bd3f8b",
          5344 => x"56800b82",
          5345 => x"8cdc0824",
          5346 => x"8bf83882",
          5347 => x"8cdc0884",
          5348 => x"29828d8c",
          5349 => x"05700851",
          5350 => x"5574802e",
          5351 => x"84388075",
          5352 => x"34828cdc",
          5353 => x"0881ff06",
          5354 => x"5f81527e",
          5355 => x"51ffa0d0",
          5356 => x"3f828cdc",
          5357 => x"0881ff06",
          5358 => x"70810656",
          5359 => x"57835674",
          5360 => x"8bc03876",
          5361 => x"822a7081",
          5362 => x"0651558a",
          5363 => x"56748bb2",
          5364 => x"38993dfc",
          5365 => x"05538352",
          5366 => x"7e51ffa4",
          5367 => x"f03f828c",
          5368 => x"dc089938",
          5369 => x"67557480",
          5370 => x"2e923874",
          5371 => x"82808026",
          5372 => x"8b38ff15",
          5373 => x"75065574",
          5374 => x"802e8338",
          5375 => x"81487880",
          5376 => x"2e873884",
          5377 => x"80792692",
          5378 => x"38788180",
          5379 => x"0a268b38",
          5380 => x"ff197906",
          5381 => x"5574802e",
          5382 => x"86389356",
          5383 => x"8ae43978",
          5384 => x"892a6e89",
          5385 => x"2a70892b",
          5386 => x"77594843",
          5387 => x"597a8338",
          5388 => x"81566130",
          5389 => x"70802577",
          5390 => x"07515591",
          5391 => x"56748ac2",
          5392 => x"38993df8",
          5393 => x"05538152",
          5394 => x"7e51ffa4",
          5395 => x"803f8156",
          5396 => x"828cdc08",
          5397 => x"8aac3877",
          5398 => x"832a7077",
          5399 => x"06828cdc",
          5400 => x"08435645",
          5401 => x"748338bf",
          5402 => x"4166558e",
          5403 => x"56607526",
          5404 => x"8a903874",
          5405 => x"61317048",
          5406 => x"5580ff75",
          5407 => x"278a8338",
          5408 => x"93567881",
          5409 => x"802689fa",
          5410 => x"3877812a",
          5411 => x"70810656",
          5412 => x"4374802e",
          5413 => x"95387787",
          5414 => x"06557482",
          5415 => x"2e838d38",
          5416 => x"77810655",
          5417 => x"74802e83",
          5418 => x"83387781",
          5419 => x"06559356",
          5420 => x"825e7480",
          5421 => x"2e89cb38",
          5422 => x"785a7d83",
          5423 => x"2e098106",
          5424 => x"80e13878",
          5425 => x"ae386691",
          5426 => x"2a57810b",
          5427 => x"81fc9022",
          5428 => x"565a7480",
          5429 => x"2e9d3874",
          5430 => x"77269838",
          5431 => x"81fc9056",
          5432 => x"79108217",
          5433 => x"70225757",
          5434 => x"5a74802e",
          5435 => x"86387675",
          5436 => x"27ee3879",
          5437 => x"526651fe",
          5438 => x"e0e13f82",
          5439 => x"8cdc0884",
          5440 => x"29848705",
          5441 => x"70892a5e",
          5442 => x"55a05c80",
          5443 => x"0b828cdc",
          5444 => x"08fc808a",
          5445 => x"055644fd",
          5446 => x"fff00a75",
          5447 => x"2780ec38",
          5448 => x"88d33978",
          5449 => x"ae38668c",
          5450 => x"2a57810b",
          5451 => x"81fc8022",
          5452 => x"565a7480",
          5453 => x"2e9d3874",
          5454 => x"77269838",
          5455 => x"81fc8056",
          5456 => x"79108217",
          5457 => x"70225757",
          5458 => x"5a74802e",
          5459 => x"86387675",
          5460 => x"27ee3879",
          5461 => x"526651fe",
          5462 => x"e0813f82",
          5463 => x"8cdc0810",
          5464 => x"84055782",
          5465 => x"8cdc089f",
          5466 => x"f5269638",
          5467 => x"810b828c",
          5468 => x"dc081082",
          5469 => x"8cdc0805",
          5470 => x"7111722a",
          5471 => x"83055956",
          5472 => x"5e83ff17",
          5473 => x"892a5d81",
          5474 => x"5ca04460",
          5475 => x"1c7d1165",
          5476 => x"05697012",
          5477 => x"ff057130",
          5478 => x"70720674",
          5479 => x"315c5259",
          5480 => x"5759407d",
          5481 => x"832e0981",
          5482 => x"06893876",
          5483 => x"1c601841",
          5484 => x"5c843976",
          5485 => x"1d5d7990",
          5486 => x"29187062",
          5487 => x"31685851",
          5488 => x"55747626",
          5489 => x"87af3875",
          5490 => x"7c317d31",
          5491 => x"7a537065",
          5492 => x"315255fe",
          5493 => x"df853f82",
          5494 => x"8cdc0858",
          5495 => x"7d832e09",
          5496 => x"81069b38",
          5497 => x"828cdc08",
          5498 => x"83fff526",
          5499 => x"80dd3878",
          5500 => x"87833879",
          5501 => x"812a5978",
          5502 => x"fdbe3886",
          5503 => x"f8397d82",
          5504 => x"2e098106",
          5505 => x"80c53883",
          5506 => x"fff50b82",
          5507 => x"8cdc0827",
          5508 => x"a038788f",
          5509 => x"38791a55",
          5510 => x"7480c026",
          5511 => x"86387459",
          5512 => x"fd963962",
          5513 => x"81065574",
          5514 => x"802e8f38",
          5515 => x"835efd88",
          5516 => x"39828cdc",
          5517 => x"089ff526",
          5518 => x"92387886",
          5519 => x"b838791a",
          5520 => x"59818079",
          5521 => x"27fcf138",
          5522 => x"86ab3980",
          5523 => x"557d812e",
          5524 => x"09810683",
          5525 => x"387d559f",
          5526 => x"f578278b",
          5527 => x"38748106",
          5528 => x"558e5674",
          5529 => x"869c3884",
          5530 => x"80538052",
          5531 => x"7a51ffa2",
          5532 => x"b93f8b53",
          5533 => x"81faa852",
          5534 => x"7a51ffa2",
          5535 => x"8a3f8480",
          5536 => x"528b1b51",
          5537 => x"ffa1b33f",
          5538 => x"798d1c34",
          5539 => x"7b83ffff",
          5540 => x"06528e1b",
          5541 => x"51ffa1a2",
          5542 => x"3f810b90",
          5543 => x"1c347d83",
          5544 => x"32703070",
          5545 => x"962a8480",
          5546 => x"06545155",
          5547 => x"911b51ff",
          5548 => x"a1883f66",
          5549 => x"557483ff",
          5550 => x"ff269038",
          5551 => x"7483ffff",
          5552 => x"0652931b",
          5553 => x"51ffa0f2",
          5554 => x"3f8a3974",
          5555 => x"52a01b51",
          5556 => x"ffa1853f",
          5557 => x"f80b951c",
          5558 => x"34bf5298",
          5559 => x"1b51ffa0",
          5560 => x"d93f81ff",
          5561 => x"529a1b51",
          5562 => x"ffa0cf3f",
          5563 => x"60529c1b",
          5564 => x"51ffa0e4",
          5565 => x"3f7d832e",
          5566 => x"09810680",
          5567 => x"cb388288",
          5568 => x"b20a5280",
          5569 => x"c31b51ff",
          5570 => x"a0ce3f7c",
          5571 => x"52a41b51",
          5572 => x"ffa0c53f",
          5573 => x"8252ac1b",
          5574 => x"51ffa0bc",
          5575 => x"3f8152b0",
          5576 => x"1b51ffa0",
          5577 => x"953f8652",
          5578 => x"b21b51ff",
          5579 => x"a08c3fff",
          5580 => x"800b80c0",
          5581 => x"1c34a90b",
          5582 => x"80c21c34",
          5583 => x"935381fa",
          5584 => x"b45280c7",
          5585 => x"1b51ae39",
          5586 => x"8288b20a",
          5587 => x"52a71b51",
          5588 => x"ffa0853f",
          5589 => x"7c83ffff",
          5590 => x"0652961b",
          5591 => x"51ff9fda",
          5592 => x"3fff800b",
          5593 => x"a41c34a9",
          5594 => x"0ba61c34",
          5595 => x"935381fa",
          5596 => x"c852ab1b",
          5597 => x"51ffa08f",
          5598 => x"3f82d4d5",
          5599 => x"5283fe1b",
          5600 => x"705259ff",
          5601 => x"9fb43f81",
          5602 => x"5460537a",
          5603 => x"527e51ff",
          5604 => x"9bd73f81",
          5605 => x"56828cdc",
          5606 => x"0883e738",
          5607 => x"7d832e09",
          5608 => x"810680ee",
          5609 => x"38755460",
          5610 => x"8605537a",
          5611 => x"527e51ff",
          5612 => x"9bb73f84",
          5613 => x"80538052",
          5614 => x"7a51ff9f",
          5615 => x"ed3f848b",
          5616 => x"85a4d252",
          5617 => x"7a51ff9f",
          5618 => x"8f3f868a",
          5619 => x"85e4f252",
          5620 => x"83e41b51",
          5621 => x"ff9f813f",
          5622 => x"ff185283",
          5623 => x"e81b51ff",
          5624 => x"9ef63f82",
          5625 => x"5283ec1b",
          5626 => x"51ff9eec",
          5627 => x"3f82d4d5",
          5628 => x"527851ff",
          5629 => x"9ec43f75",
          5630 => x"54608705",
          5631 => x"537a527e",
          5632 => x"51ff9ae5",
          5633 => x"3f755460",
          5634 => x"16537a52",
          5635 => x"7e51ff9a",
          5636 => x"d83f6553",
          5637 => x"80527a51",
          5638 => x"ff9f8f3f",
          5639 => x"7f568058",
          5640 => x"7d832e09",
          5641 => x"81069a38",
          5642 => x"f8527a51",
          5643 => x"ff9ea93f",
          5644 => x"ff52841b",
          5645 => x"51ff9ea0",
          5646 => x"3ff00a52",
          5647 => x"881b5191",
          5648 => x"3987ffff",
          5649 => x"f8557d81",
          5650 => x"2e8338f8",
          5651 => x"5574527a",
          5652 => x"51ff9e84",
          5653 => x"3f7c5561",
          5654 => x"57746226",
          5655 => x"83387457",
          5656 => x"76547553",
          5657 => x"7a527e51",
          5658 => x"ff99fe3f",
          5659 => x"828cdc08",
          5660 => x"82873884",
          5661 => x"8053828c",
          5662 => x"dc08527a",
          5663 => x"51ff9eaa",
          5664 => x"3f761675",
          5665 => x"78315656",
          5666 => x"74cd3881",
          5667 => x"18587780",
          5668 => x"2eff8d38",
          5669 => x"79557d83",
          5670 => x"2e833863",
          5671 => x"55615774",
          5672 => x"62268338",
          5673 => x"74577654",
          5674 => x"75537a52",
          5675 => x"7e51ff99",
          5676 => x"b83f828c",
          5677 => x"dc0881c1",
          5678 => x"38761675",
          5679 => x"78315656",
          5680 => x"74db388c",
          5681 => x"567d832e",
          5682 => x"93388656",
          5683 => x"6683ffff",
          5684 => x"268a3884",
          5685 => x"567d822e",
          5686 => x"83388156",
          5687 => x"64810658",
          5688 => x"7780fe38",
          5689 => x"84805377",
          5690 => x"527a51ff",
          5691 => x"9dbc3f82",
          5692 => x"d4d55278",
          5693 => x"51ff9cc2",
          5694 => x"3f83be1b",
          5695 => x"55777534",
          5696 => x"810b8116",
          5697 => x"34810b82",
          5698 => x"16347783",
          5699 => x"16347584",
          5700 => x"16346067",
          5701 => x"055680fd",
          5702 => x"c1527551",
          5703 => x"fed8bc3f",
          5704 => x"fe0b8516",
          5705 => x"34828cdc",
          5706 => x"08822abf",
          5707 => x"07567586",
          5708 => x"1634828c",
          5709 => x"dc088716",
          5710 => x"34605283",
          5711 => x"c61b51ff",
          5712 => x"9c963f66",
          5713 => x"5283ca1b",
          5714 => x"51ff9c8c",
          5715 => x"3f815477",
          5716 => x"537a527e",
          5717 => x"51ff9891",
          5718 => x"3f815682",
          5719 => x"8cdc08a2",
          5720 => x"38805380",
          5721 => x"527e51ff",
          5722 => x"99e33f81",
          5723 => x"56828cdc",
          5724 => x"08903889",
          5725 => x"398e568a",
          5726 => x"39815686",
          5727 => x"39828cdc",
          5728 => x"08567582",
          5729 => x"8cdc0c99",
          5730 => x"3d0d04f5",
          5731 => x"3d0d7d60",
          5732 => x"5b598079",
          5733 => x"60ff055a",
          5734 => x"57577678",
          5735 => x"25b4388d",
          5736 => x"3df81155",
          5737 => x"558153fc",
          5738 => x"15527951",
          5739 => x"c9dc3f7a",
          5740 => x"812e0981",
          5741 => x"069c388c",
          5742 => x"3d335574",
          5743 => x"8d2edb38",
          5744 => x"74767081",
          5745 => x"05583481",
          5746 => x"1757748a",
          5747 => x"2e098106",
          5748 => x"c9388076",
          5749 => x"34785576",
          5750 => x"83387655",
          5751 => x"74828cdc",
          5752 => x"0c8d3d0d",
          5753 => x"04f73d0d",
          5754 => x"7b028405",
          5755 => x"b3053359",
          5756 => x"57778a2e",
          5757 => x"09810687",
          5758 => x"388d5276",
          5759 => x"51e73f84",
          5760 => x"17085680",
          5761 => x"7624be38",
          5762 => x"88170877",
          5763 => x"178c0556",
          5764 => x"59777534",
          5765 => x"811656bb",
          5766 => x"7625a138",
          5767 => x"8b3dfc05",
          5768 => x"5475538c",
          5769 => x"17527608",
          5770 => x"51cbdc3f",
          5771 => x"79763270",
          5772 => x"30707207",
          5773 => x"9f2a7030",
          5774 => x"53515656",
          5775 => x"7584180c",
          5776 => x"81198818",
          5777 => x"0c8b3d0d",
          5778 => x"04f93d0d",
          5779 => x"79841108",
          5780 => x"56568075",
          5781 => x"24a73889",
          5782 => x"3dfc0554",
          5783 => x"74538c16",
          5784 => x"52750851",
          5785 => x"cba13f82",
          5786 => x"8cdc0891",
          5787 => x"38841608",
          5788 => x"782e0981",
          5789 => x"06873888",
          5790 => x"16085583",
          5791 => x"39ff5574",
          5792 => x"828cdc0c",
          5793 => x"893d0d04",
          5794 => x"fd3d0d75",
          5795 => x"5480cc53",
          5796 => x"80527351",
          5797 => x"ff9a933f",
          5798 => x"76740c85",
          5799 => x"3d0d04ea",
          5800 => x"3d0d0280",
          5801 => x"e305336a",
          5802 => x"53863d70",
          5803 => x"535454d8",
          5804 => x"3f735272",
          5805 => x"51feae3f",
          5806 => x"7251ff8d",
          5807 => x"3f983d0d",
          5808 => x"04f83d0d",
          5809 => x"7a700870",
          5810 => x"56565974",
          5811 => x"802e80e1",
          5812 => x"388c3977",
          5813 => x"15790c85",
          5814 => x"16335480",
          5815 => x"d4397433",
          5816 => x"5473a02e",
          5817 => x"09810686",
          5818 => x"38811555",
          5819 => x"f1398057",
          5820 => x"76902982",
          5821 => x"89cc0570",
          5822 => x"085256fe",
          5823 => x"daf03f82",
          5824 => x"8cdc0882",
          5825 => x"8cdc0854",
          5826 => x"75537608",
          5827 => x"5258fedb",
          5828 => x"be3f828c",
          5829 => x"dc088b38",
          5830 => x"84163354",
          5831 => x"73812eff",
          5832 => x"b2388117",
          5833 => x"7081ff06",
          5834 => x"58549877",
          5835 => x"27c238ff",
          5836 => x"5473828c",
          5837 => x"dc0c8a3d",
          5838 => x"0d04ff3d",
          5839 => x"0d735271",
          5840 => x"9326818e",
          5841 => x"38718429",
          5842 => x"81f19405",
          5843 => x"52710804",
          5844 => x"81fdc851",
          5845 => x"81803981",
          5846 => x"fdd45180",
          5847 => x"f93981fd",
          5848 => x"e85180f2",
          5849 => x"3981fdfc",
          5850 => x"5180eb39",
          5851 => x"81fe8c51",
          5852 => x"80e43981",
          5853 => x"fe9c5180",
          5854 => x"dd3981fe",
          5855 => x"b05180d6",
          5856 => x"3981fec0",
          5857 => x"5180cf39",
          5858 => x"81fed851",
          5859 => x"80c83981",
          5860 => x"fef05180",
          5861 => x"c13981ff",
          5862 => x"8851bb39",
          5863 => x"81ffa451",
          5864 => x"b53981ff",
          5865 => x"b851af39",
          5866 => x"81ffe451",
          5867 => x"a93981ff",
          5868 => x"f851a339",
          5869 => x"82809851",
          5870 => x"9d398280",
          5871 => x"ac519739",
          5872 => x"8280c451",
          5873 => x"91398280",
          5874 => x"dc518b39",
          5875 => x"8280f451",
          5876 => x"85398281",
          5877 => x"8051fef2",
          5878 => x"ae3f833d",
          5879 => x"0d04fb3d",
          5880 => x"0d777956",
          5881 => x"567487e7",
          5882 => x"268a3874",
          5883 => x"527587e8",
          5884 => x"29519139",
          5885 => x"87e85274",
          5886 => x"51fed2df",
          5887 => x"3f828cdc",
          5888 => x"08527551",
          5889 => x"fed2d43f",
          5890 => x"828cdc08",
          5891 => x"54795375",
          5892 => x"52828190",
          5893 => x"51fef7d3",
          5894 => x"3f873d0d",
          5895 => x"04ec3d0d",
          5896 => x"66028405",
          5897 => x"80e30533",
          5898 => x"5b578068",
          5899 => x"7830707a",
          5900 => x"07732551",
          5901 => x"57595978",
          5902 => x"567787ff",
          5903 => x"26833881",
          5904 => x"56747607",
          5905 => x"7081ff06",
          5906 => x"51559356",
          5907 => x"74818038",
          5908 => x"81537652",
          5909 => x"8c3d7052",
          5910 => x"56ffbfc9",
          5911 => x"3f828cdc",
          5912 => x"0857828c",
          5913 => x"dc08b838",
          5914 => x"828cdc08",
          5915 => x"87c09888",
          5916 => x"0c828cdc",
          5917 => x"0859963d",
          5918 => x"d4055484",
          5919 => x"80537752",
          5920 => x"7551c486",
          5921 => x"3f828cdc",
          5922 => x"0857828c",
          5923 => x"dc089038",
          5924 => x"7a557480",
          5925 => x"2e893874",
          5926 => x"19751959",
          5927 => x"59d83996",
          5928 => x"3dd80551",
          5929 => x"cbf03f76",
          5930 => x"30707807",
          5931 => x"80257b30",
          5932 => x"709f2a72",
          5933 => x"06515751",
          5934 => x"5674802e",
          5935 => x"90388281",
          5936 => x"b45387c0",
          5937 => x"98880852",
          5938 => x"7851fe92",
          5939 => x"3f765675",
          5940 => x"828cdc0c",
          5941 => x"963d0d04",
          5942 => x"f93d0d7b",
          5943 => x"028405b3",
          5944 => x"05335758",
          5945 => x"ff578053",
          5946 => x"7a527951",
          5947 => x"feaf3f82",
          5948 => x"8cdc08a4",
          5949 => x"3875802e",
          5950 => x"88387581",
          5951 => x"2e983898",
          5952 => x"3960557f",
          5953 => x"54828cdc",
          5954 => x"537e527d",
          5955 => x"51772d82",
          5956 => x"8cdc0857",
          5957 => x"83397704",
          5958 => x"76828cdc",
          5959 => x"0c893d0d",
          5960 => x"04f33d0d",
          5961 => x"7f616302",
          5962 => x"8c0580cf",
          5963 => x"05337373",
          5964 => x"1568415f",
          5965 => x"5c5c5e5e",
          5966 => x"5e7a5282",
          5967 => x"81bc51fe",
          5968 => x"f5a93f82",
          5969 => x"81c451fe",
          5970 => x"efbd3f80",
          5971 => x"55747927",
          5972 => x"80fc387b",
          5973 => x"902e8938",
          5974 => x"7ba02ea7",
          5975 => x"3880c639",
          5976 => x"74185372",
          5977 => x"7a278e38",
          5978 => x"72225282",
          5979 => x"81c851fe",
          5980 => x"f4f93f89",
          5981 => x"398281d4",
          5982 => x"51feef8b",
          5983 => x"3f821555",
          5984 => x"80c33974",
          5985 => x"1853727a",
          5986 => x"278e3872",
          5987 => x"08528281",
          5988 => x"bc51fef4",
          5989 => x"d63f8939",
          5990 => x"8281d051",
          5991 => x"feeee83f",
          5992 => x"841555a1",
          5993 => x"39741853",
          5994 => x"727a278e",
          5995 => x"38723352",
          5996 => x"8281dc51",
          5997 => x"fef4b43f",
          5998 => x"89398281",
          5999 => x"e451feee",
          6000 => x"c63f8115",
          6001 => x"55a051fe",
          6002 => x"ede03fff",
          6003 => x"80398281",
          6004 => x"e851feee",
          6005 => x"b23f8055",
          6006 => x"747927bc",
          6007 => x"38741870",
          6008 => x"33555380",
          6009 => x"56727a27",
          6010 => x"83388156",
          6011 => x"80539f74",
          6012 => x"27833881",
          6013 => x"53757306",
          6014 => x"7081ff06",
          6015 => x"51537280",
          6016 => x"2e8b3873",
          6017 => x"80fe2685",
          6018 => x"38735183",
          6019 => x"39a051fe",
          6020 => x"ed983f81",
          6021 => x"1555c139",
          6022 => x"8281ec51",
          6023 => x"feede83f",
          6024 => x"7818791c",
          6025 => x"5c58fede",
          6026 => x"d53f828c",
          6027 => x"dc08982b",
          6028 => x"70982c51",
          6029 => x"5776a02e",
          6030 => x"098106ab",
          6031 => x"38fedebe",
          6032 => x"3f828cdc",
          6033 => x"08982b70",
          6034 => x"982c70a0",
          6035 => x"32703072",
          6036 => x"9b327030",
          6037 => x"70720773",
          6038 => x"75070651",
          6039 => x"58585957",
          6040 => x"51578073",
          6041 => x"24d73876",
          6042 => x"9b2e0981",
          6043 => x"06853880",
          6044 => x"538c397c",
          6045 => x"1e537278",
          6046 => x"26fdbe38",
          6047 => x"ff537282",
          6048 => x"8cdc0c8f",
          6049 => x"3d0d04fc",
          6050 => x"3d0d029b",
          6051 => x"05338281",
          6052 => x"f0538281",
          6053 => x"f45255fe",
          6054 => x"f2d13f82",
          6055 => x"888c2251",
          6056 => x"fee7963f",
          6057 => x"82828054",
          6058 => x"82828c53",
          6059 => x"82888d33",
          6060 => x"52828294",
          6061 => x"51fef2b3",
          6062 => x"3f74802e",
          6063 => x"8538fee2",
          6064 => x"e13f863d",
          6065 => x"0d04fe3d",
          6066 => x"0d87c096",
          6067 => x"800853fe",
          6068 => x"e7b13f81",
          6069 => x"51fed9ba",
          6070 => x"3f8282b0",
          6071 => x"51fedbb2",
          6072 => x"3f8051fe",
          6073 => x"d9ac3f72",
          6074 => x"812a7081",
          6075 => x"06515271",
          6076 => x"802e9538",
          6077 => x"8151fed9",
          6078 => x"993f8282",
          6079 => x"c851fedb",
          6080 => x"913f8051",
          6081 => x"fed98b3f",
          6082 => x"72822a70",
          6083 => x"81065152",
          6084 => x"71802e95",
          6085 => x"388151fe",
          6086 => x"d8f83f82",
          6087 => x"82dc51fe",
          6088 => x"daf03f80",
          6089 => x"51fed8ea",
          6090 => x"3f72832a",
          6091 => x"70810651",
          6092 => x"5271802e",
          6093 => x"95388151",
          6094 => x"fed8d73f",
          6095 => x"8282ec51",
          6096 => x"fedacf3f",
          6097 => x"8051fed8",
          6098 => x"c93f7284",
          6099 => x"2a708106",
          6100 => x"51527180",
          6101 => x"2e953881",
          6102 => x"51fed8b6",
          6103 => x"3f828380",
          6104 => x"51fedaae",
          6105 => x"3f8051fe",
          6106 => x"d8a83f72",
          6107 => x"852a7081",
          6108 => x"06515271",
          6109 => x"802e9538",
          6110 => x"8151fed8",
          6111 => x"953f8283",
          6112 => x"9451feda",
          6113 => x"8d3f8051",
          6114 => x"fed8873f",
          6115 => x"72862a70",
          6116 => x"81065152",
          6117 => x"71802e95",
          6118 => x"388151fe",
          6119 => x"d7f43f82",
          6120 => x"83a851fe",
          6121 => x"d9ec3f80",
          6122 => x"51fed7e6",
          6123 => x"3f72872a",
          6124 => x"70810651",
          6125 => x"5271802e",
          6126 => x"95388151",
          6127 => x"fed7d33f",
          6128 => x"8283bc51",
          6129 => x"fed9cb3f",
          6130 => x"8051fed7",
          6131 => x"c53f7288",
          6132 => x"2a708106",
          6133 => x"51527180",
          6134 => x"2e953881",
          6135 => x"51fed7b2",
          6136 => x"3f8283d0",
          6137 => x"51fed9aa",
          6138 => x"3f8051fe",
          6139 => x"d7a43ffe",
          6140 => x"e5993f84",
          6141 => x"3d0d04fb",
          6142 => x"3d0d7702",
          6143 => x"8405a305",
          6144 => x"33705556",
          6145 => x"56805275",
          6146 => x"51fecee2",
          6147 => x"3f8289c8",
          6148 => x"335473a7",
          6149 => x"38815382",
          6150 => x"84905282",
          6151 => x"a3f451ff",
          6152 => x"b8833f82",
          6153 => x"8cdc0830",
          6154 => x"70828cdc",
          6155 => x"08078025",
          6156 => x"82713151",
          6157 => x"51547382",
          6158 => x"89c83482",
          6159 => x"89c83354",
          6160 => x"73812e09",
          6161 => x"8106ac38",
          6162 => x"82a3f453",
          6163 => x"74527551",
          6164 => x"f2b93f82",
          6165 => x"8cdc0880",
          6166 => x"2e8c3882",
          6167 => x"8cdc0851",
          6168 => x"fee9a43f",
          6169 => x"8e3982a3",
          6170 => x"f451c4aa",
          6171 => x"3f820b82",
          6172 => x"89c83482",
          6173 => x"89c83354",
          6174 => x"73822e09",
          6175 => x"81068938",
          6176 => x"74527551",
          6177 => x"fefae43f",
          6178 => x"800b828c",
          6179 => x"dc0c873d",
          6180 => x"0d04ce3d",
          6181 => x"0d807071",
          6182 => x"82a3f00c",
          6183 => x"5f5d8152",
          6184 => x"7c51ff86",
          6185 => x"db3f828c",
          6186 => x"dc0881ff",
          6187 => x"0659787d",
          6188 => x"2e098106",
          6189 => x"a2388284",
          6190 => x"a052963d",
          6191 => x"705259fe",
          6192 => x"eebf3f7c",
          6193 => x"53785282",
          6194 => x"8ea051ff",
          6195 => x"b5f63f82",
          6196 => x"8cdc087d",
          6197 => x"2e883882",
          6198 => x"84a4518d",
          6199 => x"bc398170",
          6200 => x"5f5d8284",
          6201 => x"dc51fee8",
          6202 => x"9e3f963d",
          6203 => x"70465a80",
          6204 => x"f8527951",
          6205 => x"fe813fb4",
          6206 => x"3dff8405",
          6207 => x"51f3c23f",
          6208 => x"828cdc08",
          6209 => x"902b7090",
          6210 => x"2c515978",
          6211 => x"80c22e87",
          6212 => x"b3387880",
          6213 => x"c224b238",
          6214 => x"78bd2e81",
          6215 => x"d53878bd",
          6216 => x"24903878",
          6217 => x"802effba",
          6218 => x"3878bc2e",
          6219 => x"80da388a",
          6220 => x"e9397880",
          6221 => x"c02e83a1",
          6222 => x"387880c0",
          6223 => x"2485dd38",
          6224 => x"78bf2e82",
          6225 => x"92388ad2",
          6226 => x"397880f9",
          6227 => x"2e89ea38",
          6228 => x"7880f924",
          6229 => x"92387880",
          6230 => x"c32e8898",
          6231 => x"387880f8",
          6232 => x"2e89b138",
          6233 => x"8ab43978",
          6234 => x"81832e8a",
          6235 => x"99387881",
          6236 => x"83248b38",
          6237 => x"7881822e",
          6238 => x"89fd388a",
          6239 => x"9d397881",
          6240 => x"852e8a8f",
          6241 => x"388a9339",
          6242 => x"b43dff80",
          6243 => x"1153ff84",
          6244 => x"0551feee",
          6245 => x"cb3f828c",
          6246 => x"dc08802e",
          6247 => x"fec438b4",
          6248 => x"3dfefc11",
          6249 => x"53ff8405",
          6250 => x"51feeeb4",
          6251 => x"3f828cdc",
          6252 => x"08802efe",
          6253 => x"ad38b43d",
          6254 => x"fef81153",
          6255 => x"ff840551",
          6256 => x"feee9d3f",
          6257 => x"828cdc08",
          6258 => x"8638828c",
          6259 => x"dc084282",
          6260 => x"84e051fe",
          6261 => x"e6b13f63",
          6262 => x"635c5a79",
          6263 => x"7b2781f2",
          6264 => x"38615978",
          6265 => x"7a708405",
          6266 => x"5c0c7a7a",
          6267 => x"26f53881",
          6268 => x"e139b43d",
          6269 => x"ff801153",
          6270 => x"ff840551",
          6271 => x"feede13f",
          6272 => x"828cdc08",
          6273 => x"802efdda",
          6274 => x"38b43dfe",
          6275 => x"fc1153ff",
          6276 => x"840551fe",
          6277 => x"edca3f82",
          6278 => x"8cdc0880",
          6279 => x"2efdc338",
          6280 => x"b43dfef8",
          6281 => x"1153ff84",
          6282 => x"0551feed",
          6283 => x"b33f828c",
          6284 => x"dc08802e",
          6285 => x"fdac3882",
          6286 => x"84f051fe",
          6287 => x"e5c93f63",
          6288 => x"5a796327",
          6289 => x"818c3861",
          6290 => x"59797081",
          6291 => x"055b3379",
          6292 => x"34618105",
          6293 => x"42eb39b4",
          6294 => x"3dff8011",
          6295 => x"53ff8405",
          6296 => x"51feecfc",
          6297 => x"3f828cdc",
          6298 => x"08802efc",
          6299 => x"f538b43d",
          6300 => x"fefc1153",
          6301 => x"ff840551",
          6302 => x"feece53f",
          6303 => x"828cdc08",
          6304 => x"802efcde",
          6305 => x"38b43dfe",
          6306 => x"f81153ff",
          6307 => x"840551fe",
          6308 => x"ecce3f82",
          6309 => x"8cdc0880",
          6310 => x"2efcc738",
          6311 => x"8284fc51",
          6312 => x"fee4e43f",
          6313 => x"635a7963",
          6314 => x"27a83861",
          6315 => x"70337b33",
          6316 => x"5e5a5b78",
          6317 => x"7c2e9238",
          6318 => x"78557a54",
          6319 => x"79335379",
          6320 => x"5282858c",
          6321 => x"51feeaa3",
          6322 => x"3f811a62",
          6323 => x"8105435a",
          6324 => x"d5398285",
          6325 => x"a45182bd",
          6326 => x"39b43dff",
          6327 => x"801153ff",
          6328 => x"840551fe",
          6329 => x"ebfa3f82",
          6330 => x"8cdc0880",
          6331 => x"df388288",
          6332 => x"a0335978",
          6333 => x"802e8938",
          6334 => x"8287d808",
          6335 => x"4480cd39",
          6336 => x"8288a133",
          6337 => x"5978802e",
          6338 => x"88388287",
          6339 => x"e00844bc",
          6340 => x"398288a2",
          6341 => x"33597880",
          6342 => x"2e883882",
          6343 => x"87e80844",
          6344 => x"ab398288",
          6345 => x"a3335978",
          6346 => x"802e8838",
          6347 => x"8287f008",
          6348 => x"449a3982",
          6349 => x"889e3359",
          6350 => x"78802e88",
          6351 => x"388287f8",
          6352 => x"08448939",
          6353 => x"82888808",
          6354 => x"fc800544",
          6355 => x"b43dfefc",
          6356 => x"1153ff84",
          6357 => x"0551feeb",
          6358 => x"873f828c",
          6359 => x"dc0880de",
          6360 => x"388288a0",
          6361 => x"33597880",
          6362 => x"2e893882",
          6363 => x"87dc0843",
          6364 => x"80cc3982",
          6365 => x"88a13359",
          6366 => x"78802e88",
          6367 => x"388287e4",
          6368 => x"0843bb39",
          6369 => x"8288a233",
          6370 => x"5978802e",
          6371 => x"88388287",
          6372 => x"ec0843aa",
          6373 => x"398288a3",
          6374 => x"33597880",
          6375 => x"2e883882",
          6376 => x"87f40843",
          6377 => x"99398288",
          6378 => x"9e335978",
          6379 => x"802e8838",
          6380 => x"8287fc08",
          6381 => x"43883982",
          6382 => x"88880888",
          6383 => x"0543b43d",
          6384 => x"fef81153",
          6385 => x"ff840551",
          6386 => x"feea953f",
          6387 => x"828cdc08",
          6388 => x"802ea738",
          6389 => x"80625c5c",
          6390 => x"7a882e83",
          6391 => x"38815c7a",
          6392 => x"90327030",
          6393 => x"7072079f",
          6394 => x"2a707f06",
          6395 => x"51515a5a",
          6396 => x"78802e88",
          6397 => x"387aa02e",
          6398 => x"83388842",
          6399 => x"8285a851",
          6400 => x"fee2843f",
          6401 => x"a0556354",
          6402 => x"61536252",
          6403 => x"6351f291",
          6404 => x"3f8285b8",
          6405 => x"51fee1ef",
          6406 => x"3ff9c739",
          6407 => x"b43dff80",
          6408 => x"1153ff84",
          6409 => x"0551fee9",
          6410 => x"b73f828c",
          6411 => x"dc08802e",
          6412 => x"f9b038b4",
          6413 => x"3dfefc11",
          6414 => x"53ff8405",
          6415 => x"51fee9a0",
          6416 => x"3f828cdc",
          6417 => x"08802ea5",
          6418 => x"38635902",
          6419 => x"80cb0533",
          6420 => x"79346381",
          6421 => x"0544b43d",
          6422 => x"fefc1153",
          6423 => x"ff840551",
          6424 => x"fee8fd3f",
          6425 => x"828cdc08",
          6426 => x"e038f8f6",
          6427 => x"39637033",
          6428 => x"54528285",
          6429 => x"c451fee6",
          6430 => x"f23f80f8",
          6431 => x"527951fe",
          6432 => x"e7c33f79",
          6433 => x"45793359",
          6434 => x"78ae2ef8",
          6435 => x"d5389f79",
          6436 => x"27a038b4",
          6437 => x"3dfefc11",
          6438 => x"53ff8405",
          6439 => x"51fee8c0",
          6440 => x"3f828cdc",
          6441 => x"08802e91",
          6442 => x"38635902",
          6443 => x"80cb0533",
          6444 => x"79346381",
          6445 => x"0544ffb5",
          6446 => x"398285d0",
          6447 => x"51fee0c7",
          6448 => x"3fffaa39",
          6449 => x"b43dfef4",
          6450 => x"1153ff84",
          6451 => x"0551feea",
          6452 => x"813f828c",
          6453 => x"dc08802e",
          6454 => x"f88838b4",
          6455 => x"3dfef011",
          6456 => x"53ff8405",
          6457 => x"51fee9ea",
          6458 => x"3f828cdc",
          6459 => x"08802ea6",
          6460 => x"38605902",
          6461 => x"be052279",
          6462 => x"7082055b",
          6463 => x"237841b4",
          6464 => x"3dfef011",
          6465 => x"53ff8405",
          6466 => x"51fee9c6",
          6467 => x"3f828cdc",
          6468 => x"08df38f7",
          6469 => x"cd396070",
          6470 => x"22545282",
          6471 => x"85d851fe",
          6472 => x"e5c93f80",
          6473 => x"f8527951",
          6474 => x"fee69a3f",
          6475 => x"79457933",
          6476 => x"5978ae2e",
          6477 => x"f7ac3878",
          6478 => x"9f268738",
          6479 => x"60820541",
          6480 => x"d539b43d",
          6481 => x"fef01153",
          6482 => x"ff840551",
          6483 => x"fee9833f",
          6484 => x"828cdc08",
          6485 => x"802e9238",
          6486 => x"605902be",
          6487 => x"05227970",
          6488 => x"82055b23",
          6489 => x"7841ffae",
          6490 => x"398285d0",
          6491 => x"51fedf97",
          6492 => x"3fffa339",
          6493 => x"b43dfef4",
          6494 => x"1153ff84",
          6495 => x"0551fee8",
          6496 => x"d13f828c",
          6497 => x"dc08802e",
          6498 => x"f6d838b4",
          6499 => x"3dfef011",
          6500 => x"53ff8405",
          6501 => x"51fee8ba",
          6502 => x"3f828cdc",
          6503 => x"08802ea1",
          6504 => x"38606071",
          6505 => x"0c596084",
          6506 => x"0541b43d",
          6507 => x"fef01153",
          6508 => x"ff840551",
          6509 => x"fee89b3f",
          6510 => x"828cdc08",
          6511 => x"e438f6a2",
          6512 => x"39607008",
          6513 => x"54528285",
          6514 => x"e451fee4",
          6515 => x"9e3f80f8",
          6516 => x"527951fe",
          6517 => x"e4ef3f79",
          6518 => x"45793359",
          6519 => x"78ae2ef6",
          6520 => x"81389f79",
          6521 => x"279c38b4",
          6522 => x"3dfef011",
          6523 => x"53ff8405",
          6524 => x"51fee7de",
          6525 => x"3f828cdc",
          6526 => x"08802e8d",
          6527 => x"38606071",
          6528 => x"0c596084",
          6529 => x"0541ffb9",
          6530 => x"398285d0",
          6531 => x"51feddf7",
          6532 => x"3fffae39",
          6533 => x"b43dff80",
          6534 => x"1153ff84",
          6535 => x"0551fee5",
          6536 => x"bf3f828c",
          6537 => x"dc08802e",
          6538 => x"f5b83863",
          6539 => x"528285f0",
          6540 => x"51fee3b7",
          6541 => x"3f635978",
          6542 => x"04b43dff",
          6543 => x"801153ff",
          6544 => x"840551fe",
          6545 => x"e59a3f82",
          6546 => x"8cdc0880",
          6547 => x"2ef59338",
          6548 => x"63528286",
          6549 => x"8c51fee3",
          6550 => x"923f6359",
          6551 => x"782d828c",
          6552 => x"dc08802e",
          6553 => x"f4fc3882",
          6554 => x"8cdc0852",
          6555 => x"8286a851",
          6556 => x"fee2f83f",
          6557 => x"f4ec3982",
          6558 => x"86c451fe",
          6559 => x"dd893ffe",
          6560 => x"bdb93ff4",
          6561 => x"dd398286",
          6562 => x"e051fedc",
          6563 => x"fa3f8059",
          6564 => x"ffa539fe",
          6565 => x"d38c3ff4",
          6566 => x"c9397945",
          6567 => x"79335978",
          6568 => x"802ef4be",
          6569 => x"387d7d06",
          6570 => x"5978802e",
          6571 => x"81d338b4",
          6572 => x"3dff8405",
          6573 => x"51fec68b",
          6574 => x"3f828cdc",
          6575 => x"085c815b",
          6576 => x"7a822eb2",
          6577 => x"387a8224",
          6578 => x"89387a81",
          6579 => x"2e8c3880",
          6580 => x"cd397a83",
          6581 => x"2eb03880",
          6582 => x"c5398286",
          6583 => x"f4567b55",
          6584 => x"8286f854",
          6585 => x"80538286",
          6586 => x"fc52b43d",
          6587 => x"ffb00551",
          6588 => x"fee28e3f",
          6589 => x"bb398287",
          6590 => x"9c52b43d",
          6591 => x"ffb00551",
          6592 => x"fee1fe3f",
          6593 => x"ab397b55",
          6594 => x"8286f854",
          6595 => x"80538287",
          6596 => x"8c52b43d",
          6597 => x"ffb00551",
          6598 => x"fee1e63f",
          6599 => x"93397b54",
          6600 => x"80538287",
          6601 => x"9852b43d",
          6602 => x"ffb00551",
          6603 => x"fee1d23f",
          6604 => x"8287d858",
          6605 => x"828da457",
          6606 => x"80566455",
          6607 => x"80548380",
          6608 => x"80538380",
          6609 => x"8052b43d",
          6610 => x"ffb00551",
          6611 => x"eb8a3f82",
          6612 => x"8cdc0882",
          6613 => x"8cdc0809",
          6614 => x"70307072",
          6615 => x"07802551",
          6616 => x"5b5b5f80",
          6617 => x"5a7a8326",
          6618 => x"8338815a",
          6619 => x"787a0659",
          6620 => x"78802e8d",
          6621 => x"38811b70",
          6622 => x"81ff065c",
          6623 => x"597afec0",
          6624 => x"387d8132",
          6625 => x"7d813207",
          6626 => x"59788a38",
          6627 => x"7eff2e09",
          6628 => x"8106f2ce",
          6629 => x"388287a0",
          6630 => x"51fee0cf",
          6631 => x"3ff2c339",
          6632 => x"fc3d0d80",
          6633 => x"0b828da4",
          6634 => x"3487c094",
          6635 => x"8c700854",
          6636 => x"55878480",
          6637 => x"527251fe",
          6638 => x"bba13f82",
          6639 => x"8cdc0890",
          6640 => x"2b750855",
          6641 => x"53878480",
          6642 => x"527351fe",
          6643 => x"bb8d3f72",
          6644 => x"828cdc08",
          6645 => x"07750c87",
          6646 => x"c0949c70",
          6647 => x"08545587",
          6648 => x"84805272",
          6649 => x"51febaf3",
          6650 => x"3f828cdc",
          6651 => x"08902b75",
          6652 => x"08555387",
          6653 => x"84805273",
          6654 => x"51febadf",
          6655 => x"3f72828c",
          6656 => x"dc080775",
          6657 => x"0c8c8083",
          6658 => x"0b87c094",
          6659 => x"840c8c80",
          6660 => x"830b87c0",
          6661 => x"94940cb7",
          6662 => x"ac0b828c",
          6663 => x"f00cbaad",
          6664 => x"0b828cf4",
          6665 => x"0cfecbae",
          6666 => x"3ffed4d7",
          6667 => x"3f8287b0",
          6668 => x"51fed9d3",
          6669 => x"3f8287bc",
          6670 => x"51fed9cb",
          6671 => x"3f81ddc6",
          6672 => x"51fed4ba",
          6673 => x"3f8151ec",
          6674 => x"be3ff0c6",
          6675 => x"3f800400",
          6676 => x"00002255",
          6677 => x"0000225b",
          6678 => x"00002261",
          6679 => x"00002267",
          6680 => x"0000226d",
          6681 => x"00002fd8",
          6682 => x"000030b4",
          6683 => x"00003157",
          6684 => x"00003197",
          6685 => x"000031ba",
          6686 => x"00003247",
          6687 => x"00002ead",
          6688 => x"00002ead",
          6689 => x"00003284",
          6690 => x"000032fa",
          6691 => x"00003385",
          6692 => x"000033ae",
          6693 => x"00006bcc",
          6694 => x"00006b50",
          6695 => x"00006b57",
          6696 => x"00006b5e",
          6697 => x"00006b65",
          6698 => x"00006b6c",
          6699 => x"00006b73",
          6700 => x"00006b7a",
          6701 => x"00006b81",
          6702 => x"00006b88",
          6703 => x"00006b8f",
          6704 => x"00006b96",
          6705 => x"00006b9c",
          6706 => x"00006ba2",
          6707 => x"00006ba8",
          6708 => x"00006bae",
          6709 => x"00006bb4",
          6710 => x"00006bba",
          6711 => x"00006bc0",
          6712 => x"00006bc6",
          6713 => x"25642f25",
          6714 => x"642f2564",
          6715 => x"2025643a",
          6716 => x"25643a25",
          6717 => x"642e2564",
          6718 => x"25640a00",
          6719 => x"536f4320",
          6720 => x"436f6e66",
          6721 => x"69677572",
          6722 => x"6174696f",
          6723 => x"6e000000",
          6724 => x"20286672",
          6725 => x"6f6d2053",
          6726 => x"6f432063",
          6727 => x"6f6e6669",
          6728 => x"67290000",
          6729 => x"3a0a4465",
          6730 => x"76696365",
          6731 => x"7320696d",
          6732 => x"706c656d",
          6733 => x"656e7465",
          6734 => x"643a0a00",
          6735 => x"20202020",
          6736 => x"57422053",
          6737 => x"4452414d",
          6738 => x"20202825",
          6739 => x"3038583a",
          6740 => x"25303858",
          6741 => x"292e0a00",
          6742 => x"20202020",
          6743 => x"53445241",
          6744 => x"4d202020",
          6745 => x"20202825",
          6746 => x"3038583a",
          6747 => x"25303858",
          6748 => x"292e0a00",
          6749 => x"20202020",
          6750 => x"494e534e",
          6751 => x"20425241",
          6752 => x"4d202825",
          6753 => x"3038583a",
          6754 => x"25303858",
          6755 => x"292e0a00",
          6756 => x"20202020",
          6757 => x"4252414d",
          6758 => x"20202020",
          6759 => x"20202825",
          6760 => x"3038583a",
          6761 => x"25303858",
          6762 => x"292e0a00",
          6763 => x"20202020",
          6764 => x"52414d20",
          6765 => x"20202020",
          6766 => x"20202825",
          6767 => x"3038583a",
          6768 => x"25303858",
          6769 => x"292e0a00",
          6770 => x"20202020",
          6771 => x"53442043",
          6772 => x"41524420",
          6773 => x"20202844",
          6774 => x"65766963",
          6775 => x"6573203d",
          6776 => x"25303264",
          6777 => x"292e0a00",
          6778 => x"20202020",
          6779 => x"54494d45",
          6780 => x"52312020",
          6781 => x"20202854",
          6782 => x"696d6572",
          6783 => x"7320203d",
          6784 => x"25303264",
          6785 => x"292e0a00",
          6786 => x"20202020",
          6787 => x"494e5452",
          6788 => x"20435452",
          6789 => x"4c202843",
          6790 => x"68616e6e",
          6791 => x"656c733d",
          6792 => x"25303264",
          6793 => x"292e0a00",
          6794 => x"20202020",
          6795 => x"57495348",
          6796 => x"424f4e45",
          6797 => x"20425553",
          6798 => x"0a000000",
          6799 => x"20202020",
          6800 => x"57422049",
          6801 => x"32430a00",
          6802 => x"20202020",
          6803 => x"494f4354",
          6804 => x"4c0a0000",
          6805 => x"20202020",
          6806 => x"5053320a",
          6807 => x"00000000",
          6808 => x"20202020",
          6809 => x"5350490a",
          6810 => x"00000000",
          6811 => x"41646472",
          6812 => x"65737365",
          6813 => x"733a0a00",
          6814 => x"20202020",
          6815 => x"43505520",
          6816 => x"52657365",
          6817 => x"74205665",
          6818 => x"63746f72",
          6819 => x"20416464",
          6820 => x"72657373",
          6821 => x"203d2025",
          6822 => x"3038580a",
          6823 => x"00000000",
          6824 => x"20202020",
          6825 => x"43505520",
          6826 => x"4d656d6f",
          6827 => x"72792053",
          6828 => x"74617274",
          6829 => x"20416464",
          6830 => x"72657373",
          6831 => x"203d2025",
          6832 => x"3038580a",
          6833 => x"00000000",
          6834 => x"20202020",
          6835 => x"53746163",
          6836 => x"6b205374",
          6837 => x"61727420",
          6838 => x"41646472",
          6839 => x"65737320",
          6840 => x"20202020",
          6841 => x"203d2025",
          6842 => x"3038580a",
          6843 => x"00000000",
          6844 => x"4d697363",
          6845 => x"3a0a0000",
          6846 => x"20202020",
          6847 => x"5a505520",
          6848 => x"49642020",
          6849 => x"20202020",
          6850 => x"20202020",
          6851 => x"20202020",
          6852 => x"20202020",
          6853 => x"203d2025",
          6854 => x"3034580a",
          6855 => x"00000000",
          6856 => x"20202020",
          6857 => x"53797374",
          6858 => x"656d2043",
          6859 => x"6c6f636b",
          6860 => x"20467265",
          6861 => x"71202020",
          6862 => x"20202020",
          6863 => x"203d2025",
          6864 => x"642e2530",
          6865 => x"34644d48",
          6866 => x"7a0a0000",
          6867 => x"20202020",
          6868 => x"53445241",
          6869 => x"4d20436c",
          6870 => x"6f636b20",
          6871 => x"46726571",
          6872 => x"20202020",
          6873 => x"20202020",
          6874 => x"203d2025",
          6875 => x"642e2530",
          6876 => x"34644d48",
          6877 => x"7a0a0000",
          6878 => x"20202020",
          6879 => x"57697368",
          6880 => x"626f6e65",
          6881 => x"20534452",
          6882 => x"414d2043",
          6883 => x"6c6f636b",
          6884 => x"20467265",
          6885 => x"713d2025",
          6886 => x"642e2530",
          6887 => x"34644d48",
          6888 => x"7a0a0000",
          6889 => x"536d616c",
          6890 => x"6c000000",
          6891 => x"4d656469",
          6892 => x"756d0000",
          6893 => x"466c6578",
          6894 => x"00000000",
          6895 => x"45564f00",
          6896 => x"45564f6d",
          6897 => x"696e0000",
          6898 => x"556e6b6e",
          6899 => x"6f776e00",
          6900 => x"68697374",
          6901 => x"6f72792e",
          6902 => x"74787400",
          6903 => x"68697374",
          6904 => x"6f727900",
          6905 => x"68697374",
          6906 => x"00000000",
          6907 => x"21000000",
          6908 => x"25303464",
          6909 => x"20202573",
          6910 => x"0a000000",
          6911 => x"4661696c",
          6912 => x"65642074",
          6913 => x"6f207265",
          6914 => x"73657420",
          6915 => x"74686520",
          6916 => x"68697374",
          6917 => x"6f727920",
          6918 => x"66696c65",
          6919 => x"20746f20",
          6920 => x"454f462e",
          6921 => x"0a000000",
          6922 => x"43616e6e",
          6923 => x"6f74206f",
          6924 => x"70656e2f",
          6925 => x"63726561",
          6926 => x"74652068",
          6927 => x"6973746f",
          6928 => x"72792066",
          6929 => x"696c652c",
          6930 => x"20646973",
          6931 => x"61626c69",
          6932 => x"6e672e0a",
          6933 => x"00000000",
          6934 => x"00007d04",
          6935 => x"01000000",
          6936 => x"00000001",
          6937 => x"00007d00",
          6938 => x"01000000",
          6939 => x"00000002",
          6940 => x"00007cfc",
          6941 => x"04000000",
          6942 => x"00000003",
          6943 => x"00007cf8",
          6944 => x"04000000",
          6945 => x"00000004",
          6946 => x"00007cf4",
          6947 => x"04000000",
          6948 => x"00000005",
          6949 => x"00007cf0",
          6950 => x"04000000",
          6951 => x"00000006",
          6952 => x"00007cec",
          6953 => x"04000000",
          6954 => x"00000007",
          6955 => x"00007ce8",
          6956 => x"03000000",
          6957 => x"00000008",
          6958 => x"00007ce4",
          6959 => x"03000000",
          6960 => x"00000009",
          6961 => x"00007ce0",
          6962 => x"03000000",
          6963 => x"0000000a",
          6964 => x"00007cdc",
          6965 => x"03000000",
          6966 => x"0000000b",
          6967 => x"1b5b4400",
          6968 => x"1b5b4300",
          6969 => x"1b5b4200",
          6970 => x"1b5b4100",
          6971 => x"1b5b367e",
          6972 => x"1b5b357e",
          6973 => x"1b5b347e",
          6974 => x"1b5b337e",
          6975 => x"1b5b317e",
          6976 => x"0d000000",
          6977 => x"08000000",
          6978 => x"53440000",
          6979 => x"222a2b2c",
          6980 => x"3a3b3c3d",
          6981 => x"3e3f5b5d",
          6982 => x"7c7f0000",
          6983 => x"46415400",
          6984 => x"46415433",
          6985 => x"32000000",
          6986 => x"ebfe904d",
          6987 => x"53444f53",
          6988 => x"352e3000",
          6989 => x"4e4f204e",
          6990 => x"414d4520",
          6991 => x"20202046",
          6992 => x"41543332",
          6993 => x"20202000",
          6994 => x"4e4f204e",
          6995 => x"414d4520",
          6996 => x"20202046",
          6997 => x"41542020",
          6998 => x"20202000",
          6999 => x"00007d08",
          7000 => x"00000000",
          7001 => x"00000000",
          7002 => x"00000000",
          7003 => x"809a4541",
          7004 => x"8e418f80",
          7005 => x"45454549",
          7006 => x"49498e8f",
          7007 => x"9092924f",
          7008 => x"994f5555",
          7009 => x"59999a9b",
          7010 => x"9c9d9e9f",
          7011 => x"41494f55",
          7012 => x"a5a5a6a7",
          7013 => x"a8a9aaab",
          7014 => x"acadaeaf",
          7015 => x"b0b1b2b3",
          7016 => x"b4b5b6b7",
          7017 => x"b8b9babb",
          7018 => x"bcbdbebf",
          7019 => x"c0c1c2c3",
          7020 => x"c4c5c6c7",
          7021 => x"c8c9cacb",
          7022 => x"cccdcecf",
          7023 => x"d0d1d2d3",
          7024 => x"d4d5d6d7",
          7025 => x"d8d9dadb",
          7026 => x"dcdddedf",
          7027 => x"e0e1e2e3",
          7028 => x"e4e5e6e7",
          7029 => x"e8e9eaeb",
          7030 => x"ecedeeef",
          7031 => x"f0f1f2f3",
          7032 => x"f4f5f6f7",
          7033 => x"f8f9fafb",
          7034 => x"fcfdfeff",
          7035 => x"2b2e2c3b",
          7036 => x"3d5b5d2f",
          7037 => x"5c222a3a",
          7038 => x"3c3e3f7c",
          7039 => x"7f000000",
          7040 => x"00010004",
          7041 => x"00100040",
          7042 => x"01000200",
          7043 => x"00000000",
          7044 => x"00010002",
          7045 => x"00040008",
          7046 => x"00100020",
          7047 => x"00000000",
          7048 => x"64696e69",
          7049 => x"74000000",
          7050 => x"64696f63",
          7051 => x"746c0000",
          7052 => x"66696e69",
          7053 => x"74000000",
          7054 => x"666c6f61",
          7055 => x"64000000",
          7056 => x"66657865",
          7057 => x"63000000",
          7058 => x"6d636c65",
          7059 => x"61720000",
          7060 => x"6d636f70",
          7061 => x"79000000",
          7062 => x"6d646966",
          7063 => x"66000000",
          7064 => x"6d64756d",
          7065 => x"70000000",
          7066 => x"6d656200",
          7067 => x"6d656800",
          7068 => x"6d657700",
          7069 => x"68696400",
          7070 => x"68696500",
          7071 => x"68666400",
          7072 => x"68666500",
          7073 => x"63616c6c",
          7074 => x"00000000",
          7075 => x"6a6d7000",
          7076 => x"72657374",
          7077 => x"61727400",
          7078 => x"72657365",
          7079 => x"74000000",
          7080 => x"696e666f",
          7081 => x"00000000",
          7082 => x"74657374",
          7083 => x"00000000",
          7084 => x"74626173",
          7085 => x"69630000",
          7086 => x"6d626173",
          7087 => x"69630000",
          7088 => x"6b696c6f",
          7089 => x"00000000",
          7090 => x"4469736b",
          7091 => x"20457272",
          7092 => x"6f720a00",
          7093 => x"496e7465",
          7094 => x"726e616c",
          7095 => x"20657272",
          7096 => x"6f722e0a",
          7097 => x"00000000",
          7098 => x"4469736b",
          7099 => x"206e6f74",
          7100 => x"20726561",
          7101 => x"64792e0a",
          7102 => x"00000000",
          7103 => x"4e6f2066",
          7104 => x"696c6520",
          7105 => x"666f756e",
          7106 => x"642e0a00",
          7107 => x"4e6f2070",
          7108 => x"61746820",
          7109 => x"666f756e",
          7110 => x"642e0a00",
          7111 => x"496e7661",
          7112 => x"6c696420",
          7113 => x"66696c65",
          7114 => x"6e616d65",
          7115 => x"2e0a0000",
          7116 => x"41636365",
          7117 => x"73732064",
          7118 => x"656e6965",
          7119 => x"642e0a00",
          7120 => x"46696c65",
          7121 => x"20616c72",
          7122 => x"65616479",
          7123 => x"20657869",
          7124 => x"7374732e",
          7125 => x"0a000000",
          7126 => x"46696c65",
          7127 => x"2068616e",
          7128 => x"646c6520",
          7129 => x"696e7661",
          7130 => x"6c69642e",
          7131 => x"0a000000",
          7132 => x"53442069",
          7133 => x"73207772",
          7134 => x"69746520",
          7135 => x"70726f74",
          7136 => x"65637465",
          7137 => x"642e0a00",
          7138 => x"44726976",
          7139 => x"65206e75",
          7140 => x"6d626572",
          7141 => x"20697320",
          7142 => x"696e7661",
          7143 => x"6c69642e",
          7144 => x"0a000000",
          7145 => x"4469736b",
          7146 => x"206e6f74",
          7147 => x"20656e61",
          7148 => x"626c6564",
          7149 => x"2e0a0000",
          7150 => x"4e6f2063",
          7151 => x"6f6d7061",
          7152 => x"7469626c",
          7153 => x"65206669",
          7154 => x"6c657379",
          7155 => x"7374656d",
          7156 => x"20666f75",
          7157 => x"6e64206f",
          7158 => x"6e206469",
          7159 => x"736b2e0a",
          7160 => x"00000000",
          7161 => x"466f726d",
          7162 => x"61742061",
          7163 => x"626f7274",
          7164 => x"65642e0a",
          7165 => x"00000000",
          7166 => x"54696d65",
          7167 => x"6f75742c",
          7168 => x"206f7065",
          7169 => x"72617469",
          7170 => x"6f6e2063",
          7171 => x"616e6365",
          7172 => x"6c6c6564",
          7173 => x"2e0a0000",
          7174 => x"46696c65",
          7175 => x"20697320",
          7176 => x"6c6f636b",
          7177 => x"65642e0a",
          7178 => x"00000000",
          7179 => x"496e7375",
          7180 => x"66666963",
          7181 => x"69656e74",
          7182 => x"206d656d",
          7183 => x"6f72792e",
          7184 => x"0a000000",
          7185 => x"546f6f20",
          7186 => x"6d616e79",
          7187 => x"206f7065",
          7188 => x"6e206669",
          7189 => x"6c65732e",
          7190 => x"0a000000",
          7191 => x"50617261",
          7192 => x"6d657465",
          7193 => x"72732069",
          7194 => x"6e636f72",
          7195 => x"72656374",
          7196 => x"2e0a0000",
          7197 => x"53756363",
          7198 => x"6573732e",
          7199 => x"0a000000",
          7200 => x"556e6b6e",
          7201 => x"6f776e20",
          7202 => x"6572726f",
          7203 => x"722e0a00",
          7204 => x"0a256c75",
          7205 => x"20627974",
          7206 => x"65732025",
          7207 => x"73206174",
          7208 => x"20256c75",
          7209 => x"20627974",
          7210 => x"65732f73",
          7211 => x"65632e0a",
          7212 => x"00000000",
          7213 => x"72656164",
          7214 => x"00000000",
          7215 => x"25303858",
          7216 => x"00000000",
          7217 => x"3a202000",
          7218 => x"25303458",
          7219 => x"00000000",
          7220 => x"20202020",
          7221 => x"20202020",
          7222 => x"00000000",
          7223 => x"25303258",
          7224 => x"00000000",
          7225 => x"20200000",
          7226 => x"207c0000",
          7227 => x"7c0d0a00",
          7228 => x"7a4f5300",
          7229 => x"0a2a2a20",
          7230 => x"25732028",
          7231 => x"00000000",
          7232 => x"31372f30",
          7233 => x"342f3230",
          7234 => x"32300000",
          7235 => x"76312e30",
          7236 => x"31000000",
          7237 => x"205a5055",
          7238 => x"2c207265",
          7239 => x"76202530",
          7240 => x"32782920",
          7241 => x"25732025",
          7242 => x"73202a2a",
          7243 => x"0a0a0000",
          7244 => x"5a505520",
          7245 => x"496e7465",
          7246 => x"72727570",
          7247 => x"74204861",
          7248 => x"6e646c65",
          7249 => x"720a0000",
          7250 => x"54696d65",
          7251 => x"7220696e",
          7252 => x"74657272",
          7253 => x"7570740a",
          7254 => x"00000000",
          7255 => x"50533220",
          7256 => x"696e7465",
          7257 => x"72727570",
          7258 => x"740a0000",
          7259 => x"494f4354",
          7260 => x"4c205244",
          7261 => x"20696e74",
          7262 => x"65727275",
          7263 => x"70740a00",
          7264 => x"494f4354",
          7265 => x"4c205752",
          7266 => x"20696e74",
          7267 => x"65727275",
          7268 => x"70740a00",
          7269 => x"55415254",
          7270 => x"30205258",
          7271 => x"20696e74",
          7272 => x"65727275",
          7273 => x"70740a00",
          7274 => x"55415254",
          7275 => x"30205458",
          7276 => x"20696e74",
          7277 => x"65727275",
          7278 => x"70740a00",
          7279 => x"55415254",
          7280 => x"31205258",
          7281 => x"20696e74",
          7282 => x"65727275",
          7283 => x"70740a00",
          7284 => x"55415254",
          7285 => x"31205458",
          7286 => x"20696e74",
          7287 => x"65727275",
          7288 => x"70740a00",
          7289 => x"53657474",
          7290 => x"696e6720",
          7291 => x"75702074",
          7292 => x"696d6572",
          7293 => x"2e2e2e0a",
          7294 => x"00000000",
          7295 => x"456e6162",
          7296 => x"6c696e67",
          7297 => x"2074696d",
          7298 => x"65722e2e",
          7299 => x"2e0a0000",
          7300 => x"6175746f",
          7301 => x"65786563",
          7302 => x"2e626174",
          7303 => x"00000000",
          7304 => x"303a0000",
          7305 => x"4661696c",
          7306 => x"65642074",
          7307 => x"6f20696e",
          7308 => x"69746961",
          7309 => x"6c697365",
          7310 => x"20736420",
          7311 => x"63617264",
          7312 => x"20302c20",
          7313 => x"706c6561",
          7314 => x"73652069",
          7315 => x"6e697420",
          7316 => x"6d616e75",
          7317 => x"616c6c79",
          7318 => x"2e0a0000",
          7319 => x"2a200000",
          7320 => x"436c6561",
          7321 => x"72696e67",
          7322 => x"2e2e2e2e",
          7323 => x"00000000",
          7324 => x"436f7079",
          7325 => x"696e672e",
          7326 => x"2e2e0000",
          7327 => x"436f6d70",
          7328 => x"6172696e",
          7329 => x"672e2e2e",
          7330 => x"00000000",
          7331 => x"2530386c",
          7332 => x"78282530",
          7333 => x"3878292d",
          7334 => x"3e253038",
          7335 => x"6c782825",
          7336 => x"30387829",
          7337 => x"0a000000",
          7338 => x"44756d70",
          7339 => x"204d656d",
          7340 => x"6f72790a",
          7341 => x"00000000",
          7342 => x"0a436f6d",
          7343 => x"706c6574",
          7344 => x"652e0a00",
          7345 => x"25303858",
          7346 => x"20253032",
          7347 => x"582d0000",
          7348 => x"3f3f3f0a",
          7349 => x"00000000",
          7350 => x"25303858",
          7351 => x"20253034",
          7352 => x"582d0000",
          7353 => x"25303858",
          7354 => x"20253038",
          7355 => x"582d0000",
          7356 => x"45786563",
          7357 => x"7574696e",
          7358 => x"6720636f",
          7359 => x"64652040",
          7360 => x"20253038",
          7361 => x"78202e2e",
          7362 => x"2e0a0000",
          7363 => x"43616c6c",
          7364 => x"696e6720",
          7365 => x"636f6465",
          7366 => x"20402025",
          7367 => x"30387820",
          7368 => x"2e2e2e0a",
          7369 => x"00000000",
          7370 => x"43616c6c",
          7371 => x"20726574",
          7372 => x"75726e65",
          7373 => x"6420636f",
          7374 => x"64652028",
          7375 => x"2564292e",
          7376 => x"0a000000",
          7377 => x"52657374",
          7378 => x"61727469",
          7379 => x"6e672061",
          7380 => x"70706c69",
          7381 => x"63617469",
          7382 => x"6f6e2e2e",
          7383 => x"2e0a0000",
          7384 => x"436f6c64",
          7385 => x"20726562",
          7386 => x"6f6f7469",
          7387 => x"6e672e2e",
          7388 => x"2e0a0000",
          7389 => x"5a505500",
          7390 => x"62696e00",
          7391 => x"25643a5c",
          7392 => x"25735c25",
          7393 => x"732e2573",
          7394 => x"00000000",
          7395 => x"25643a5c",
          7396 => x"25735c25",
          7397 => x"73000000",
          7398 => x"25643a5c",
          7399 => x"25730000",
          7400 => x"42616420",
          7401 => x"636f6d6d",
          7402 => x"616e642e",
          7403 => x"0a000000",
          7404 => x"52756e6e",
          7405 => x"696e672e",
          7406 => x"2e2e0a00",
          7407 => x"456e6162",
          7408 => x"6c696e67",
          7409 => x"20696e74",
          7410 => x"65727275",
          7411 => x"7074732e",
          7412 => x"2e2e0a00",
          7413 => x"00000000",
          7414 => x"00000000",
          7415 => x"00007fff",
          7416 => x"00000000",
          7417 => x"00007fff",
          7418 => x"00010000",
          7419 => x"00007fff",
          7420 => x"00010000",
          7421 => x"00810000",
          7422 => x"01000000",
          7423 => x"017fffff",
          7424 => x"00000000",
          7425 => x"00000000",
          7426 => x"00007800",
          7427 => x"00000000",
          7428 => x"05f5e100",
          7429 => x"05f5e100",
          7430 => x"05f5e100",
          7431 => x"00000000",
          7432 => x"01010101",
          7433 => x"01010101",
          7434 => x"01011001",
          7435 => x"01000000",
          7436 => x"00000000",
          7437 => x"00000002",
          7438 => x"00000000",
          7439 => x"00008434",
          7440 => x"00008434",
          7441 => x"00008434",
          7442 => x"00008434",
          7443 => x"00007bd0",
          7444 => x"00000000",
          7445 => x"00000000",
          7446 => x"00000000",
          7447 => x"00000000",
          7448 => x"00000000",
          7449 => x"00000000",
          7450 => x"00000000",
          7451 => x"00000000",
          7452 => x"00000000",
          7453 => x"00000000",
          7454 => x"00000000",
          7455 => x"00000000",
          7456 => x"00000000",
          7457 => x"00000000",
          7458 => x"00000000",
          7459 => x"00000000",
          7460 => x"00000000",
          7461 => x"00000000",
          7462 => x"00000000",
          7463 => x"00000000",
          7464 => x"00000000",
          7465 => x"00000000",
          7466 => x"00000000",
          7467 => x"00007bdc",
          7468 => x"01000000",
          7469 => x"00007be4",
          7470 => x"01000000",
          7471 => x"00007bec",
          7472 => x"02000000",
          7473 => x"01000000",
          7474 => x"00000000",
          7475 => x"00007e20",
          7476 => x"01020100",
          7477 => x"00000000",
          7478 => x"00000000",
          7479 => x"00007e28",
          7480 => x"01040100",
          7481 => x"00000000",
          7482 => x"00000000",
          7483 => x"00007e30",
          7484 => x"01140300",
          7485 => x"00000000",
          7486 => x"00000000",
          7487 => x"00007e38",
          7488 => x"012b0300",
          7489 => x"00000000",
          7490 => x"00000000",
          7491 => x"00007e40",
          7492 => x"01300300",
          7493 => x"00000000",
          7494 => x"00000000",
          7495 => x"00007e48",
          7496 => x"013c0400",
          7497 => x"00000000",
          7498 => x"00000000",
          7499 => x"00007e50",
          7500 => x"013d0400",
          7501 => x"00000000",
          7502 => x"00000000",
          7503 => x"00007e58",
          7504 => x"013f0400",
          7505 => x"00000000",
          7506 => x"00000000",
          7507 => x"00007e60",
          7508 => x"01400400",
          7509 => x"00000000",
          7510 => x"00000000",
          7511 => x"00007e68",
          7512 => x"01410400",
          7513 => x"00000000",
          7514 => x"00000000",
          7515 => x"00007e6c",
          7516 => x"01420400",
          7517 => x"00000000",
          7518 => x"00000000",
          7519 => x"00007e70",
          7520 => x"01430400",
          7521 => x"00000000",
          7522 => x"00000000",
          7523 => x"00007e74",
          7524 => x"01500500",
          7525 => x"00000000",
          7526 => x"00000000",
          7527 => x"00007e78",
          7528 => x"01510500",
          7529 => x"00000000",
          7530 => x"00000000",
          7531 => x"00007e7c",
          7532 => x"01540500",
          7533 => x"00000000",
          7534 => x"00000000",
          7535 => x"00007e80",
          7536 => x"01550500",
          7537 => x"00000000",
          7538 => x"00000000",
          7539 => x"00007e84",
          7540 => x"01790700",
          7541 => x"00000000",
          7542 => x"00000000",
          7543 => x"00007e8c",
          7544 => x"01780700",
          7545 => x"00000000",
          7546 => x"00000000",
          7547 => x"00007e90",
          7548 => x"01820800",
          7549 => x"00000000",
          7550 => x"00000000",
          7551 => x"00007e98",
          7552 => x"01830800",
          7553 => x"00000000",
          7554 => x"00000000",
          7555 => x"00007ea0",
          7556 => x"01850800",
          7557 => x"00000000",
          7558 => x"00000000",
          7559 => x"00007ea8",
          7560 => x"01870800",
          7561 => x"00000000",
          7562 => x"00000000",
          7563 => x"00007eb0",
          7564 => x"018c0900",
          7565 => x"00000000",
          7566 => x"00000000",
          7567 => x"00007eb8",
          7568 => x"018d0900",
          7569 => x"00000000",
          7570 => x"00000000",
          7571 => x"00007ec0",
          7572 => x"018e0900",
          7573 => x"00000000",
          7574 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

