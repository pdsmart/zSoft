-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"93",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"e0",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"e8",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"eb",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"ed",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"d8",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"2d",
           407 => x"08",
           408 => x"04",
           409 => x"0c",
           410 => x"2d",
           411 => x"08",
           412 => x"04",
           413 => x"0c",
           414 => x"2d",
           415 => x"08",
           416 => x"04",
           417 => x"0c",
           418 => x"2d",
           419 => x"08",
           420 => x"04",
           421 => x"0c",
           422 => x"2d",
           423 => x"08",
           424 => x"04",
           425 => x"0c",
           426 => x"2d",
           427 => x"08",
           428 => x"04",
           429 => x"0c",
           430 => x"2d",
           431 => x"08",
           432 => x"04",
           433 => x"0c",
           434 => x"2d",
           435 => x"08",
           436 => x"04",
           437 => x"0c",
           438 => x"2d",
           439 => x"08",
           440 => x"04",
           441 => x"0c",
           442 => x"2d",
           443 => x"08",
           444 => x"04",
           445 => x"0c",
           446 => x"82",
           447 => x"82",
           448 => x"82",
           449 => x"ba",
           450 => x"87",
           451 => x"a0",
           452 => x"87",
           453 => x"fd",
           454 => x"d8",
           455 => x"90",
           456 => x"d8",
           457 => x"97",
           458 => x"d8",
           459 => x"90",
           460 => x"d8",
           461 => x"88",
           462 => x"d8",
           463 => x"90",
           464 => x"d8",
           465 => x"fc",
           466 => x"d8",
           467 => x"90",
           468 => x"d8",
           469 => x"f9",
           470 => x"d8",
           471 => x"90",
           472 => x"d8",
           473 => x"97",
           474 => x"d8",
           475 => x"90",
           476 => x"d8",
           477 => x"f7",
           478 => x"d8",
           479 => x"90",
           480 => x"d8",
           481 => x"ea",
           482 => x"d8",
           483 => x"90",
           484 => x"d8",
           485 => x"b6",
           486 => x"d8",
           487 => x"90",
           488 => x"d8",
           489 => x"d5",
           490 => x"d8",
           491 => x"90",
           492 => x"d8",
           493 => x"f4",
           494 => x"d8",
           495 => x"90",
           496 => x"d8",
           497 => x"de",
           498 => x"d8",
           499 => x"90",
           500 => x"d8",
           501 => x"c4",
           502 => x"d8",
           503 => x"90",
           504 => x"d8",
           505 => x"b2",
           506 => x"d8",
           507 => x"90",
           508 => x"d8",
           509 => x"f8",
           510 => x"d8",
           511 => x"90",
           512 => x"d8",
           513 => x"b2",
           514 => x"d8",
           515 => x"90",
           516 => x"d8",
           517 => x"b3",
           518 => x"d8",
           519 => x"90",
           520 => x"d8",
           521 => x"e8",
           522 => x"d8",
           523 => x"90",
           524 => x"d8",
           525 => x"c1",
           526 => x"d8",
           527 => x"90",
           528 => x"d8",
           529 => x"ec",
           530 => x"d8",
           531 => x"90",
           532 => x"d8",
           533 => x"cf",
           534 => x"d8",
           535 => x"90",
           536 => x"d8",
           537 => x"a4",
           538 => x"d8",
           539 => x"90",
           540 => x"d8",
           541 => x"ae",
           542 => x"d8",
           543 => x"90",
           544 => x"d8",
           545 => x"f0",
           546 => x"d8",
           547 => x"90",
           548 => x"d8",
           549 => x"b6",
           550 => x"d8",
           551 => x"90",
           552 => x"d8",
           553 => x"dc",
           554 => x"d8",
           555 => x"90",
           556 => x"d8",
           557 => x"91",
           558 => x"d8",
           559 => x"90",
           560 => x"d8",
           561 => x"fd",
           562 => x"d8",
           563 => x"90",
           564 => x"d8",
           565 => x"f2",
           566 => x"d8",
           567 => x"90",
           568 => x"d8",
           569 => x"dc",
           570 => x"d8",
           571 => x"90",
           572 => x"d8",
           573 => x"c0",
           574 => x"d8",
           575 => x"90",
           576 => x"d8",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"82",
           582 => x"82",
           583 => x"82",
           584 => x"bd",
           585 => x"87",
           586 => x"a0",
           587 => x"87",
           588 => x"f4",
           589 => x"d8",
           590 => x"90",
           591 => x"00",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"00",
           601 => x"ff",
           602 => x"06",
           603 => x"83",
           604 => x"10",
           605 => x"fc",
           606 => x"51",
           607 => x"80",
           608 => x"ff",
           609 => x"06",
           610 => x"52",
           611 => x"0a",
           612 => x"38",
           613 => x"51",
           614 => x"cc",
           615 => x"88",
           616 => x"80",
           617 => x"05",
           618 => x"0b",
           619 => x"04",
           620 => x"b7",
           621 => x"82",
           622 => x"02",
           623 => x"0c",
           624 => x"82",
           625 => x"88",
           626 => x"87",
           627 => x"05",
           628 => x"d8",
           629 => x"08",
           630 => x"82",
           631 => x"fc",
           632 => x"05",
           633 => x"08",
           634 => x"70",
           635 => x"51",
           636 => x"2e",
           637 => x"39",
           638 => x"08",
           639 => x"ff",
           640 => x"d8",
           641 => x"0c",
           642 => x"08",
           643 => x"82",
           644 => x"88",
           645 => x"70",
           646 => x"0c",
           647 => x"0d",
           648 => x"0c",
           649 => x"d8",
           650 => x"87",
           651 => x"3d",
           652 => x"d8",
           653 => x"08",
           654 => x"08",
           655 => x"82",
           656 => x"8c",
           657 => x"71",
           658 => x"d8",
           659 => x"08",
           660 => x"87",
           661 => x"05",
           662 => x"d8",
           663 => x"08",
           664 => x"72",
           665 => x"d8",
           666 => x"08",
           667 => x"87",
           668 => x"05",
           669 => x"ff",
           670 => x"80",
           671 => x"ff",
           672 => x"87",
           673 => x"05",
           674 => x"87",
           675 => x"84",
           676 => x"87",
           677 => x"82",
           678 => x"02",
           679 => x"0c",
           680 => x"82",
           681 => x"88",
           682 => x"87",
           683 => x"05",
           684 => x"d8",
           685 => x"08",
           686 => x"08",
           687 => x"82",
           688 => x"90",
           689 => x"2e",
           690 => x"82",
           691 => x"90",
           692 => x"05",
           693 => x"08",
           694 => x"82",
           695 => x"90",
           696 => x"05",
           697 => x"08",
           698 => x"82",
           699 => x"90",
           700 => x"2e",
           701 => x"87",
           702 => x"05",
           703 => x"33",
           704 => x"08",
           705 => x"81",
           706 => x"d8",
           707 => x"0c",
           708 => x"08",
           709 => x"52",
           710 => x"34",
           711 => x"08",
           712 => x"81",
           713 => x"d8",
           714 => x"0c",
           715 => x"82",
           716 => x"88",
           717 => x"82",
           718 => x"51",
           719 => x"82",
           720 => x"04",
           721 => x"08",
           722 => x"d8",
           723 => x"0d",
           724 => x"08",
           725 => x"80",
           726 => x"38",
           727 => x"08",
           728 => x"52",
           729 => x"87",
           730 => x"05",
           731 => x"82",
           732 => x"8c",
           733 => x"87",
           734 => x"05",
           735 => x"72",
           736 => x"53",
           737 => x"71",
           738 => x"38",
           739 => x"82",
           740 => x"88",
           741 => x"71",
           742 => x"d8",
           743 => x"08",
           744 => x"87",
           745 => x"05",
           746 => x"ff",
           747 => x"70",
           748 => x"0b",
           749 => x"08",
           750 => x"81",
           751 => x"87",
           752 => x"05",
           753 => x"82",
           754 => x"90",
           755 => x"87",
           756 => x"05",
           757 => x"84",
           758 => x"39",
           759 => x"08",
           760 => x"80",
           761 => x"38",
           762 => x"08",
           763 => x"70",
           764 => x"70",
           765 => x"0b",
           766 => x"08",
           767 => x"80",
           768 => x"87",
           769 => x"05",
           770 => x"82",
           771 => x"8c",
           772 => x"87",
           773 => x"05",
           774 => x"52",
           775 => x"38",
           776 => x"87",
           777 => x"05",
           778 => x"82",
           779 => x"88",
           780 => x"33",
           781 => x"08",
           782 => x"70",
           783 => x"31",
           784 => x"d8",
           785 => x"0c",
           786 => x"52",
           787 => x"80",
           788 => x"d8",
           789 => x"0c",
           790 => x"08",
           791 => x"82",
           792 => x"85",
           793 => x"87",
           794 => x"82",
           795 => x"02",
           796 => x"0c",
           797 => x"82",
           798 => x"88",
           799 => x"87",
           800 => x"05",
           801 => x"d8",
           802 => x"08",
           803 => x"d4",
           804 => x"d8",
           805 => x"08",
           806 => x"87",
           807 => x"05",
           808 => x"d8",
           809 => x"08",
           810 => x"87",
           811 => x"05",
           812 => x"d8",
           813 => x"08",
           814 => x"38",
           815 => x"08",
           816 => x"51",
           817 => x"d8",
           818 => x"08",
           819 => x"71",
           820 => x"d8",
           821 => x"08",
           822 => x"87",
           823 => x"05",
           824 => x"39",
           825 => x"08",
           826 => x"70",
           827 => x"0c",
           828 => x"0d",
           829 => x"0c",
           830 => x"0d",
           831 => x"70",
           832 => x"74",
           833 => x"e3",
           834 => x"75",
           835 => x"a7",
           836 => x"cc",
           837 => x"0c",
           838 => x"54",
           839 => x"74",
           840 => x"a0",
           841 => x"06",
           842 => x"15",
           843 => x"80",
           844 => x"29",
           845 => x"05",
           846 => x"56",
           847 => x"82",
           848 => x"53",
           849 => x"08",
           850 => x"3f",
           851 => x"08",
           852 => x"16",
           853 => x"81",
           854 => x"38",
           855 => x"81",
           856 => x"54",
           857 => x"c9",
           858 => x"73",
           859 => x"0c",
           860 => x"04",
           861 => x"73",
           862 => x"26",
           863 => x"71",
           864 => x"e8",
           865 => x"71",
           866 => x"eb",
           867 => x"80",
           868 => x"b8",
           869 => x"39",
           870 => x"51",
           871 => x"81",
           872 => x"80",
           873 => x"eb",
           874 => x"e4",
           875 => x"80",
           876 => x"39",
           877 => x"51",
           878 => x"81",
           879 => x"80",
           880 => x"ec",
           881 => x"c8",
           882 => x"d4",
           883 => x"39",
           884 => x"51",
           885 => x"ed",
           886 => x"39",
           887 => x"51",
           888 => x"ed",
           889 => x"39",
           890 => x"51",
           891 => x"ed",
           892 => x"39",
           893 => x"51",
           894 => x"ee",
           895 => x"39",
           896 => x"51",
           897 => x"ee",
           898 => x"39",
           899 => x"51",
           900 => x"83",
           901 => x"fb",
           902 => x"79",
           903 => x"87",
           904 => x"38",
           905 => x"87",
           906 => x"91",
           907 => x"52",
           908 => x"cf",
           909 => x"87",
           910 => x"75",
           911 => x"ab",
           912 => x"cc",
           913 => x"53",
           914 => x"ee",
           915 => x"b4",
           916 => x"0d",
           917 => x"0d",
           918 => x"05",
           919 => x"33",
           920 => x"68",
           921 => x"7a",
           922 => x"51",
           923 => x"78",
           924 => x"ff",
           925 => x"81",
           926 => x"07",
           927 => x"06",
           928 => x"56",
           929 => x"38",
           930 => x"52",
           931 => x"52",
           932 => x"83",
           933 => x"cc",
           934 => x"87",
           935 => x"38",
           936 => x"08",
           937 => x"88",
           938 => x"cc",
           939 => x"3d",
           940 => x"84",
           941 => x"52",
           942 => x"92",
           943 => x"87",
           944 => x"82",
           945 => x"90",
           946 => x"74",
           947 => x"38",
           948 => x"19",
           949 => x"39",
           950 => x"05",
           951 => x"a8",
           952 => x"70",
           953 => x"25",
           954 => x"9f",
           955 => x"51",
           956 => x"74",
           957 => x"38",
           958 => x"53",
           959 => x"88",
           960 => x"51",
           961 => x"76",
           962 => x"87",
           963 => x"3d",
           964 => x"3d",
           965 => x"84",
           966 => x"33",
           967 => x"57",
           968 => x"52",
           969 => x"ad",
           970 => x"cc",
           971 => x"75",
           972 => x"38",
           973 => x"98",
           974 => x"60",
           975 => x"82",
           976 => x"7e",
           977 => x"77",
           978 => x"cc",
           979 => x"39",
           980 => x"82",
           981 => x"89",
           982 => x"f3",
           983 => x"61",
           984 => x"05",
           985 => x"33",
           986 => x"68",
           987 => x"5c",
           988 => x"7a",
           989 => x"a0",
           990 => x"3f",
           991 => x"51",
           992 => x"80",
           993 => x"27",
           994 => x"7b",
           995 => x"38",
           996 => x"a4",
           997 => x"39",
           998 => x"72",
           999 => x"38",
          1000 => x"81",
          1001 => x"b2",
          1002 => x"39",
          1003 => x"51",
          1004 => x"82",
          1005 => x"39",
          1006 => x"72",
          1007 => x"38",
          1008 => x"81",
          1009 => x"b2",
          1010 => x"39",
          1011 => x"51",
          1012 => x"84",
          1013 => x"39",
          1014 => x"72",
          1015 => x"38",
          1016 => x"81",
          1017 => x"b2",
          1018 => x"39",
          1019 => x"51",
          1020 => x"81",
          1021 => x"51",
          1022 => x"ff",
          1023 => x"ef",
          1024 => x"9c",
          1025 => x"74",
          1026 => x"38",
          1027 => x"33",
          1028 => x"56",
          1029 => x"83",
          1030 => x"80",
          1031 => x"27",
          1032 => x"53",
          1033 => x"70",
          1034 => x"51",
          1035 => x"2e",
          1036 => x"80",
          1037 => x"38",
          1038 => x"39",
          1039 => x"83",
          1040 => x"55",
          1041 => x"ef",
          1042 => x"d4",
          1043 => x"79",
          1044 => x"a0",
          1045 => x"87",
          1046 => x"2b",
          1047 => x"51",
          1048 => x"2e",
          1049 => x"aa",
          1050 => x"3f",
          1051 => x"08",
          1052 => x"98",
          1053 => x"32",
          1054 => x"9b",
          1055 => x"70",
          1056 => x"75",
          1057 => x"58",
          1058 => x"51",
          1059 => x"24",
          1060 => x"9b",
          1061 => x"06",
          1062 => x"53",
          1063 => x"1e",
          1064 => x"26",
          1065 => x"ff",
          1066 => x"87",
          1067 => x"3d",
          1068 => x"3d",
          1069 => x"05",
          1070 => x"d4",
          1071 => x"dc",
          1072 => x"c0",
          1073 => x"a4",
          1074 => x"dc",
          1075 => x"e8",
          1076 => x"f4",
          1077 => x"a5",
          1078 => x"ef",
          1079 => x"a4",
          1080 => x"2e",
          1081 => x"a9",
          1082 => x"0d",
          1083 => x"0d",
          1084 => x"80",
          1085 => x"b9",
          1086 => x"9b",
          1087 => x"f0",
          1088 => x"83",
          1089 => x"9b",
          1090 => x"81",
          1091 => x"06",
          1092 => x"80",
          1093 => x"81",
          1094 => x"3f",
          1095 => x"51",
          1096 => x"80",
          1097 => x"3f",
          1098 => x"70",
          1099 => x"52",
          1100 => x"92",
          1101 => x"9a",
          1102 => x"f0",
          1103 => x"c7",
          1104 => x"9a",
          1105 => x"83",
          1106 => x"06",
          1107 => x"80",
          1108 => x"81",
          1109 => x"3f",
          1110 => x"51",
          1111 => x"80",
          1112 => x"3f",
          1113 => x"70",
          1114 => x"52",
          1115 => x"92",
          1116 => x"9a",
          1117 => x"f0",
          1118 => x"8b",
          1119 => x"9a",
          1120 => x"85",
          1121 => x"06",
          1122 => x"80",
          1123 => x"81",
          1124 => x"3f",
          1125 => x"51",
          1126 => x"80",
          1127 => x"3f",
          1128 => x"70",
          1129 => x"52",
          1130 => x"92",
          1131 => x"99",
          1132 => x"f1",
          1133 => x"cf",
          1134 => x"99",
          1135 => x"87",
          1136 => x"06",
          1137 => x"80",
          1138 => x"81",
          1139 => x"3f",
          1140 => x"51",
          1141 => x"80",
          1142 => x"3f",
          1143 => x"70",
          1144 => x"52",
          1145 => x"92",
          1146 => x"99",
          1147 => x"f1",
          1148 => x"93",
          1149 => x"99",
          1150 => x"bd",
          1151 => x"0d",
          1152 => x"0d",
          1153 => x"05",
          1154 => x"70",
          1155 => x"80",
          1156 => x"f4",
          1157 => x"0b",
          1158 => x"33",
          1159 => x"38",
          1160 => x"f1",
          1161 => x"9e",
          1162 => x"86",
          1163 => x"87",
          1164 => x"70",
          1165 => x"08",
          1166 => x"82",
          1167 => x"51",
          1168 => x"0b",
          1169 => x"34",
          1170 => x"82",
          1171 => x"73",
          1172 => x"81",
          1173 => x"82",
          1174 => x"74",
          1175 => x"81",
          1176 => x"82",
          1177 => x"80",
          1178 => x"82",
          1179 => x"51",
          1180 => x"91",
          1181 => x"ac",
          1182 => x"8c",
          1183 => x"0b",
          1184 => x"c8",
          1185 => x"82",
          1186 => x"54",
          1187 => x"09",
          1188 => x"38",
          1189 => x"53",
          1190 => x"51",
          1191 => x"80",
          1192 => x"cc",
          1193 => x"0d",
          1194 => x"0d",
          1195 => x"82",
          1196 => x"5f",
          1197 => x"7c",
          1198 => x"b7",
          1199 => x"cc",
          1200 => x"06",
          1201 => x"2e",
          1202 => x"a1",
          1203 => x"98",
          1204 => x"70",
          1205 => x"c2",
          1206 => x"78",
          1207 => x"d8",
          1208 => x"d2",
          1209 => x"cc",
          1210 => x"88",
          1211 => x"9c",
          1212 => x"39",
          1213 => x"5d",
          1214 => x"51",
          1215 => x"96",
          1216 => x"5a",
          1217 => x"79",
          1218 => x"3f",
          1219 => x"84",
          1220 => x"e5",
          1221 => x"cc",
          1222 => x"70",
          1223 => x"59",
          1224 => x"2e",
          1225 => x"78",
          1226 => x"80",
          1227 => x"ab",
          1228 => x"38",
          1229 => x"a4",
          1230 => x"2e",
          1231 => x"78",
          1232 => x"38",
          1233 => x"ff",
          1234 => x"e1",
          1235 => x"2e",
          1236 => x"78",
          1237 => x"ad",
          1238 => x"39",
          1239 => x"84",
          1240 => x"bd",
          1241 => x"78",
          1242 => x"a5",
          1243 => x"2e",
          1244 => x"8e",
          1245 => x"bf",
          1246 => x"38",
          1247 => x"2e",
          1248 => x"8e",
          1249 => x"80",
          1250 => x"88",
          1251 => x"d5",
          1252 => x"78",
          1253 => x"8c",
          1254 => x"80",
          1255 => x"38",
          1256 => x"2e",
          1257 => x"78",
          1258 => x"8b",
          1259 => x"fd",
          1260 => x"d1",
          1261 => x"38",
          1262 => x"2e",
          1263 => x"8d",
          1264 => x"81",
          1265 => x"c6",
          1266 => x"82",
          1267 => x"78",
          1268 => x"8c",
          1269 => x"80",
          1270 => x"f7",
          1271 => x"39",
          1272 => x"2e",
          1273 => x"78",
          1274 => x"8d",
          1275 => x"bd",
          1276 => x"ff",
          1277 => x"ff",
          1278 => x"ab",
          1279 => x"87",
          1280 => x"38",
          1281 => x"51",
          1282 => x"b4",
          1283 => x"11",
          1284 => x"05",
          1285 => x"3f",
          1286 => x"08",
          1287 => x"38",
          1288 => x"83",
          1289 => x"02",
          1290 => x"33",
          1291 => x"cf",
          1292 => x"80",
          1293 => x"82",
          1294 => x"81",
          1295 => x"78",
          1296 => x"f2",
          1297 => x"d8",
          1298 => x"fd",
          1299 => x"f2",
          1300 => x"9d",
          1301 => x"ff",
          1302 => x"ff",
          1303 => x"ab",
          1304 => x"87",
          1305 => x"2e",
          1306 => x"80",
          1307 => x"02",
          1308 => x"33",
          1309 => x"c8",
          1310 => x"cc",
          1311 => x"f3",
          1312 => x"84",
          1313 => x"ff",
          1314 => x"ff",
          1315 => x"aa",
          1316 => x"87",
          1317 => x"2e",
          1318 => x"89",
          1319 => x"38",
          1320 => x"fc",
          1321 => x"84",
          1322 => x"cd",
          1323 => x"cc",
          1324 => x"82",
          1325 => x"43",
          1326 => x"f3",
          1327 => x"51",
          1328 => x"02",
          1329 => x"33",
          1330 => x"63",
          1331 => x"82",
          1332 => x"51",
          1333 => x"3f",
          1334 => x"08",
          1335 => x"81",
          1336 => x"a2",
          1337 => x"5d",
          1338 => x"b4",
          1339 => x"05",
          1340 => x"3f",
          1341 => x"08",
          1342 => x"84",
          1343 => x"90",
          1344 => x"53",
          1345 => x"08",
          1346 => x"f2",
          1347 => x"d1",
          1348 => x"ff",
          1349 => x"8e",
          1350 => x"87",
          1351 => x"3d",
          1352 => x"52",
          1353 => x"3f",
          1354 => x"08",
          1355 => x"84",
          1356 => x"8f",
          1357 => x"87",
          1358 => x"3d",
          1359 => x"52",
          1360 => x"3f",
          1361 => x"58",
          1362 => x"57",
          1363 => x"55",
          1364 => x"08",
          1365 => x"54",
          1366 => x"52",
          1367 => x"b2",
          1368 => x"cc",
          1369 => x"fb",
          1370 => x"87",
          1371 => x"f0",
          1372 => x"84",
          1373 => x"ff",
          1374 => x"ff",
          1375 => x"a8",
          1376 => x"87",
          1377 => x"2e",
          1378 => x"b4",
          1379 => x"11",
          1380 => x"05",
          1381 => x"3f",
          1382 => x"08",
          1383 => x"d8",
          1384 => x"fe",
          1385 => x"ff",
          1386 => x"a8",
          1387 => x"87",
          1388 => x"38",
          1389 => x"08",
          1390 => x"9c",
          1391 => x"3f",
          1392 => x"5a",
          1393 => x"81",
          1394 => x"59",
          1395 => x"84",
          1396 => x"7a",
          1397 => x"38",
          1398 => x"b4",
          1399 => x"11",
          1400 => x"05",
          1401 => x"3f",
          1402 => x"08",
          1403 => x"88",
          1404 => x"fe",
          1405 => x"ff",
          1406 => x"a7",
          1407 => x"87",
          1408 => x"2e",
          1409 => x"b4",
          1410 => x"11",
          1411 => x"05",
          1412 => x"3f",
          1413 => x"08",
          1414 => x"dc",
          1415 => x"ac",
          1416 => x"3f",
          1417 => x"63",
          1418 => x"38",
          1419 => x"70",
          1420 => x"33",
          1421 => x"81",
          1422 => x"39",
          1423 => x"80",
          1424 => x"84",
          1425 => x"b1",
          1426 => x"cc",
          1427 => x"f9",
          1428 => x"3d",
          1429 => x"53",
          1430 => x"51",
          1431 => x"82",
          1432 => x"80",
          1433 => x"38",
          1434 => x"f8",
          1435 => x"84",
          1436 => x"85",
          1437 => x"cc",
          1438 => x"f8",
          1439 => x"f3",
          1440 => x"9c",
          1441 => x"79",
          1442 => x"38",
          1443 => x"7b",
          1444 => x"5b",
          1445 => x"91",
          1446 => x"7a",
          1447 => x"53",
          1448 => x"f3",
          1449 => x"dc",
          1450 => x"62",
          1451 => x"5a",
          1452 => x"f2",
          1453 => x"b9",
          1454 => x"ff",
          1455 => x"ff",
          1456 => x"a6",
          1457 => x"87",
          1458 => x"df",
          1459 => x"b8",
          1460 => x"80",
          1461 => x"82",
          1462 => x"44",
          1463 => x"82",
          1464 => x"59",
          1465 => x"88",
          1466 => x"f8",
          1467 => x"39",
          1468 => x"33",
          1469 => x"2e",
          1470 => x"86",
          1471 => x"ab",
          1472 => x"bb",
          1473 => x"80",
          1474 => x"82",
          1475 => x"44",
          1476 => x"86",
          1477 => x"78",
          1478 => x"38",
          1479 => x"08",
          1480 => x"82",
          1481 => x"fc",
          1482 => x"b4",
          1483 => x"11",
          1484 => x"05",
          1485 => x"3f",
          1486 => x"08",
          1487 => x"82",
          1488 => x"59",
          1489 => x"89",
          1490 => x"f4",
          1491 => x"cc",
          1492 => x"b9",
          1493 => x"80",
          1494 => x"82",
          1495 => x"43",
          1496 => x"86",
          1497 => x"78",
          1498 => x"38",
          1499 => x"08",
          1500 => x"82",
          1501 => x"59",
          1502 => x"88",
          1503 => x"8c",
          1504 => x"39",
          1505 => x"33",
          1506 => x"2e",
          1507 => x"86",
          1508 => x"88",
          1509 => x"a0",
          1510 => x"43",
          1511 => x"f8",
          1512 => x"84",
          1513 => x"d1",
          1514 => x"cc",
          1515 => x"a7",
          1516 => x"5c",
          1517 => x"2e",
          1518 => x"5c",
          1519 => x"70",
          1520 => x"07",
          1521 => x"7f",
          1522 => x"5a",
          1523 => x"2e",
          1524 => x"a0",
          1525 => x"88",
          1526 => x"e4",
          1527 => x"3f",
          1528 => x"54",
          1529 => x"52",
          1530 => x"ef",
          1531 => x"f4",
          1532 => x"3f",
          1533 => x"b4",
          1534 => x"11",
          1535 => x"05",
          1536 => x"3f",
          1537 => x"08",
          1538 => x"ec",
          1539 => x"fe",
          1540 => x"ff",
          1541 => x"a3",
          1542 => x"87",
          1543 => x"2e",
          1544 => x"59",
          1545 => x"05",
          1546 => x"63",
          1547 => x"b4",
          1548 => x"11",
          1549 => x"05",
          1550 => x"3f",
          1551 => x"08",
          1552 => x"b4",
          1553 => x"33",
          1554 => x"f4",
          1555 => x"b4",
          1556 => x"52",
          1557 => x"86",
          1558 => x"79",
          1559 => x"ae",
          1560 => x"38",
          1561 => x"9f",
          1562 => x"fe",
          1563 => x"ff",
          1564 => x"a3",
          1565 => x"87",
          1566 => x"2e",
          1567 => x"59",
          1568 => x"05",
          1569 => x"63",
          1570 => x"ff",
          1571 => x"f4",
          1572 => x"8c",
          1573 => x"39",
          1574 => x"f4",
          1575 => x"84",
          1576 => x"c7",
          1577 => x"cc",
          1578 => x"f4",
          1579 => x"3d",
          1580 => x"53",
          1581 => x"51",
          1582 => x"82",
          1583 => x"80",
          1584 => x"60",
          1585 => x"05",
          1586 => x"82",
          1587 => x"78",
          1588 => x"fe",
          1589 => x"ff",
          1590 => x"a4",
          1591 => x"87",
          1592 => x"38",
          1593 => x"60",
          1594 => x"52",
          1595 => x"51",
          1596 => x"80",
          1597 => x"51",
          1598 => x"79",
          1599 => x"59",
          1600 => x"f3",
          1601 => x"9f",
          1602 => x"60",
          1603 => x"d7",
          1604 => x"fe",
          1605 => x"ff",
          1606 => x"a3",
          1607 => x"87",
          1608 => x"2e",
          1609 => x"59",
          1610 => x"22",
          1611 => x"05",
          1612 => x"41",
          1613 => x"81",
          1614 => x"99",
          1615 => x"a7",
          1616 => x"fe",
          1617 => x"ff",
          1618 => x"a3",
          1619 => x"87",
          1620 => x"2e",
          1621 => x"b4",
          1622 => x"11",
          1623 => x"05",
          1624 => x"3f",
          1625 => x"08",
          1626 => x"38",
          1627 => x"0c",
          1628 => x"05",
          1629 => x"fe",
          1630 => x"ff",
          1631 => x"a2",
          1632 => x"87",
          1633 => x"38",
          1634 => x"60",
          1635 => x"52",
          1636 => x"51",
          1637 => x"80",
          1638 => x"51",
          1639 => x"79",
          1640 => x"59",
          1641 => x"f2",
          1642 => x"79",
          1643 => x"b4",
          1644 => x"11",
          1645 => x"05",
          1646 => x"3f",
          1647 => x"08",
          1648 => x"38",
          1649 => x"0c",
          1650 => x"05",
          1651 => x"39",
          1652 => x"51",
          1653 => x"ff",
          1654 => x"f4",
          1655 => x"c0",
          1656 => x"97",
          1657 => x"90",
          1658 => x"c4",
          1659 => x"3f",
          1660 => x"fc",
          1661 => x"39",
          1662 => x"51",
          1663 => x"84",
          1664 => x"87",
          1665 => x"0c",
          1666 => x"0b",
          1667 => x"94",
          1668 => x"39",
          1669 => x"51",
          1670 => x"8c",
          1671 => x"87",
          1672 => x"0c",
          1673 => x"0b",
          1674 => x"94",
          1675 => x"39",
          1676 => x"80",
          1677 => x"84",
          1678 => x"bd",
          1679 => x"cc",
          1680 => x"f1",
          1681 => x"52",
          1682 => x"51",
          1683 => x"63",
          1684 => x"b4",
          1685 => x"11",
          1686 => x"05",
          1687 => x"3f",
          1688 => x"08",
          1689 => x"90",
          1690 => x"81",
          1691 => x"9d",
          1692 => x"59",
          1693 => x"87",
          1694 => x"2e",
          1695 => x"82",
          1696 => x"52",
          1697 => x"51",
          1698 => x"f0",
          1699 => x"f5",
          1700 => x"8c",
          1701 => x"3f",
          1702 => x"81",
          1703 => x"96",
          1704 => x"59",
          1705 => x"90",
          1706 => x"cc",
          1707 => x"79",
          1708 => x"80",
          1709 => x"38",
          1710 => x"59",
          1711 => x"81",
          1712 => x"3d",
          1713 => x"51",
          1714 => x"82",
          1715 => x"5b",
          1716 => x"82",
          1717 => x"7b",
          1718 => x"38",
          1719 => x"8c",
          1720 => x"39",
          1721 => x"ae",
          1722 => x"39",
          1723 => x"56",
          1724 => x"f6",
          1725 => x"53",
          1726 => x"52",
          1727 => x"b0",
          1728 => x"96",
          1729 => x"81",
          1730 => x"b4",
          1731 => x"05",
          1732 => x"3f",
          1733 => x"55",
          1734 => x"54",
          1735 => x"f6",
          1736 => x"3d",
          1737 => x"51",
          1738 => x"92",
          1739 => x"80",
          1740 => x"ac",
          1741 => x"ff",
          1742 => x"9b",
          1743 => x"85",
          1744 => x"87",
          1745 => x"56",
          1746 => x"54",
          1747 => x"53",
          1748 => x"52",
          1749 => x"b0",
          1750 => x"b6",
          1751 => x"cc",
          1752 => x"cc",
          1753 => x"30",
          1754 => x"80",
          1755 => x"5b",
          1756 => x"7b",
          1757 => x"38",
          1758 => x"7a",
          1759 => x"80",
          1760 => x"81",
          1761 => x"ff",
          1762 => x"7b",
          1763 => x"7d",
          1764 => x"81",
          1765 => x"78",
          1766 => x"ff",
          1767 => x"06",
          1768 => x"81",
          1769 => x"9a",
          1770 => x"cc",
          1771 => x"0d",
          1772 => x"87",
          1773 => x"c0",
          1774 => x"08",
          1775 => x"84",
          1776 => x"51",
          1777 => x"82",
          1778 => x"90",
          1779 => x"55",
          1780 => x"80",
          1781 => x"b4",
          1782 => x"82",
          1783 => x"07",
          1784 => x"c0",
          1785 => x"08",
          1786 => x"84",
          1787 => x"51",
          1788 => x"82",
          1789 => x"90",
          1790 => x"55",
          1791 => x"80",
          1792 => x"b3",
          1793 => x"82",
          1794 => x"07",
          1795 => x"80",
          1796 => x"c0",
          1797 => x"8c",
          1798 => x"87",
          1799 => x"0c",
          1800 => x"82",
          1801 => x"80",
          1802 => x"82",
          1803 => x"89",
          1804 => x"fd",
          1805 => x"c4",
          1806 => x"3f",
          1807 => x"51",
          1808 => x"a1",
          1809 => x"a3",
          1810 => x"e8",
          1811 => x"d9",
          1812 => x"fe",
          1813 => x"52",
          1814 => x"88",
          1815 => x"c0",
          1816 => x"cc",
          1817 => x"06",
          1818 => x"14",
          1819 => x"80",
          1820 => x"71",
          1821 => x"0c",
          1822 => x"04",
          1823 => x"76",
          1824 => x"55",
          1825 => x"54",
          1826 => x"81",
          1827 => x"33",
          1828 => x"2e",
          1829 => x"86",
          1830 => x"53",
          1831 => x"33",
          1832 => x"2e",
          1833 => x"86",
          1834 => x"53",
          1835 => x"52",
          1836 => x"09",
          1837 => x"38",
          1838 => x"12",
          1839 => x"33",
          1840 => x"a2",
          1841 => x"81",
          1842 => x"2e",
          1843 => x"ea",
          1844 => x"81",
          1845 => x"72",
          1846 => x"70",
          1847 => x"38",
          1848 => x"80",
          1849 => x"73",
          1850 => x"72",
          1851 => x"70",
          1852 => x"81",
          1853 => x"81",
          1854 => x"32",
          1855 => x"80",
          1856 => x"51",
          1857 => x"80",
          1858 => x"80",
          1859 => x"05",
          1860 => x"75",
          1861 => x"70",
          1862 => x"0c",
          1863 => x"04",
          1864 => x"76",
          1865 => x"80",
          1866 => x"86",
          1867 => x"52",
          1868 => x"b7",
          1869 => x"cc",
          1870 => x"80",
          1871 => x"74",
          1872 => x"87",
          1873 => x"3d",
          1874 => x"3d",
          1875 => x"11",
          1876 => x"52",
          1877 => x"70",
          1878 => x"98",
          1879 => x"33",
          1880 => x"82",
          1881 => x"26",
          1882 => x"84",
          1883 => x"83",
          1884 => x"26",
          1885 => x"85",
          1886 => x"84",
          1887 => x"26",
          1888 => x"86",
          1889 => x"85",
          1890 => x"26",
          1891 => x"88",
          1892 => x"86",
          1893 => x"e7",
          1894 => x"38",
          1895 => x"54",
          1896 => x"87",
          1897 => x"cc",
          1898 => x"87",
          1899 => x"0c",
          1900 => x"c0",
          1901 => x"82",
          1902 => x"c0",
          1903 => x"83",
          1904 => x"c0",
          1905 => x"84",
          1906 => x"c0",
          1907 => x"85",
          1908 => x"c0",
          1909 => x"86",
          1910 => x"c0",
          1911 => x"74",
          1912 => x"a4",
          1913 => x"c0",
          1914 => x"80",
          1915 => x"98",
          1916 => x"52",
          1917 => x"cc",
          1918 => x"0d",
          1919 => x"0d",
          1920 => x"c0",
          1921 => x"81",
          1922 => x"c0",
          1923 => x"5e",
          1924 => x"87",
          1925 => x"08",
          1926 => x"1c",
          1927 => x"98",
          1928 => x"79",
          1929 => x"87",
          1930 => x"08",
          1931 => x"1c",
          1932 => x"98",
          1933 => x"79",
          1934 => x"87",
          1935 => x"08",
          1936 => x"1c",
          1937 => x"98",
          1938 => x"7b",
          1939 => x"87",
          1940 => x"08",
          1941 => x"1c",
          1942 => x"0c",
          1943 => x"ff",
          1944 => x"83",
          1945 => x"58",
          1946 => x"57",
          1947 => x"56",
          1948 => x"55",
          1949 => x"54",
          1950 => x"53",
          1951 => x"ff",
          1952 => x"f6",
          1953 => x"fc",
          1954 => x"0d",
          1955 => x"0d",
          1956 => x"33",
          1957 => x"9f",
          1958 => x"52",
          1959 => x"ec",
          1960 => x"0d",
          1961 => x"0d",
          1962 => x"ec",
          1963 => x"ff",
          1964 => x"56",
          1965 => x"84",
          1966 => x"2e",
          1967 => x"c0",
          1968 => x"70",
          1969 => x"2a",
          1970 => x"53",
          1971 => x"80",
          1972 => x"71",
          1973 => x"81",
          1974 => x"70",
          1975 => x"81",
          1976 => x"06",
          1977 => x"80",
          1978 => x"71",
          1979 => x"81",
          1980 => x"70",
          1981 => x"73",
          1982 => x"51",
          1983 => x"80",
          1984 => x"2e",
          1985 => x"c0",
          1986 => x"75",
          1987 => x"82",
          1988 => x"87",
          1989 => x"fb",
          1990 => x"9f",
          1991 => x"85",
          1992 => x"81",
          1993 => x"55",
          1994 => x"94",
          1995 => x"80",
          1996 => x"87",
          1997 => x"51",
          1998 => x"96",
          1999 => x"06",
          2000 => x"70",
          2001 => x"38",
          2002 => x"70",
          2003 => x"51",
          2004 => x"72",
          2005 => x"81",
          2006 => x"70",
          2007 => x"38",
          2008 => x"70",
          2009 => x"51",
          2010 => x"38",
          2011 => x"06",
          2012 => x"94",
          2013 => x"80",
          2014 => x"87",
          2015 => x"52",
          2016 => x"87",
          2017 => x"f9",
          2018 => x"54",
          2019 => x"70",
          2020 => x"53",
          2021 => x"77",
          2022 => x"38",
          2023 => x"06",
          2024 => x"85",
          2025 => x"81",
          2026 => x"57",
          2027 => x"c0",
          2028 => x"75",
          2029 => x"38",
          2030 => x"94",
          2031 => x"70",
          2032 => x"81",
          2033 => x"52",
          2034 => x"8c",
          2035 => x"2a",
          2036 => x"51",
          2037 => x"38",
          2038 => x"70",
          2039 => x"51",
          2040 => x"8d",
          2041 => x"2a",
          2042 => x"51",
          2043 => x"be",
          2044 => x"ff",
          2045 => x"c0",
          2046 => x"70",
          2047 => x"38",
          2048 => x"90",
          2049 => x"0c",
          2050 => x"33",
          2051 => x"06",
          2052 => x"70",
          2053 => x"76",
          2054 => x"0c",
          2055 => x"04",
          2056 => x"82",
          2057 => x"70",
          2058 => x"54",
          2059 => x"94",
          2060 => x"80",
          2061 => x"87",
          2062 => x"51",
          2063 => x"82",
          2064 => x"06",
          2065 => x"70",
          2066 => x"38",
          2067 => x"06",
          2068 => x"94",
          2069 => x"80",
          2070 => x"87",
          2071 => x"52",
          2072 => x"81",
          2073 => x"87",
          2074 => x"84",
          2075 => x"fe",
          2076 => x"85",
          2077 => x"81",
          2078 => x"53",
          2079 => x"84",
          2080 => x"2e",
          2081 => x"c0",
          2082 => x"71",
          2083 => x"2a",
          2084 => x"51",
          2085 => x"52",
          2086 => x"a0",
          2087 => x"ff",
          2088 => x"c0",
          2089 => x"70",
          2090 => x"38",
          2091 => x"90",
          2092 => x"70",
          2093 => x"98",
          2094 => x"51",
          2095 => x"cc",
          2096 => x"0d",
          2097 => x"0d",
          2098 => x"80",
          2099 => x"2a",
          2100 => x"51",
          2101 => x"84",
          2102 => x"c0",
          2103 => x"82",
          2104 => x"87",
          2105 => x"08",
          2106 => x"0c",
          2107 => x"94",
          2108 => x"f8",
          2109 => x"9e",
          2110 => x"85",
          2111 => x"c0",
          2112 => x"82",
          2113 => x"87",
          2114 => x"08",
          2115 => x"0c",
          2116 => x"ac",
          2117 => x"88",
          2118 => x"9e",
          2119 => x"86",
          2120 => x"c0",
          2121 => x"82",
          2122 => x"87",
          2123 => x"08",
          2124 => x"0c",
          2125 => x"bc",
          2126 => x"98",
          2127 => x"9e",
          2128 => x"86",
          2129 => x"c0",
          2130 => x"82",
          2131 => x"87",
          2132 => x"08",
          2133 => x"86",
          2134 => x"c0",
          2135 => x"82",
          2136 => x"87",
          2137 => x"08",
          2138 => x"0c",
          2139 => x"8c",
          2140 => x"b0",
          2141 => x"82",
          2142 => x"80",
          2143 => x"9e",
          2144 => x"84",
          2145 => x"51",
          2146 => x"80",
          2147 => x"81",
          2148 => x"86",
          2149 => x"0b",
          2150 => x"90",
          2151 => x"80",
          2152 => x"52",
          2153 => x"2e",
          2154 => x"52",
          2155 => x"b6",
          2156 => x"87",
          2157 => x"08",
          2158 => x"0a",
          2159 => x"52",
          2160 => x"83",
          2161 => x"71",
          2162 => x"34",
          2163 => x"c0",
          2164 => x"70",
          2165 => x"06",
          2166 => x"70",
          2167 => x"38",
          2168 => x"82",
          2169 => x"80",
          2170 => x"9e",
          2171 => x"a0",
          2172 => x"51",
          2173 => x"80",
          2174 => x"81",
          2175 => x"86",
          2176 => x"0b",
          2177 => x"90",
          2178 => x"80",
          2179 => x"52",
          2180 => x"2e",
          2181 => x"52",
          2182 => x"ba",
          2183 => x"87",
          2184 => x"08",
          2185 => x"80",
          2186 => x"52",
          2187 => x"83",
          2188 => x"71",
          2189 => x"34",
          2190 => x"c0",
          2191 => x"70",
          2192 => x"06",
          2193 => x"70",
          2194 => x"38",
          2195 => x"82",
          2196 => x"80",
          2197 => x"9e",
          2198 => x"81",
          2199 => x"51",
          2200 => x"80",
          2201 => x"81",
          2202 => x"86",
          2203 => x"0b",
          2204 => x"90",
          2205 => x"c0",
          2206 => x"52",
          2207 => x"2e",
          2208 => x"52",
          2209 => x"be",
          2210 => x"87",
          2211 => x"08",
          2212 => x"06",
          2213 => x"70",
          2214 => x"38",
          2215 => x"82",
          2216 => x"87",
          2217 => x"08",
          2218 => x"06",
          2219 => x"51",
          2220 => x"82",
          2221 => x"80",
          2222 => x"9e",
          2223 => x"84",
          2224 => x"52",
          2225 => x"2e",
          2226 => x"52",
          2227 => x"c1",
          2228 => x"9e",
          2229 => x"83",
          2230 => x"84",
          2231 => x"51",
          2232 => x"c2",
          2233 => x"87",
          2234 => x"08",
          2235 => x"51",
          2236 => x"80",
          2237 => x"81",
          2238 => x"86",
          2239 => x"c0",
          2240 => x"70",
          2241 => x"51",
          2242 => x"c4",
          2243 => x"0d",
          2244 => x"0d",
          2245 => x"51",
          2246 => x"82",
          2247 => x"54",
          2248 => x"88",
          2249 => x"94",
          2250 => x"3f",
          2251 => x"51",
          2252 => x"82",
          2253 => x"54",
          2254 => x"93",
          2255 => x"90",
          2256 => x"94",
          2257 => x"52",
          2258 => x"51",
          2259 => x"82",
          2260 => x"54",
          2261 => x"93",
          2262 => x"88",
          2263 => x"8c",
          2264 => x"52",
          2265 => x"51",
          2266 => x"82",
          2267 => x"54",
          2268 => x"93",
          2269 => x"f0",
          2270 => x"f4",
          2271 => x"52",
          2272 => x"51",
          2273 => x"82",
          2274 => x"54",
          2275 => x"93",
          2276 => x"f8",
          2277 => x"fc",
          2278 => x"52",
          2279 => x"51",
          2280 => x"82",
          2281 => x"54",
          2282 => x"93",
          2283 => x"80",
          2284 => x"84",
          2285 => x"52",
          2286 => x"51",
          2287 => x"82",
          2288 => x"54",
          2289 => x"8d",
          2290 => x"c0",
          2291 => x"f8",
          2292 => x"b0",
          2293 => x"c3",
          2294 => x"80",
          2295 => x"82",
          2296 => x"52",
          2297 => x"51",
          2298 => x"82",
          2299 => x"54",
          2300 => x"8d",
          2301 => x"c2",
          2302 => x"f9",
          2303 => x"84",
          2304 => x"b5",
          2305 => x"80",
          2306 => x"81",
          2307 => x"84",
          2308 => x"86",
          2309 => x"73",
          2310 => x"38",
          2311 => x"51",
          2312 => x"82",
          2313 => x"54",
          2314 => x"88",
          2315 => x"cc",
          2316 => x"3f",
          2317 => x"33",
          2318 => x"2e",
          2319 => x"f9",
          2320 => x"dc",
          2321 => x"be",
          2322 => x"80",
          2323 => x"81",
          2324 => x"83",
          2325 => x"f9",
          2326 => x"c4",
          2327 => x"98",
          2328 => x"f9",
          2329 => x"9c",
          2330 => x"9c",
          2331 => x"fa",
          2332 => x"90",
          2333 => x"a0",
          2334 => x"fa",
          2335 => x"84",
          2336 => x"f4",
          2337 => x"3f",
          2338 => x"22",
          2339 => x"fc",
          2340 => x"3f",
          2341 => x"08",
          2342 => x"c0",
          2343 => x"a2",
          2344 => x"87",
          2345 => x"84",
          2346 => x"71",
          2347 => x"82",
          2348 => x"52",
          2349 => x"51",
          2350 => x"82",
          2351 => x"54",
          2352 => x"a8",
          2353 => x"ac",
          2354 => x"84",
          2355 => x"51",
          2356 => x"82",
          2357 => x"bd",
          2358 => x"76",
          2359 => x"54",
          2360 => x"08",
          2361 => x"d0",
          2362 => x"3f",
          2363 => x"33",
          2364 => x"2e",
          2365 => x"86",
          2366 => x"bd",
          2367 => x"75",
          2368 => x"3f",
          2369 => x"08",
          2370 => x"29",
          2371 => x"54",
          2372 => x"cc",
          2373 => x"fb",
          2374 => x"e8",
          2375 => x"e4",
          2376 => x"3f",
          2377 => x"04",
          2378 => x"02",
          2379 => x"ff",
          2380 => x"84",
          2381 => x"71",
          2382 => x"e9",
          2383 => x"71",
          2384 => x"fc",
          2385 => x"39",
          2386 => x"51",
          2387 => x"fc",
          2388 => x"39",
          2389 => x"51",
          2390 => x"fc",
          2391 => x"39",
          2392 => x"51",
          2393 => x"84",
          2394 => x"71",
          2395 => x"04",
          2396 => x"87",
          2397 => x"70",
          2398 => x"80",
          2399 => x"74",
          2400 => x"86",
          2401 => x"0c",
          2402 => x"04",
          2403 => x"87",
          2404 => x"70",
          2405 => x"c8",
          2406 => x"72",
          2407 => x"70",
          2408 => x"08",
          2409 => x"86",
          2410 => x"0c",
          2411 => x"0d",
          2412 => x"87",
          2413 => x"0c",
          2414 => x"c8",
          2415 => x"96",
          2416 => x"fe",
          2417 => x"93",
          2418 => x"72",
          2419 => x"81",
          2420 => x"8d",
          2421 => x"82",
          2422 => x"52",
          2423 => x"90",
          2424 => x"34",
          2425 => x"08",
          2426 => x"9e",
          2427 => x"39",
          2428 => x"08",
          2429 => x"2e",
          2430 => x"51",
          2431 => x"3d",
          2432 => x"3d",
          2433 => x"05",
          2434 => x"d4",
          2435 => x"9e",
          2436 => x"51",
          2437 => x"72",
          2438 => x"0c",
          2439 => x"04",
          2440 => x"75",
          2441 => x"70",
          2442 => x"53",
          2443 => x"2e",
          2444 => x"81",
          2445 => x"81",
          2446 => x"87",
          2447 => x"85",
          2448 => x"fc",
          2449 => x"82",
          2450 => x"78",
          2451 => x"0c",
          2452 => x"33",
          2453 => x"06",
          2454 => x"80",
          2455 => x"72",
          2456 => x"51",
          2457 => x"fe",
          2458 => x"39",
          2459 => x"d4",
          2460 => x"0d",
          2461 => x"0d",
          2462 => x"59",
          2463 => x"05",
          2464 => x"75",
          2465 => x"f8",
          2466 => x"2e",
          2467 => x"82",
          2468 => x"70",
          2469 => x"05",
          2470 => x"5b",
          2471 => x"2e",
          2472 => x"85",
          2473 => x"8b",
          2474 => x"2e",
          2475 => x"8a",
          2476 => x"78",
          2477 => x"5a",
          2478 => x"aa",
          2479 => x"06",
          2480 => x"84",
          2481 => x"7b",
          2482 => x"5d",
          2483 => x"59",
          2484 => x"d0",
          2485 => x"89",
          2486 => x"7a",
          2487 => x"10",
          2488 => x"d0",
          2489 => x"81",
          2490 => x"57",
          2491 => x"75",
          2492 => x"70",
          2493 => x"07",
          2494 => x"80",
          2495 => x"30",
          2496 => x"80",
          2497 => x"53",
          2498 => x"55",
          2499 => x"2e",
          2500 => x"84",
          2501 => x"81",
          2502 => x"57",
          2503 => x"2e",
          2504 => x"75",
          2505 => x"76",
          2506 => x"e0",
          2507 => x"ff",
          2508 => x"73",
          2509 => x"81",
          2510 => x"80",
          2511 => x"38",
          2512 => x"2e",
          2513 => x"73",
          2514 => x"8b",
          2515 => x"c2",
          2516 => x"38",
          2517 => x"73",
          2518 => x"81",
          2519 => x"8f",
          2520 => x"d5",
          2521 => x"38",
          2522 => x"24",
          2523 => x"80",
          2524 => x"38",
          2525 => x"73",
          2526 => x"80",
          2527 => x"ef",
          2528 => x"19",
          2529 => x"59",
          2530 => x"33",
          2531 => x"75",
          2532 => x"81",
          2533 => x"70",
          2534 => x"55",
          2535 => x"79",
          2536 => x"90",
          2537 => x"16",
          2538 => x"7b",
          2539 => x"a0",
          2540 => x"3f",
          2541 => x"53",
          2542 => x"e9",
          2543 => x"fc",
          2544 => x"81",
          2545 => x"72",
          2546 => x"b0",
          2547 => x"fb",
          2548 => x"39",
          2549 => x"83",
          2550 => x"59",
          2551 => x"82",
          2552 => x"88",
          2553 => x"8a",
          2554 => x"90",
          2555 => x"75",
          2556 => x"3f",
          2557 => x"79",
          2558 => x"81",
          2559 => x"72",
          2560 => x"38",
          2561 => x"59",
          2562 => x"84",
          2563 => x"58",
          2564 => x"80",
          2565 => x"30",
          2566 => x"80",
          2567 => x"55",
          2568 => x"25",
          2569 => x"80",
          2570 => x"74",
          2571 => x"07",
          2572 => x"0b",
          2573 => x"57",
          2574 => x"51",
          2575 => x"82",
          2576 => x"81",
          2577 => x"53",
          2578 => x"9b",
          2579 => x"87",
          2580 => x"89",
          2581 => x"38",
          2582 => x"75",
          2583 => x"84",
          2584 => x"53",
          2585 => x"06",
          2586 => x"53",
          2587 => x"81",
          2588 => x"81",
          2589 => x"70",
          2590 => x"2a",
          2591 => x"76",
          2592 => x"38",
          2593 => x"38",
          2594 => x"70",
          2595 => x"53",
          2596 => x"8e",
          2597 => x"77",
          2598 => x"53",
          2599 => x"81",
          2600 => x"7a",
          2601 => x"55",
          2602 => x"83",
          2603 => x"79",
          2604 => x"81",
          2605 => x"72",
          2606 => x"17",
          2607 => x"27",
          2608 => x"51",
          2609 => x"75",
          2610 => x"72",
          2611 => x"81",
          2612 => x"7a",
          2613 => x"38",
          2614 => x"05",
          2615 => x"ff",
          2616 => x"70",
          2617 => x"57",
          2618 => x"76",
          2619 => x"81",
          2620 => x"72",
          2621 => x"84",
          2622 => x"f9",
          2623 => x"39",
          2624 => x"04",
          2625 => x"86",
          2626 => x"84",
          2627 => x"55",
          2628 => x"fa",
          2629 => x"3d",
          2630 => x"3d",
          2631 => x"9e",
          2632 => x"3d",
          2633 => x"75",
          2634 => x"3f",
          2635 => x"08",
          2636 => x"34",
          2637 => x"9e",
          2638 => x"3d",
          2639 => x"3d",
          2640 => x"d4",
          2641 => x"9e",
          2642 => x"3d",
          2643 => x"77",
          2644 => x"a1",
          2645 => x"9e",
          2646 => x"3d",
          2647 => x"3d",
          2648 => x"82",
          2649 => x"70",
          2650 => x"55",
          2651 => x"80",
          2652 => x"38",
          2653 => x"08",
          2654 => x"82",
          2655 => x"81",
          2656 => x"72",
          2657 => x"cb",
          2658 => x"2e",
          2659 => x"88",
          2660 => x"70",
          2661 => x"51",
          2662 => x"2e",
          2663 => x"80",
          2664 => x"ff",
          2665 => x"39",
          2666 => x"c8",
          2667 => x"52",
          2668 => x"c0",
          2669 => x"52",
          2670 => x"81",
          2671 => x"51",
          2672 => x"ff",
          2673 => x"15",
          2674 => x"34",
          2675 => x"f3",
          2676 => x"72",
          2677 => x"0c",
          2678 => x"04",
          2679 => x"82",
          2680 => x"75",
          2681 => x"0c",
          2682 => x"52",
          2683 => x"3f",
          2684 => x"d8",
          2685 => x"0d",
          2686 => x"0d",
          2687 => x"56",
          2688 => x"0c",
          2689 => x"70",
          2690 => x"73",
          2691 => x"81",
          2692 => x"81",
          2693 => x"ed",
          2694 => x"2e",
          2695 => x"8e",
          2696 => x"08",
          2697 => x"76",
          2698 => x"56",
          2699 => x"b0",
          2700 => x"06",
          2701 => x"75",
          2702 => x"76",
          2703 => x"70",
          2704 => x"73",
          2705 => x"8b",
          2706 => x"73",
          2707 => x"85",
          2708 => x"82",
          2709 => x"76",
          2710 => x"70",
          2711 => x"ac",
          2712 => x"a0",
          2713 => x"fa",
          2714 => x"53",
          2715 => x"57",
          2716 => x"98",
          2717 => x"39",
          2718 => x"80",
          2719 => x"26",
          2720 => x"86",
          2721 => x"80",
          2722 => x"57",
          2723 => x"74",
          2724 => x"38",
          2725 => x"27",
          2726 => x"14",
          2727 => x"06",
          2728 => x"14",
          2729 => x"06",
          2730 => x"74",
          2731 => x"f9",
          2732 => x"ff",
          2733 => x"89",
          2734 => x"38",
          2735 => x"c5",
          2736 => x"29",
          2737 => x"81",
          2738 => x"76",
          2739 => x"56",
          2740 => x"ba",
          2741 => x"2e",
          2742 => x"30",
          2743 => x"0c",
          2744 => x"82",
          2745 => x"8a",
          2746 => x"f8",
          2747 => x"7c",
          2748 => x"70",
          2749 => x"75",
          2750 => x"55",
          2751 => x"2e",
          2752 => x"87",
          2753 => x"76",
          2754 => x"73",
          2755 => x"81",
          2756 => x"81",
          2757 => x"77",
          2758 => x"70",
          2759 => x"58",
          2760 => x"09",
          2761 => x"c2",
          2762 => x"81",
          2763 => x"75",
          2764 => x"55",
          2765 => x"e2",
          2766 => x"90",
          2767 => x"f8",
          2768 => x"8f",
          2769 => x"81",
          2770 => x"75",
          2771 => x"55",
          2772 => x"81",
          2773 => x"27",
          2774 => x"d0",
          2775 => x"55",
          2776 => x"73",
          2777 => x"80",
          2778 => x"14",
          2779 => x"72",
          2780 => x"e0",
          2781 => x"80",
          2782 => x"39",
          2783 => x"55",
          2784 => x"80",
          2785 => x"e0",
          2786 => x"38",
          2787 => x"81",
          2788 => x"53",
          2789 => x"81",
          2790 => x"53",
          2791 => x"8e",
          2792 => x"70",
          2793 => x"55",
          2794 => x"27",
          2795 => x"77",
          2796 => x"74",
          2797 => x"76",
          2798 => x"77",
          2799 => x"70",
          2800 => x"55",
          2801 => x"77",
          2802 => x"38",
          2803 => x"74",
          2804 => x"55",
          2805 => x"cc",
          2806 => x"0d",
          2807 => x"0d",
          2808 => x"70",
          2809 => x"98",
          2810 => x"2c",
          2811 => x"70",
          2812 => x"53",
          2813 => x"51",
          2814 => x"fc",
          2815 => x"55",
          2816 => x"25",
          2817 => x"fc",
          2818 => x"12",
          2819 => x"97",
          2820 => x"33",
          2821 => x"70",
          2822 => x"81",
          2823 => x"81",
          2824 => x"87",
          2825 => x"3d",
          2826 => x"3d",
          2827 => x"84",
          2828 => x"33",
          2829 => x"55",
          2830 => x"2e",
          2831 => x"51",
          2832 => x"a0",
          2833 => x"3f",
          2834 => x"f7",
          2835 => x"ff",
          2836 => x"73",
          2837 => x"ff",
          2838 => x"39",
          2839 => x"c0",
          2840 => x"34",
          2841 => x"04",
          2842 => x"7c",
          2843 => x"b7",
          2844 => x"88",
          2845 => x"33",
          2846 => x"33",
          2847 => x"82",
          2848 => x"70",
          2849 => x"59",
          2850 => x"74",
          2851 => x"38",
          2852 => x"83",
          2853 => x"a4",
          2854 => x"29",
          2855 => x"05",
          2856 => x"54",
          2857 => x"a1",
          2858 => x"87",
          2859 => x"0c",
          2860 => x"33",
          2861 => x"82",
          2862 => x"70",
          2863 => x"5a",
          2864 => x"a7",
          2865 => x"78",
          2866 => x"ff",
          2867 => x"82",
          2868 => x"81",
          2869 => x"82",
          2870 => x"74",
          2871 => x"55",
          2872 => x"87",
          2873 => x"82",
          2874 => x"77",
          2875 => x"38",
          2876 => x"08",
          2877 => x"2e",
          2878 => x"87",
          2879 => x"74",
          2880 => x"3d",
          2881 => x"76",
          2882 => x"75",
          2883 => x"e9",
          2884 => x"a0",
          2885 => x"51",
          2886 => x"3f",
          2887 => x"08",
          2888 => x"c6",
          2889 => x"0d",
          2890 => x"0d",
          2891 => x"53",
          2892 => x"08",
          2893 => x"2e",
          2894 => x"51",
          2895 => x"80",
          2896 => x"14",
          2897 => x"54",
          2898 => x"e6",
          2899 => x"82",
          2900 => x"82",
          2901 => x"52",
          2902 => x"95",
          2903 => x"80",
          2904 => x"82",
          2905 => x"51",
          2906 => x"80",
          2907 => x"a0",
          2908 => x"0d",
          2909 => x"0d",
          2910 => x"52",
          2911 => x"08",
          2912 => x"93",
          2913 => x"cc",
          2914 => x"38",
          2915 => x"08",
          2916 => x"52",
          2917 => x"52",
          2918 => x"e1",
          2919 => x"cc",
          2920 => x"b9",
          2921 => x"ff",
          2922 => x"82",
          2923 => x"55",
          2924 => x"87",
          2925 => x"9c",
          2926 => x"cc",
          2927 => x"70",
          2928 => x"80",
          2929 => x"53",
          2930 => x"17",
          2931 => x"52",
          2932 => x"3f",
          2933 => x"09",
          2934 => x"b0",
          2935 => x"0d",
          2936 => x"0d",
          2937 => x"ad",
          2938 => x"5a",
          2939 => x"58",
          2940 => x"87",
          2941 => x"80",
          2942 => x"82",
          2943 => x"81",
          2944 => x"0b",
          2945 => x"08",
          2946 => x"f8",
          2947 => x"70",
          2948 => x"89",
          2949 => x"87",
          2950 => x"2e",
          2951 => x"51",
          2952 => x"3f",
          2953 => x"08",
          2954 => x"55",
          2955 => x"87",
          2956 => x"8e",
          2957 => x"cc",
          2958 => x"70",
          2959 => x"80",
          2960 => x"09",
          2961 => x"72",
          2962 => x"51",
          2963 => x"77",
          2964 => x"73",
          2965 => x"82",
          2966 => x"8c",
          2967 => x"51",
          2968 => x"3f",
          2969 => x"08",
          2970 => x"38",
          2971 => x"51",
          2972 => x"78",
          2973 => x"81",
          2974 => x"75",
          2975 => x"ff",
          2976 => x"79",
          2977 => x"af",
          2978 => x"08",
          2979 => x"cc",
          2980 => x"80",
          2981 => x"87",
          2982 => x"3d",
          2983 => x"3d",
          2984 => x"71",
          2985 => x"33",
          2986 => x"58",
          2987 => x"09",
          2988 => x"38",
          2989 => x"05",
          2990 => x"27",
          2991 => x"17",
          2992 => x"71",
          2993 => x"55",
          2994 => x"09",
          2995 => x"38",
          2996 => x"ea",
          2997 => x"73",
          2998 => x"87",
          2999 => x"08",
          3000 => x"b5",
          3001 => x"87",
          3002 => x"79",
          3003 => x"51",
          3004 => x"3f",
          3005 => x"08",
          3006 => x"84",
          3007 => x"74",
          3008 => x"38",
          3009 => x"88",
          3010 => x"fc",
          3011 => x"39",
          3012 => x"8c",
          3013 => x"53",
          3014 => x"f5",
          3015 => x"87",
          3016 => x"2e",
          3017 => x"1b",
          3018 => x"77",
          3019 => x"3f",
          3020 => x"08",
          3021 => x"55",
          3022 => x"74",
          3023 => x"81",
          3024 => x"ff",
          3025 => x"82",
          3026 => x"8b",
          3027 => x"73",
          3028 => x"0c",
          3029 => x"04",
          3030 => x"b0",
          3031 => x"3d",
          3032 => x"08",
          3033 => x"80",
          3034 => x"34",
          3035 => x"33",
          3036 => x"08",
          3037 => x"81",
          3038 => x"82",
          3039 => x"55",
          3040 => x"38",
          3041 => x"80",
          3042 => x"38",
          3043 => x"06",
          3044 => x"80",
          3045 => x"38",
          3046 => x"91",
          3047 => x"cc",
          3048 => x"a0",
          3049 => x"cc",
          3050 => x"81",
          3051 => x"53",
          3052 => x"87",
          3053 => x"80",
          3054 => x"82",
          3055 => x"80",
          3056 => x"82",
          3057 => x"f2",
          3058 => x"f7",
          3059 => x"cc",
          3060 => x"87",
          3061 => x"80",
          3062 => x"3d",
          3063 => x"81",
          3064 => x"82",
          3065 => x"56",
          3066 => x"08",
          3067 => x"81",
          3068 => x"38",
          3069 => x"08",
          3070 => x"bb",
          3071 => x"cc",
          3072 => x"0b",
          3073 => x"08",
          3074 => x"82",
          3075 => x"ff",
          3076 => x"55",
          3077 => x"34",
          3078 => x"81",
          3079 => x"75",
          3080 => x"3f",
          3081 => x"81",
          3082 => x"54",
          3083 => x"83",
          3084 => x"74",
          3085 => x"81",
          3086 => x"38",
          3087 => x"82",
          3088 => x"76",
          3089 => x"87",
          3090 => x"2e",
          3091 => x"d9",
          3092 => x"5d",
          3093 => x"82",
          3094 => x"98",
          3095 => x"2c",
          3096 => x"ff",
          3097 => x"78",
          3098 => x"82",
          3099 => x"70",
          3100 => x"98",
          3101 => x"e0",
          3102 => x"2b",
          3103 => x"71",
          3104 => x"70",
          3105 => x"fc",
          3106 => x"08",
          3107 => x"51",
          3108 => x"59",
          3109 => x"5d",
          3110 => x"73",
          3111 => x"e9",
          3112 => x"27",
          3113 => x"81",
          3114 => x"81",
          3115 => x"70",
          3116 => x"55",
          3117 => x"80",
          3118 => x"53",
          3119 => x"51",
          3120 => x"82",
          3121 => x"81",
          3122 => x"73",
          3123 => x"38",
          3124 => x"e0",
          3125 => x"b1",
          3126 => x"80",
          3127 => x"80",
          3128 => x"98",
          3129 => x"ff",
          3130 => x"55",
          3131 => x"97",
          3132 => x"74",
          3133 => x"f5",
          3134 => x"87",
          3135 => x"ff",
          3136 => x"cc",
          3137 => x"80",
          3138 => x"2e",
          3139 => x"81",
          3140 => x"82",
          3141 => x"74",
          3142 => x"98",
          3143 => x"e0",
          3144 => x"2b",
          3145 => x"70",
          3146 => x"82",
          3147 => x"d8",
          3148 => x"51",
          3149 => x"58",
          3150 => x"77",
          3151 => x"06",
          3152 => x"81",
          3153 => x"08",
          3154 => x"0b",
          3155 => x"34",
          3156 => x"9e",
          3157 => x"39",
          3158 => x"e4",
          3159 => x"9e",
          3160 => x"af",
          3161 => x"7d",
          3162 => x"73",
          3163 => x"e1",
          3164 => x"29",
          3165 => x"05",
          3166 => x"04",
          3167 => x"33",
          3168 => x"2e",
          3169 => x"82",
          3170 => x"55",
          3171 => x"ab",
          3172 => x"2b",
          3173 => x"51",
          3174 => x"24",
          3175 => x"1a",
          3176 => x"81",
          3177 => x"81",
          3178 => x"81",
          3179 => x"70",
          3180 => x"9e",
          3181 => x"51",
          3182 => x"82",
          3183 => x"81",
          3184 => x"74",
          3185 => x"34",
          3186 => x"ae",
          3187 => x"34",
          3188 => x"33",
          3189 => x"25",
          3190 => x"14",
          3191 => x"9e",
          3192 => x"9e",
          3193 => x"81",
          3194 => x"81",
          3195 => x"70",
          3196 => x"9e",
          3197 => x"51",
          3198 => x"77",
          3199 => x"74",
          3200 => x"52",
          3201 => x"3f",
          3202 => x"0a",
          3203 => x"0a",
          3204 => x"2c",
          3205 => x"33",
          3206 => x"73",
          3207 => x"38",
          3208 => x"33",
          3209 => x"70",
          3210 => x"9e",
          3211 => x"51",
          3212 => x"77",
          3213 => x"38",
          3214 => x"87",
          3215 => x"80",
          3216 => x"80",
          3217 => x"98",
          3218 => x"e8",
          3219 => x"55",
          3220 => x"e4",
          3221 => x"39",
          3222 => x"80",
          3223 => x"34",
          3224 => x"53",
          3225 => x"f5",
          3226 => x"be",
          3227 => x"39",
          3228 => x"33",
          3229 => x"06",
          3230 => x"80",
          3231 => x"38",
          3232 => x"33",
          3233 => x"73",
          3234 => x"34",
          3235 => x"73",
          3236 => x"34",
          3237 => x"ab",
          3238 => x"ec",
          3239 => x"2b",
          3240 => x"82",
          3241 => x"57",
          3242 => x"74",
          3243 => x"38",
          3244 => x"81",
          3245 => x"34",
          3246 => x"e6",
          3247 => x"81",
          3248 => x"81",
          3249 => x"70",
          3250 => x"9e",
          3251 => x"51",
          3252 => x"24",
          3253 => x"51",
          3254 => x"82",
          3255 => x"70",
          3256 => x"98",
          3257 => x"e8",
          3258 => x"56",
          3259 => x"24",
          3260 => x"88",
          3261 => x"3f",
          3262 => x"0a",
          3263 => x"0a",
          3264 => x"2c",
          3265 => x"33",
          3266 => x"75",
          3267 => x"38",
          3268 => x"82",
          3269 => x"7a",
          3270 => x"74",
          3271 => x"e5",
          3272 => x"9e",
          3273 => x"51",
          3274 => x"82",
          3275 => x"81",
          3276 => x"73",
          3277 => x"9e",
          3278 => x"73",
          3279 => x"38",
          3280 => x"52",
          3281 => x"a0",
          3282 => x"80",
          3283 => x"0b",
          3284 => x"34",
          3285 => x"9e",
          3286 => x"82",
          3287 => x"af",
          3288 => x"82",
          3289 => x"54",
          3290 => x"f9",
          3291 => x"51",
          3292 => x"82",
          3293 => x"ff",
          3294 => x"82",
          3295 => x"73",
          3296 => x"54",
          3297 => x"9e",
          3298 => x"9e",
          3299 => x"55",
          3300 => x"f9",
          3301 => x"14",
          3302 => x"9e",
          3303 => x"98",
          3304 => x"2c",
          3305 => x"06",
          3306 => x"74",
          3307 => x"38",
          3308 => x"81",
          3309 => x"34",
          3310 => x"e4",
          3311 => x"81",
          3312 => x"81",
          3313 => x"70",
          3314 => x"9e",
          3315 => x"51",
          3316 => x"24",
          3317 => x"51",
          3318 => x"82",
          3319 => x"70",
          3320 => x"98",
          3321 => x"e8",
          3322 => x"56",
          3323 => x"24",
          3324 => x"88",
          3325 => x"3f",
          3326 => x"0a",
          3327 => x"0a",
          3328 => x"2c",
          3329 => x"33",
          3330 => x"75",
          3331 => x"38",
          3332 => x"82",
          3333 => x"70",
          3334 => x"82",
          3335 => x"59",
          3336 => x"77",
          3337 => x"38",
          3338 => x"73",
          3339 => x"34",
          3340 => x"33",
          3341 => x"8b",
          3342 => x"ec",
          3343 => x"ff",
          3344 => x"e8",
          3345 => x"54",
          3346 => x"dc",
          3347 => x"39",
          3348 => x"53",
          3349 => x"f5",
          3350 => x"ce",
          3351 => x"82",
          3352 => x"80",
          3353 => x"e8",
          3354 => x"39",
          3355 => x"82",
          3356 => x"55",
          3357 => x"a6",
          3358 => x"ff",
          3359 => x"82",
          3360 => x"82",
          3361 => x"82",
          3362 => x"81",
          3363 => x"05",
          3364 => x"79",
          3365 => x"ff",
          3366 => x"81",
          3367 => x"84",
          3368 => x"cc",
          3369 => x"08",
          3370 => x"80",
          3371 => x"74",
          3372 => x"83",
          3373 => x"cc",
          3374 => x"e8",
          3375 => x"cc",
          3376 => x"06",
          3377 => x"74",
          3378 => x"ff",
          3379 => x"ff",
          3380 => x"fa",
          3381 => x"55",
          3382 => x"f6",
          3383 => x"51",
          3384 => x"3f",
          3385 => x"93",
          3386 => x"06",
          3387 => x"86",
          3388 => x"74",
          3389 => x"38",
          3390 => x"a9",
          3391 => x"87",
          3392 => x"9e",
          3393 => x"87",
          3394 => x"ff",
          3395 => x"53",
          3396 => x"51",
          3397 => x"3f",
          3398 => x"7a",
          3399 => x"86",
          3400 => x"08",
          3401 => x"80",
          3402 => x"74",
          3403 => x"87",
          3404 => x"cc",
          3405 => x"e8",
          3406 => x"cc",
          3407 => x"06",
          3408 => x"74",
          3409 => x"ff",
          3410 => x"81",
          3411 => x"81",
          3412 => x"89",
          3413 => x"9e",
          3414 => x"7a",
          3415 => x"ec",
          3416 => x"e8",
          3417 => x"51",
          3418 => x"f5",
          3419 => x"9e",
          3420 => x"81",
          3421 => x"9e",
          3422 => x"56",
          3423 => x"27",
          3424 => x"81",
          3425 => x"82",
          3426 => x"74",
          3427 => x"52",
          3428 => x"3f",
          3429 => x"82",
          3430 => x"54",
          3431 => x"f5",
          3432 => x"51",
          3433 => x"82",
          3434 => x"ff",
          3435 => x"82",
          3436 => x"f5",
          3437 => x"3d",
          3438 => x"2c",
          3439 => x"79",
          3440 => x"32",
          3441 => x"7c",
          3442 => x"32",
          3443 => x"71",
          3444 => x"55",
          3445 => x"57",
          3446 => x"82",
          3447 => x"74",
          3448 => x"82",
          3449 => x"87",
          3450 => x"fa",
          3451 => x"7a",
          3452 => x"52",
          3453 => x"8b",
          3454 => x"80",
          3455 => x"87",
          3456 => x"e0",
          3457 => x"80",
          3458 => x"74",
          3459 => x"3f",
          3460 => x"cc",
          3461 => x"80",
          3462 => x"26",
          3463 => x"74",
          3464 => x"2e",
          3465 => x"81",
          3466 => x"2a",
          3467 => x"77",
          3468 => x"54",
          3469 => x"56",
          3470 => x"a8",
          3471 => x"75",
          3472 => x"75",
          3473 => x"78",
          3474 => x"11",
          3475 => x"81",
          3476 => x"06",
          3477 => x"ff",
          3478 => x"52",
          3479 => x"56",
          3480 => x"38",
          3481 => x"07",
          3482 => x"87",
          3483 => x"3d",
          3484 => x"3d",
          3485 => x"fc",
          3486 => x"70",
          3487 => x"07",
          3488 => x"84",
          3489 => x"31",
          3490 => x"56",
          3491 => x"fe",
          3492 => x"30",
          3493 => x"83",
          3494 => x"31",
          3495 => x"59",
          3496 => x"77",
          3497 => x"70",
          3498 => x"25",
          3499 => x"71",
          3500 => x"2a",
          3501 => x"05",
          3502 => x"70",
          3503 => x"25",
          3504 => x"31",
          3505 => x"70",
          3506 => x"32",
          3507 => x"70",
          3508 => x"31",
          3509 => x"05",
          3510 => x"0c",
          3511 => x"52",
          3512 => x"53",
          3513 => x"51",
          3514 => x"53",
          3515 => x"3d",
          3516 => x"3d",
          3517 => x"70",
          3518 => x"54",
          3519 => x"3f",
          3520 => x"08",
          3521 => x"71",
          3522 => x"cc",
          3523 => x"3d",
          3524 => x"3d",
          3525 => x"57",
          3526 => x"75",
          3527 => x"38",
          3528 => x"ce",
          3529 => x"cc",
          3530 => x"12",
          3531 => x"2e",
          3532 => x"51",
          3533 => x"71",
          3534 => x"08",
          3535 => x"52",
          3536 => x"80",
          3537 => x"52",
          3538 => x"80",
          3539 => x"13",
          3540 => x"a0",
          3541 => x"71",
          3542 => x"55",
          3543 => x"72",
          3544 => x"38",
          3545 => x"9f",
          3546 => x"10",
          3547 => x"72",
          3548 => x"9f",
          3549 => x"06",
          3550 => x"75",
          3551 => x"1a",
          3552 => x"5b",
          3553 => x"54",
          3554 => x"73",
          3555 => x"87",
          3556 => x"3d",
          3557 => x"3d",
          3558 => x"80",
          3559 => x"c4",
          3560 => x"0b",
          3561 => x"23",
          3562 => x"80",
          3563 => x"80",
          3564 => x"b7",
          3565 => x"c4",
          3566 => x"58",
          3567 => x"81",
          3568 => x"15",
          3569 => x"c4",
          3570 => x"84",
          3571 => x"85",
          3572 => x"87",
          3573 => x"77",
          3574 => x"76",
          3575 => x"82",
          3576 => x"82",
          3577 => x"ff",
          3578 => x"80",
          3579 => x"ff",
          3580 => x"88",
          3581 => x"55",
          3582 => x"17",
          3583 => x"17",
          3584 => x"c0",
          3585 => x"29",
          3586 => x"08",
          3587 => x"51",
          3588 => x"82",
          3589 => x"83",
          3590 => x"3d",
          3591 => x"3d",
          3592 => x"81",
          3593 => x"27",
          3594 => x"12",
          3595 => x"11",
          3596 => x"ff",
          3597 => x"51",
          3598 => x"cc",
          3599 => x"0d",
          3600 => x"0d",
          3601 => x"22",
          3602 => x"aa",
          3603 => x"05",
          3604 => x"08",
          3605 => x"71",
          3606 => x"2b",
          3607 => x"33",
          3608 => x"71",
          3609 => x"02",
          3610 => x"05",
          3611 => x"ff",
          3612 => x"70",
          3613 => x"51",
          3614 => x"5b",
          3615 => x"54",
          3616 => x"34",
          3617 => x"34",
          3618 => x"08",
          3619 => x"2a",
          3620 => x"82",
          3621 => x"83",
          3622 => x"87",
          3623 => x"17",
          3624 => x"12",
          3625 => x"2b",
          3626 => x"2b",
          3627 => x"06",
          3628 => x"52",
          3629 => x"83",
          3630 => x"70",
          3631 => x"54",
          3632 => x"12",
          3633 => x"ff",
          3634 => x"83",
          3635 => x"87",
          3636 => x"56",
          3637 => x"72",
          3638 => x"89",
          3639 => x"fb",
          3640 => x"87",
          3641 => x"84",
          3642 => x"22",
          3643 => x"72",
          3644 => x"33",
          3645 => x"71",
          3646 => x"83",
          3647 => x"5b",
          3648 => x"52",
          3649 => x"12",
          3650 => x"33",
          3651 => x"07",
          3652 => x"54",
          3653 => x"70",
          3654 => x"73",
          3655 => x"82",
          3656 => x"70",
          3657 => x"33",
          3658 => x"71",
          3659 => x"83",
          3660 => x"59",
          3661 => x"05",
          3662 => x"87",
          3663 => x"88",
          3664 => x"88",
          3665 => x"56",
          3666 => x"13",
          3667 => x"13",
          3668 => x"c4",
          3669 => x"33",
          3670 => x"71",
          3671 => x"70",
          3672 => x"06",
          3673 => x"53",
          3674 => x"53",
          3675 => x"70",
          3676 => x"87",
          3677 => x"fa",
          3678 => x"a2",
          3679 => x"87",
          3680 => x"83",
          3681 => x"70",
          3682 => x"33",
          3683 => x"07",
          3684 => x"15",
          3685 => x"12",
          3686 => x"2b",
          3687 => x"07",
          3688 => x"55",
          3689 => x"57",
          3690 => x"80",
          3691 => x"38",
          3692 => x"ab",
          3693 => x"c4",
          3694 => x"70",
          3695 => x"33",
          3696 => x"71",
          3697 => x"74",
          3698 => x"81",
          3699 => x"88",
          3700 => x"83",
          3701 => x"f8",
          3702 => x"54",
          3703 => x"58",
          3704 => x"74",
          3705 => x"52",
          3706 => x"34",
          3707 => x"34",
          3708 => x"08",
          3709 => x"33",
          3710 => x"71",
          3711 => x"83",
          3712 => x"59",
          3713 => x"05",
          3714 => x"12",
          3715 => x"2b",
          3716 => x"ff",
          3717 => x"88",
          3718 => x"52",
          3719 => x"74",
          3720 => x"15",
          3721 => x"0d",
          3722 => x"0d",
          3723 => x"08",
          3724 => x"9e",
          3725 => x"83",
          3726 => x"82",
          3727 => x"12",
          3728 => x"2b",
          3729 => x"07",
          3730 => x"52",
          3731 => x"05",
          3732 => x"13",
          3733 => x"2b",
          3734 => x"05",
          3735 => x"71",
          3736 => x"2a",
          3737 => x"53",
          3738 => x"34",
          3739 => x"34",
          3740 => x"08",
          3741 => x"33",
          3742 => x"71",
          3743 => x"83",
          3744 => x"59",
          3745 => x"05",
          3746 => x"83",
          3747 => x"88",
          3748 => x"88",
          3749 => x"56",
          3750 => x"13",
          3751 => x"13",
          3752 => x"c4",
          3753 => x"11",
          3754 => x"33",
          3755 => x"07",
          3756 => x"0c",
          3757 => x"3d",
          3758 => x"3d",
          3759 => x"87",
          3760 => x"83",
          3761 => x"ff",
          3762 => x"53",
          3763 => x"a7",
          3764 => x"c4",
          3765 => x"2b",
          3766 => x"11",
          3767 => x"33",
          3768 => x"71",
          3769 => x"75",
          3770 => x"81",
          3771 => x"98",
          3772 => x"2b",
          3773 => x"40",
          3774 => x"58",
          3775 => x"72",
          3776 => x"38",
          3777 => x"52",
          3778 => x"9d",
          3779 => x"39",
          3780 => x"85",
          3781 => x"8b",
          3782 => x"2b",
          3783 => x"79",
          3784 => x"51",
          3785 => x"76",
          3786 => x"75",
          3787 => x"56",
          3788 => x"34",
          3789 => x"08",
          3790 => x"12",
          3791 => x"33",
          3792 => x"07",
          3793 => x"54",
          3794 => x"53",
          3795 => x"34",
          3796 => x"34",
          3797 => x"08",
          3798 => x"0b",
          3799 => x"80",
          3800 => x"34",
          3801 => x"08",
          3802 => x"14",
          3803 => x"14",
          3804 => x"c4",
          3805 => x"33",
          3806 => x"71",
          3807 => x"70",
          3808 => x"07",
          3809 => x"53",
          3810 => x"54",
          3811 => x"72",
          3812 => x"8b",
          3813 => x"ff",
          3814 => x"52",
          3815 => x"08",
          3816 => x"f2",
          3817 => x"2e",
          3818 => x"51",
          3819 => x"83",
          3820 => x"f5",
          3821 => x"7e",
          3822 => x"e2",
          3823 => x"cc",
          3824 => x"ff",
          3825 => x"c4",
          3826 => x"33",
          3827 => x"71",
          3828 => x"70",
          3829 => x"58",
          3830 => x"ff",
          3831 => x"2e",
          3832 => x"75",
          3833 => x"70",
          3834 => x"33",
          3835 => x"07",
          3836 => x"ff",
          3837 => x"70",
          3838 => x"06",
          3839 => x"52",
          3840 => x"59",
          3841 => x"27",
          3842 => x"80",
          3843 => x"75",
          3844 => x"84",
          3845 => x"16",
          3846 => x"2b",
          3847 => x"75",
          3848 => x"81",
          3849 => x"85",
          3850 => x"59",
          3851 => x"83",
          3852 => x"c4",
          3853 => x"33",
          3854 => x"71",
          3855 => x"70",
          3856 => x"06",
          3857 => x"56",
          3858 => x"75",
          3859 => x"81",
          3860 => x"79",
          3861 => x"cc",
          3862 => x"74",
          3863 => x"c4",
          3864 => x"2e",
          3865 => x"89",
          3866 => x"f8",
          3867 => x"ac",
          3868 => x"80",
          3869 => x"75",
          3870 => x"3f",
          3871 => x"08",
          3872 => x"11",
          3873 => x"33",
          3874 => x"71",
          3875 => x"53",
          3876 => x"74",
          3877 => x"70",
          3878 => x"06",
          3879 => x"5c",
          3880 => x"78",
          3881 => x"76",
          3882 => x"57",
          3883 => x"34",
          3884 => x"08",
          3885 => x"71",
          3886 => x"86",
          3887 => x"12",
          3888 => x"2b",
          3889 => x"2a",
          3890 => x"53",
          3891 => x"73",
          3892 => x"75",
          3893 => x"82",
          3894 => x"70",
          3895 => x"33",
          3896 => x"71",
          3897 => x"83",
          3898 => x"5d",
          3899 => x"05",
          3900 => x"15",
          3901 => x"15",
          3902 => x"c4",
          3903 => x"71",
          3904 => x"33",
          3905 => x"71",
          3906 => x"70",
          3907 => x"5a",
          3908 => x"54",
          3909 => x"34",
          3910 => x"34",
          3911 => x"08",
          3912 => x"54",
          3913 => x"cc",
          3914 => x"0d",
          3915 => x"0d",
          3916 => x"87",
          3917 => x"38",
          3918 => x"71",
          3919 => x"2e",
          3920 => x"51",
          3921 => x"82",
          3922 => x"53",
          3923 => x"cc",
          3924 => x"0d",
          3925 => x"0d",
          3926 => x"33",
          3927 => x"70",
          3928 => x"38",
          3929 => x"11",
          3930 => x"82",
          3931 => x"83",
          3932 => x"fc",
          3933 => x"9b",
          3934 => x"84",
          3935 => x"33",
          3936 => x"51",
          3937 => x"80",
          3938 => x"84",
          3939 => x"92",
          3940 => x"51",
          3941 => x"80",
          3942 => x"81",
          3943 => x"72",
          3944 => x"92",
          3945 => x"81",
          3946 => x"0b",
          3947 => x"8c",
          3948 => x"71",
          3949 => x"06",
          3950 => x"80",
          3951 => x"87",
          3952 => x"08",
          3953 => x"38",
          3954 => x"80",
          3955 => x"71",
          3956 => x"c0",
          3957 => x"51",
          3958 => x"87",
          3959 => x"87",
          3960 => x"82",
          3961 => x"33",
          3962 => x"87",
          3963 => x"3d",
          3964 => x"3d",
          3965 => x"64",
          3966 => x"bf",
          3967 => x"40",
          3968 => x"74",
          3969 => x"cd",
          3970 => x"cc",
          3971 => x"7a",
          3972 => x"81",
          3973 => x"72",
          3974 => x"87",
          3975 => x"11",
          3976 => x"8c",
          3977 => x"92",
          3978 => x"5a",
          3979 => x"58",
          3980 => x"c0",
          3981 => x"76",
          3982 => x"76",
          3983 => x"70",
          3984 => x"81",
          3985 => x"54",
          3986 => x"8e",
          3987 => x"52",
          3988 => x"81",
          3989 => x"81",
          3990 => x"74",
          3991 => x"53",
          3992 => x"83",
          3993 => x"78",
          3994 => x"8f",
          3995 => x"2e",
          3996 => x"c0",
          3997 => x"52",
          3998 => x"87",
          3999 => x"08",
          4000 => x"2e",
          4001 => x"84",
          4002 => x"38",
          4003 => x"87",
          4004 => x"15",
          4005 => x"70",
          4006 => x"52",
          4007 => x"ff",
          4008 => x"39",
          4009 => x"81",
          4010 => x"ff",
          4011 => x"57",
          4012 => x"90",
          4013 => x"80",
          4014 => x"71",
          4015 => x"78",
          4016 => x"38",
          4017 => x"80",
          4018 => x"80",
          4019 => x"81",
          4020 => x"72",
          4021 => x"0c",
          4022 => x"04",
          4023 => x"60",
          4024 => x"8c",
          4025 => x"33",
          4026 => x"5b",
          4027 => x"74",
          4028 => x"e1",
          4029 => x"cc",
          4030 => x"79",
          4031 => x"78",
          4032 => x"06",
          4033 => x"77",
          4034 => x"87",
          4035 => x"11",
          4036 => x"8c",
          4037 => x"92",
          4038 => x"59",
          4039 => x"85",
          4040 => x"98",
          4041 => x"7d",
          4042 => x"0c",
          4043 => x"08",
          4044 => x"70",
          4045 => x"53",
          4046 => x"2e",
          4047 => x"70",
          4048 => x"33",
          4049 => x"18",
          4050 => x"2a",
          4051 => x"51",
          4052 => x"2e",
          4053 => x"c0",
          4054 => x"52",
          4055 => x"87",
          4056 => x"08",
          4057 => x"2e",
          4058 => x"84",
          4059 => x"38",
          4060 => x"87",
          4061 => x"15",
          4062 => x"70",
          4063 => x"52",
          4064 => x"ff",
          4065 => x"39",
          4066 => x"81",
          4067 => x"80",
          4068 => x"52",
          4069 => x"90",
          4070 => x"80",
          4071 => x"71",
          4072 => x"7a",
          4073 => x"38",
          4074 => x"80",
          4075 => x"80",
          4076 => x"81",
          4077 => x"72",
          4078 => x"0c",
          4079 => x"04",
          4080 => x"7a",
          4081 => x"a3",
          4082 => x"88",
          4083 => x"33",
          4084 => x"56",
          4085 => x"3f",
          4086 => x"08",
          4087 => x"83",
          4088 => x"fe",
          4089 => x"87",
          4090 => x"0c",
          4091 => x"76",
          4092 => x"38",
          4093 => x"93",
          4094 => x"2b",
          4095 => x"8c",
          4096 => x"71",
          4097 => x"38",
          4098 => x"71",
          4099 => x"c6",
          4100 => x"39",
          4101 => x"81",
          4102 => x"06",
          4103 => x"71",
          4104 => x"38",
          4105 => x"8c",
          4106 => x"e8",
          4107 => x"98",
          4108 => x"71",
          4109 => x"73",
          4110 => x"92",
          4111 => x"72",
          4112 => x"06",
          4113 => x"f7",
          4114 => x"80",
          4115 => x"88",
          4116 => x"0c",
          4117 => x"80",
          4118 => x"56",
          4119 => x"56",
          4120 => x"82",
          4121 => x"88",
          4122 => x"fe",
          4123 => x"81",
          4124 => x"33",
          4125 => x"07",
          4126 => x"0c",
          4127 => x"3d",
          4128 => x"3d",
          4129 => x"11",
          4130 => x"33",
          4131 => x"71",
          4132 => x"81",
          4133 => x"72",
          4134 => x"75",
          4135 => x"82",
          4136 => x"52",
          4137 => x"54",
          4138 => x"0d",
          4139 => x"0d",
          4140 => x"05",
          4141 => x"52",
          4142 => x"70",
          4143 => x"34",
          4144 => x"51",
          4145 => x"83",
          4146 => x"ff",
          4147 => x"75",
          4148 => x"72",
          4149 => x"54",
          4150 => x"2a",
          4151 => x"70",
          4152 => x"34",
          4153 => x"51",
          4154 => x"81",
          4155 => x"70",
          4156 => x"70",
          4157 => x"3d",
          4158 => x"3d",
          4159 => x"77",
          4160 => x"70",
          4161 => x"38",
          4162 => x"05",
          4163 => x"70",
          4164 => x"34",
          4165 => x"eb",
          4166 => x"0d",
          4167 => x"0d",
          4168 => x"54",
          4169 => x"72",
          4170 => x"54",
          4171 => x"51",
          4172 => x"84",
          4173 => x"fc",
          4174 => x"77",
          4175 => x"53",
          4176 => x"05",
          4177 => x"70",
          4178 => x"33",
          4179 => x"ff",
          4180 => x"52",
          4181 => x"2e",
          4182 => x"80",
          4183 => x"71",
          4184 => x"0c",
          4185 => x"04",
          4186 => x"74",
          4187 => x"89",
          4188 => x"2e",
          4189 => x"11",
          4190 => x"52",
          4191 => x"70",
          4192 => x"cc",
          4193 => x"0d",
          4194 => x"82",
          4195 => x"04",
          4196 => x"87",
          4197 => x"f7",
          4198 => x"56",
          4199 => x"17",
          4200 => x"74",
          4201 => x"d6",
          4202 => x"b0",
          4203 => x"b4",
          4204 => x"81",
          4205 => x"59",
          4206 => x"82",
          4207 => x"7a",
          4208 => x"06",
          4209 => x"87",
          4210 => x"17",
          4211 => x"08",
          4212 => x"08",
          4213 => x"08",
          4214 => x"74",
          4215 => x"38",
          4216 => x"55",
          4217 => x"09",
          4218 => x"38",
          4219 => x"18",
          4220 => x"81",
          4221 => x"f9",
          4222 => x"39",
          4223 => x"82",
          4224 => x"8b",
          4225 => x"fa",
          4226 => x"7a",
          4227 => x"57",
          4228 => x"08",
          4229 => x"75",
          4230 => x"3f",
          4231 => x"08",
          4232 => x"cc",
          4233 => x"81",
          4234 => x"b4",
          4235 => x"16",
          4236 => x"be",
          4237 => x"cc",
          4238 => x"85",
          4239 => x"81",
          4240 => x"17",
          4241 => x"87",
          4242 => x"3d",
          4243 => x"3d",
          4244 => x"52",
          4245 => x"3f",
          4246 => x"08",
          4247 => x"cc",
          4248 => x"38",
          4249 => x"74",
          4250 => x"81",
          4251 => x"38",
          4252 => x"59",
          4253 => x"09",
          4254 => x"e3",
          4255 => x"53",
          4256 => x"08",
          4257 => x"70",
          4258 => x"91",
          4259 => x"d5",
          4260 => x"17",
          4261 => x"3f",
          4262 => x"a4",
          4263 => x"51",
          4264 => x"86",
          4265 => x"f2",
          4266 => x"17",
          4267 => x"3f",
          4268 => x"52",
          4269 => x"51",
          4270 => x"8c",
          4271 => x"84",
          4272 => x"fc",
          4273 => x"17",
          4274 => x"70",
          4275 => x"79",
          4276 => x"52",
          4277 => x"51",
          4278 => x"77",
          4279 => x"80",
          4280 => x"81",
          4281 => x"f9",
          4282 => x"87",
          4283 => x"2e",
          4284 => x"58",
          4285 => x"cc",
          4286 => x"0d",
          4287 => x"0d",
          4288 => x"98",
          4289 => x"05",
          4290 => x"80",
          4291 => x"27",
          4292 => x"14",
          4293 => x"29",
          4294 => x"05",
          4295 => x"82",
          4296 => x"87",
          4297 => x"f9",
          4298 => x"7a",
          4299 => x"54",
          4300 => x"27",
          4301 => x"76",
          4302 => x"27",
          4303 => x"ff",
          4304 => x"58",
          4305 => x"80",
          4306 => x"82",
          4307 => x"72",
          4308 => x"38",
          4309 => x"72",
          4310 => x"8e",
          4311 => x"39",
          4312 => x"17",
          4313 => x"a4",
          4314 => x"53",
          4315 => x"fd",
          4316 => x"87",
          4317 => x"9f",
          4318 => x"ff",
          4319 => x"11",
          4320 => x"70",
          4321 => x"18",
          4322 => x"76",
          4323 => x"53",
          4324 => x"82",
          4325 => x"80",
          4326 => x"83",
          4327 => x"b4",
          4328 => x"88",
          4329 => x"79",
          4330 => x"84",
          4331 => x"58",
          4332 => x"80",
          4333 => x"9f",
          4334 => x"80",
          4335 => x"88",
          4336 => x"08",
          4337 => x"51",
          4338 => x"82",
          4339 => x"80",
          4340 => x"10",
          4341 => x"74",
          4342 => x"51",
          4343 => x"82",
          4344 => x"83",
          4345 => x"58",
          4346 => x"87",
          4347 => x"08",
          4348 => x"51",
          4349 => x"82",
          4350 => x"9b",
          4351 => x"2b",
          4352 => x"74",
          4353 => x"51",
          4354 => x"82",
          4355 => x"f0",
          4356 => x"83",
          4357 => x"77",
          4358 => x"0c",
          4359 => x"04",
          4360 => x"7a",
          4361 => x"58",
          4362 => x"81",
          4363 => x"9e",
          4364 => x"17",
          4365 => x"96",
          4366 => x"53",
          4367 => x"81",
          4368 => x"79",
          4369 => x"72",
          4370 => x"38",
          4371 => x"72",
          4372 => x"b8",
          4373 => x"39",
          4374 => x"17",
          4375 => x"a4",
          4376 => x"53",
          4377 => x"fb",
          4378 => x"87",
          4379 => x"82",
          4380 => x"81",
          4381 => x"83",
          4382 => x"b4",
          4383 => x"78",
          4384 => x"56",
          4385 => x"76",
          4386 => x"38",
          4387 => x"9f",
          4388 => x"33",
          4389 => x"07",
          4390 => x"74",
          4391 => x"83",
          4392 => x"89",
          4393 => x"08",
          4394 => x"51",
          4395 => x"82",
          4396 => x"59",
          4397 => x"08",
          4398 => x"74",
          4399 => x"16",
          4400 => x"84",
          4401 => x"76",
          4402 => x"88",
          4403 => x"81",
          4404 => x"8f",
          4405 => x"53",
          4406 => x"80",
          4407 => x"88",
          4408 => x"08",
          4409 => x"51",
          4410 => x"82",
          4411 => x"59",
          4412 => x"08",
          4413 => x"77",
          4414 => x"06",
          4415 => x"83",
          4416 => x"05",
          4417 => x"f7",
          4418 => x"39",
          4419 => x"a4",
          4420 => x"52",
          4421 => x"ef",
          4422 => x"cc",
          4423 => x"87",
          4424 => x"38",
          4425 => x"06",
          4426 => x"83",
          4427 => x"18",
          4428 => x"54",
          4429 => x"f6",
          4430 => x"87",
          4431 => x"0a",
          4432 => x"52",
          4433 => x"83",
          4434 => x"83",
          4435 => x"82",
          4436 => x"8a",
          4437 => x"f8",
          4438 => x"7c",
          4439 => x"59",
          4440 => x"81",
          4441 => x"38",
          4442 => x"08",
          4443 => x"73",
          4444 => x"38",
          4445 => x"52",
          4446 => x"a4",
          4447 => x"cc",
          4448 => x"87",
          4449 => x"f2",
          4450 => x"82",
          4451 => x"39",
          4452 => x"e6",
          4453 => x"cc",
          4454 => x"de",
          4455 => x"78",
          4456 => x"3f",
          4457 => x"08",
          4458 => x"cc",
          4459 => x"80",
          4460 => x"87",
          4461 => x"2e",
          4462 => x"87",
          4463 => x"2e",
          4464 => x"53",
          4465 => x"51",
          4466 => x"82",
          4467 => x"c5",
          4468 => x"08",
          4469 => x"18",
          4470 => x"57",
          4471 => x"90",
          4472 => x"90",
          4473 => x"16",
          4474 => x"54",
          4475 => x"34",
          4476 => x"78",
          4477 => x"38",
          4478 => x"82",
          4479 => x"8a",
          4480 => x"f6",
          4481 => x"7e",
          4482 => x"5b",
          4483 => x"38",
          4484 => x"58",
          4485 => x"88",
          4486 => x"08",
          4487 => x"38",
          4488 => x"39",
          4489 => x"51",
          4490 => x"81",
          4491 => x"87",
          4492 => x"82",
          4493 => x"87",
          4494 => x"82",
          4495 => x"ff",
          4496 => x"38",
          4497 => x"82",
          4498 => x"26",
          4499 => x"79",
          4500 => x"08",
          4501 => x"73",
          4502 => x"b9",
          4503 => x"2e",
          4504 => x"80",
          4505 => x"1a",
          4506 => x"08",
          4507 => x"38",
          4508 => x"52",
          4509 => x"af",
          4510 => x"82",
          4511 => x"81",
          4512 => x"06",
          4513 => x"87",
          4514 => x"82",
          4515 => x"09",
          4516 => x"72",
          4517 => x"70",
          4518 => x"87",
          4519 => x"51",
          4520 => x"73",
          4521 => x"82",
          4522 => x"80",
          4523 => x"8c",
          4524 => x"81",
          4525 => x"38",
          4526 => x"08",
          4527 => x"73",
          4528 => x"75",
          4529 => x"77",
          4530 => x"56",
          4531 => x"76",
          4532 => x"82",
          4533 => x"26",
          4534 => x"75",
          4535 => x"f8",
          4536 => x"87",
          4537 => x"2e",
          4538 => x"59",
          4539 => x"08",
          4540 => x"81",
          4541 => x"82",
          4542 => x"59",
          4543 => x"08",
          4544 => x"70",
          4545 => x"25",
          4546 => x"51",
          4547 => x"73",
          4548 => x"75",
          4549 => x"81",
          4550 => x"38",
          4551 => x"f5",
          4552 => x"75",
          4553 => x"f9",
          4554 => x"87",
          4555 => x"87",
          4556 => x"70",
          4557 => x"08",
          4558 => x"51",
          4559 => x"80",
          4560 => x"73",
          4561 => x"38",
          4562 => x"52",
          4563 => x"d0",
          4564 => x"cc",
          4565 => x"a5",
          4566 => x"18",
          4567 => x"08",
          4568 => x"18",
          4569 => x"74",
          4570 => x"38",
          4571 => x"18",
          4572 => x"33",
          4573 => x"73",
          4574 => x"97",
          4575 => x"74",
          4576 => x"38",
          4577 => x"55",
          4578 => x"87",
          4579 => x"85",
          4580 => x"75",
          4581 => x"87",
          4582 => x"3d",
          4583 => x"3d",
          4584 => x"52",
          4585 => x"3f",
          4586 => x"08",
          4587 => x"82",
          4588 => x"80",
          4589 => x"52",
          4590 => x"c1",
          4591 => x"cc",
          4592 => x"cc",
          4593 => x"0c",
          4594 => x"53",
          4595 => x"15",
          4596 => x"f2",
          4597 => x"56",
          4598 => x"16",
          4599 => x"22",
          4600 => x"27",
          4601 => x"54",
          4602 => x"76",
          4603 => x"33",
          4604 => x"3f",
          4605 => x"08",
          4606 => x"38",
          4607 => x"76",
          4608 => x"70",
          4609 => x"9f",
          4610 => x"56",
          4611 => x"87",
          4612 => x"3d",
          4613 => x"3d",
          4614 => x"71",
          4615 => x"57",
          4616 => x"0a",
          4617 => x"38",
          4618 => x"53",
          4619 => x"38",
          4620 => x"0c",
          4621 => x"54",
          4622 => x"75",
          4623 => x"73",
          4624 => x"a8",
          4625 => x"73",
          4626 => x"85",
          4627 => x"0b",
          4628 => x"5a",
          4629 => x"27",
          4630 => x"a8",
          4631 => x"18",
          4632 => x"39",
          4633 => x"70",
          4634 => x"58",
          4635 => x"b2",
          4636 => x"76",
          4637 => x"3f",
          4638 => x"08",
          4639 => x"cc",
          4640 => x"bd",
          4641 => x"82",
          4642 => x"27",
          4643 => x"16",
          4644 => x"cc",
          4645 => x"38",
          4646 => x"39",
          4647 => x"55",
          4648 => x"52",
          4649 => x"d5",
          4650 => x"cc",
          4651 => x"0c",
          4652 => x"0c",
          4653 => x"53",
          4654 => x"80",
          4655 => x"85",
          4656 => x"94",
          4657 => x"2a",
          4658 => x"0c",
          4659 => x"06",
          4660 => x"9c",
          4661 => x"58",
          4662 => x"cc",
          4663 => x"0d",
          4664 => x"0d",
          4665 => x"90",
          4666 => x"05",
          4667 => x"f0",
          4668 => x"27",
          4669 => x"0b",
          4670 => x"98",
          4671 => x"84",
          4672 => x"2e",
          4673 => x"76",
          4674 => x"58",
          4675 => x"38",
          4676 => x"15",
          4677 => x"08",
          4678 => x"38",
          4679 => x"88",
          4680 => x"53",
          4681 => x"81",
          4682 => x"c0",
          4683 => x"22",
          4684 => x"89",
          4685 => x"72",
          4686 => x"74",
          4687 => x"f3",
          4688 => x"87",
          4689 => x"82",
          4690 => x"82",
          4691 => x"27",
          4692 => x"81",
          4693 => x"cc",
          4694 => x"80",
          4695 => x"16",
          4696 => x"cc",
          4697 => x"ca",
          4698 => x"38",
          4699 => x"0c",
          4700 => x"dd",
          4701 => x"08",
          4702 => x"f9",
          4703 => x"87",
          4704 => x"87",
          4705 => x"cc",
          4706 => x"80",
          4707 => x"55",
          4708 => x"08",
          4709 => x"38",
          4710 => x"87",
          4711 => x"2e",
          4712 => x"87",
          4713 => x"75",
          4714 => x"3f",
          4715 => x"08",
          4716 => x"94",
          4717 => x"52",
          4718 => x"c1",
          4719 => x"cc",
          4720 => x"0c",
          4721 => x"0c",
          4722 => x"05",
          4723 => x"80",
          4724 => x"87",
          4725 => x"3d",
          4726 => x"3d",
          4727 => x"71",
          4728 => x"57",
          4729 => x"51",
          4730 => x"82",
          4731 => x"54",
          4732 => x"08",
          4733 => x"82",
          4734 => x"56",
          4735 => x"52",
          4736 => x"83",
          4737 => x"cc",
          4738 => x"87",
          4739 => x"d2",
          4740 => x"cc",
          4741 => x"08",
          4742 => x"54",
          4743 => x"e5",
          4744 => x"06",
          4745 => x"58",
          4746 => x"08",
          4747 => x"38",
          4748 => x"75",
          4749 => x"80",
          4750 => x"81",
          4751 => x"7a",
          4752 => x"06",
          4753 => x"39",
          4754 => x"08",
          4755 => x"76",
          4756 => x"3f",
          4757 => x"08",
          4758 => x"cc",
          4759 => x"ff",
          4760 => x"84",
          4761 => x"06",
          4762 => x"54",
          4763 => x"cc",
          4764 => x"0d",
          4765 => x"0d",
          4766 => x"52",
          4767 => x"3f",
          4768 => x"08",
          4769 => x"06",
          4770 => x"51",
          4771 => x"83",
          4772 => x"06",
          4773 => x"14",
          4774 => x"3f",
          4775 => x"08",
          4776 => x"07",
          4777 => x"87",
          4778 => x"3d",
          4779 => x"3d",
          4780 => x"70",
          4781 => x"06",
          4782 => x"53",
          4783 => x"ed",
          4784 => x"33",
          4785 => x"83",
          4786 => x"06",
          4787 => x"90",
          4788 => x"15",
          4789 => x"3f",
          4790 => x"04",
          4791 => x"7b",
          4792 => x"84",
          4793 => x"58",
          4794 => x"80",
          4795 => x"38",
          4796 => x"52",
          4797 => x"8f",
          4798 => x"cc",
          4799 => x"87",
          4800 => x"f5",
          4801 => x"08",
          4802 => x"53",
          4803 => x"84",
          4804 => x"39",
          4805 => x"70",
          4806 => x"81",
          4807 => x"51",
          4808 => x"16",
          4809 => x"cc",
          4810 => x"81",
          4811 => x"38",
          4812 => x"ae",
          4813 => x"81",
          4814 => x"54",
          4815 => x"2e",
          4816 => x"8f",
          4817 => x"82",
          4818 => x"76",
          4819 => x"54",
          4820 => x"09",
          4821 => x"38",
          4822 => x"7a",
          4823 => x"80",
          4824 => x"fa",
          4825 => x"87",
          4826 => x"82",
          4827 => x"89",
          4828 => x"08",
          4829 => x"86",
          4830 => x"98",
          4831 => x"82",
          4832 => x"8b",
          4833 => x"fb",
          4834 => x"70",
          4835 => x"81",
          4836 => x"fc",
          4837 => x"87",
          4838 => x"82",
          4839 => x"b4",
          4840 => x"08",
          4841 => x"ec",
          4842 => x"87",
          4843 => x"82",
          4844 => x"a0",
          4845 => x"82",
          4846 => x"52",
          4847 => x"51",
          4848 => x"8b",
          4849 => x"52",
          4850 => x"51",
          4851 => x"81",
          4852 => x"34",
          4853 => x"cc",
          4854 => x"0d",
          4855 => x"0d",
          4856 => x"98",
          4857 => x"70",
          4858 => x"ec",
          4859 => x"87",
          4860 => x"38",
          4861 => x"53",
          4862 => x"81",
          4863 => x"34",
          4864 => x"04",
          4865 => x"78",
          4866 => x"80",
          4867 => x"34",
          4868 => x"80",
          4869 => x"38",
          4870 => x"18",
          4871 => x"9c",
          4872 => x"70",
          4873 => x"56",
          4874 => x"a0",
          4875 => x"71",
          4876 => x"81",
          4877 => x"81",
          4878 => x"89",
          4879 => x"06",
          4880 => x"73",
          4881 => x"55",
          4882 => x"55",
          4883 => x"81",
          4884 => x"81",
          4885 => x"74",
          4886 => x"75",
          4887 => x"52",
          4888 => x"13",
          4889 => x"08",
          4890 => x"33",
          4891 => x"9c",
          4892 => x"11",
          4893 => x"8a",
          4894 => x"cc",
          4895 => x"96",
          4896 => x"e7",
          4897 => x"cc",
          4898 => x"23",
          4899 => x"e7",
          4900 => x"87",
          4901 => x"17",
          4902 => x"0d",
          4903 => x"0d",
          4904 => x"5e",
          4905 => x"70",
          4906 => x"55",
          4907 => x"83",
          4908 => x"73",
          4909 => x"91",
          4910 => x"2e",
          4911 => x"1d",
          4912 => x"0c",
          4913 => x"15",
          4914 => x"70",
          4915 => x"56",
          4916 => x"09",
          4917 => x"38",
          4918 => x"80",
          4919 => x"30",
          4920 => x"78",
          4921 => x"54",
          4922 => x"73",
          4923 => x"60",
          4924 => x"54",
          4925 => x"96",
          4926 => x"0b",
          4927 => x"80",
          4928 => x"f6",
          4929 => x"87",
          4930 => x"85",
          4931 => x"3d",
          4932 => x"5c",
          4933 => x"53",
          4934 => x"51",
          4935 => x"80",
          4936 => x"88",
          4937 => x"5c",
          4938 => x"09",
          4939 => x"d4",
          4940 => x"70",
          4941 => x"71",
          4942 => x"30",
          4943 => x"73",
          4944 => x"51",
          4945 => x"57",
          4946 => x"38",
          4947 => x"75",
          4948 => x"17",
          4949 => x"75",
          4950 => x"30",
          4951 => x"51",
          4952 => x"80",
          4953 => x"38",
          4954 => x"87",
          4955 => x"26",
          4956 => x"77",
          4957 => x"a4",
          4958 => x"27",
          4959 => x"a0",
          4960 => x"39",
          4961 => x"33",
          4962 => x"57",
          4963 => x"27",
          4964 => x"75",
          4965 => x"30",
          4966 => x"32",
          4967 => x"80",
          4968 => x"25",
          4969 => x"56",
          4970 => x"80",
          4971 => x"84",
          4972 => x"58",
          4973 => x"70",
          4974 => x"55",
          4975 => x"09",
          4976 => x"38",
          4977 => x"80",
          4978 => x"30",
          4979 => x"77",
          4980 => x"54",
          4981 => x"81",
          4982 => x"ae",
          4983 => x"06",
          4984 => x"54",
          4985 => x"74",
          4986 => x"80",
          4987 => x"7b",
          4988 => x"30",
          4989 => x"70",
          4990 => x"25",
          4991 => x"07",
          4992 => x"51",
          4993 => x"a7",
          4994 => x"8b",
          4995 => x"39",
          4996 => x"54",
          4997 => x"8c",
          4998 => x"ff",
          4999 => x"94",
          5000 => x"54",
          5001 => x"e1",
          5002 => x"cc",
          5003 => x"b2",
          5004 => x"70",
          5005 => x"71",
          5006 => x"54",
          5007 => x"82",
          5008 => x"80",
          5009 => x"38",
          5010 => x"76",
          5011 => x"df",
          5012 => x"54",
          5013 => x"81",
          5014 => x"55",
          5015 => x"34",
          5016 => x"52",
          5017 => x"51",
          5018 => x"82",
          5019 => x"bf",
          5020 => x"16",
          5021 => x"26",
          5022 => x"16",
          5023 => x"06",
          5024 => x"17",
          5025 => x"34",
          5026 => x"fd",
          5027 => x"19",
          5028 => x"80",
          5029 => x"79",
          5030 => x"81",
          5031 => x"81",
          5032 => x"85",
          5033 => x"54",
          5034 => x"8f",
          5035 => x"86",
          5036 => x"39",
          5037 => x"f3",
          5038 => x"73",
          5039 => x"80",
          5040 => x"52",
          5041 => x"ce",
          5042 => x"cc",
          5043 => x"87",
          5044 => x"d7",
          5045 => x"08",
          5046 => x"e6",
          5047 => x"87",
          5048 => x"82",
          5049 => x"80",
          5050 => x"1b",
          5051 => x"55",
          5052 => x"2e",
          5053 => x"8b",
          5054 => x"06",
          5055 => x"1c",
          5056 => x"33",
          5057 => x"70",
          5058 => x"55",
          5059 => x"38",
          5060 => x"52",
          5061 => x"9f",
          5062 => x"cc",
          5063 => x"8b",
          5064 => x"7a",
          5065 => x"3f",
          5066 => x"75",
          5067 => x"57",
          5068 => x"2e",
          5069 => x"84",
          5070 => x"06",
          5071 => x"75",
          5072 => x"81",
          5073 => x"2a",
          5074 => x"73",
          5075 => x"38",
          5076 => x"54",
          5077 => x"fb",
          5078 => x"80",
          5079 => x"34",
          5080 => x"c1",
          5081 => x"06",
          5082 => x"38",
          5083 => x"39",
          5084 => x"70",
          5085 => x"54",
          5086 => x"86",
          5087 => x"84",
          5088 => x"06",
          5089 => x"73",
          5090 => x"38",
          5091 => x"83",
          5092 => x"b4",
          5093 => x"51",
          5094 => x"82",
          5095 => x"88",
          5096 => x"ea",
          5097 => x"87",
          5098 => x"3d",
          5099 => x"3d",
          5100 => x"ff",
          5101 => x"71",
          5102 => x"5c",
          5103 => x"80",
          5104 => x"38",
          5105 => x"05",
          5106 => x"a0",
          5107 => x"71",
          5108 => x"38",
          5109 => x"71",
          5110 => x"81",
          5111 => x"38",
          5112 => x"11",
          5113 => x"06",
          5114 => x"70",
          5115 => x"38",
          5116 => x"81",
          5117 => x"05",
          5118 => x"76",
          5119 => x"38",
          5120 => x"81",
          5121 => x"77",
          5122 => x"57",
          5123 => x"05",
          5124 => x"70",
          5125 => x"33",
          5126 => x"53",
          5127 => x"99",
          5128 => x"e0",
          5129 => x"ff",
          5130 => x"ff",
          5131 => x"70",
          5132 => x"38",
          5133 => x"81",
          5134 => x"51",
          5135 => x"9f",
          5136 => x"72",
          5137 => x"81",
          5138 => x"70",
          5139 => x"72",
          5140 => x"32",
          5141 => x"72",
          5142 => x"73",
          5143 => x"53",
          5144 => x"70",
          5145 => x"38",
          5146 => x"19",
          5147 => x"75",
          5148 => x"38",
          5149 => x"83",
          5150 => x"74",
          5151 => x"59",
          5152 => x"39",
          5153 => x"33",
          5154 => x"87",
          5155 => x"3d",
          5156 => x"3d",
          5157 => x"80",
          5158 => x"34",
          5159 => x"17",
          5160 => x"75",
          5161 => x"3f",
          5162 => x"87",
          5163 => x"80",
          5164 => x"16",
          5165 => x"3f",
          5166 => x"08",
          5167 => x"06",
          5168 => x"73",
          5169 => x"2e",
          5170 => x"80",
          5171 => x"0b",
          5172 => x"56",
          5173 => x"e9",
          5174 => x"06",
          5175 => x"57",
          5176 => x"32",
          5177 => x"80",
          5178 => x"51",
          5179 => x"8a",
          5180 => x"e8",
          5181 => x"06",
          5182 => x"53",
          5183 => x"52",
          5184 => x"51",
          5185 => x"82",
          5186 => x"55",
          5187 => x"08",
          5188 => x"38",
          5189 => x"80",
          5190 => x"86",
          5191 => x"97",
          5192 => x"cc",
          5193 => x"87",
          5194 => x"2e",
          5195 => x"55",
          5196 => x"cc",
          5197 => x"0d",
          5198 => x"0d",
          5199 => x"05",
          5200 => x"33",
          5201 => x"75",
          5202 => x"fc",
          5203 => x"87",
          5204 => x"8b",
          5205 => x"82",
          5206 => x"24",
          5207 => x"82",
          5208 => x"84",
          5209 => x"f0",
          5210 => x"55",
          5211 => x"73",
          5212 => x"e5",
          5213 => x"0c",
          5214 => x"06",
          5215 => x"57",
          5216 => x"ae",
          5217 => x"33",
          5218 => x"3f",
          5219 => x"08",
          5220 => x"70",
          5221 => x"55",
          5222 => x"76",
          5223 => x"b7",
          5224 => x"2a",
          5225 => x"51",
          5226 => x"72",
          5227 => x"86",
          5228 => x"74",
          5229 => x"15",
          5230 => x"81",
          5231 => x"d7",
          5232 => x"87",
          5233 => x"ff",
          5234 => x"06",
          5235 => x"56",
          5236 => x"38",
          5237 => x"8f",
          5238 => x"2a",
          5239 => x"51",
          5240 => x"72",
          5241 => x"80",
          5242 => x"52",
          5243 => x"3f",
          5244 => x"08",
          5245 => x"57",
          5246 => x"09",
          5247 => x"e2",
          5248 => x"74",
          5249 => x"56",
          5250 => x"33",
          5251 => x"72",
          5252 => x"38",
          5253 => x"51",
          5254 => x"82",
          5255 => x"57",
          5256 => x"84",
          5257 => x"ff",
          5258 => x"56",
          5259 => x"25",
          5260 => x"0b",
          5261 => x"56",
          5262 => x"05",
          5263 => x"83",
          5264 => x"2e",
          5265 => x"52",
          5266 => x"c6",
          5267 => x"cc",
          5268 => x"06",
          5269 => x"27",
          5270 => x"16",
          5271 => x"27",
          5272 => x"56",
          5273 => x"84",
          5274 => x"56",
          5275 => x"84",
          5276 => x"14",
          5277 => x"3f",
          5278 => x"08",
          5279 => x"06",
          5280 => x"80",
          5281 => x"06",
          5282 => x"80",
          5283 => x"db",
          5284 => x"87",
          5285 => x"ff",
          5286 => x"77",
          5287 => x"d8",
          5288 => x"de",
          5289 => x"cc",
          5290 => x"9c",
          5291 => x"c4",
          5292 => x"15",
          5293 => x"14",
          5294 => x"70",
          5295 => x"51",
          5296 => x"56",
          5297 => x"84",
          5298 => x"81",
          5299 => x"71",
          5300 => x"16",
          5301 => x"53",
          5302 => x"23",
          5303 => x"8b",
          5304 => x"73",
          5305 => x"80",
          5306 => x"8d",
          5307 => x"39",
          5308 => x"51",
          5309 => x"82",
          5310 => x"53",
          5311 => x"08",
          5312 => x"72",
          5313 => x"8d",
          5314 => x"cd",
          5315 => x"14",
          5316 => x"3f",
          5317 => x"08",
          5318 => x"06",
          5319 => x"38",
          5320 => x"51",
          5321 => x"82",
          5322 => x"55",
          5323 => x"51",
          5324 => x"82",
          5325 => x"83",
          5326 => x"53",
          5327 => x"80",
          5328 => x"38",
          5329 => x"78",
          5330 => x"2a",
          5331 => x"78",
          5332 => x"85",
          5333 => x"22",
          5334 => x"31",
          5335 => x"3f",
          5336 => x"08",
          5337 => x"cc",
          5338 => x"82",
          5339 => x"87",
          5340 => x"ff",
          5341 => x"26",
          5342 => x"57",
          5343 => x"f5",
          5344 => x"82",
          5345 => x"f5",
          5346 => x"81",
          5347 => x"8d",
          5348 => x"2e",
          5349 => x"82",
          5350 => x"16",
          5351 => x"16",
          5352 => x"70",
          5353 => x"7a",
          5354 => x"0c",
          5355 => x"83",
          5356 => x"06",
          5357 => x"de",
          5358 => x"af",
          5359 => x"cc",
          5360 => x"ff",
          5361 => x"56",
          5362 => x"38",
          5363 => x"38",
          5364 => x"51",
          5365 => x"82",
          5366 => x"a8",
          5367 => x"82",
          5368 => x"39",
          5369 => x"80",
          5370 => x"38",
          5371 => x"15",
          5372 => x"53",
          5373 => x"8d",
          5374 => x"15",
          5375 => x"76",
          5376 => x"51",
          5377 => x"13",
          5378 => x"8d",
          5379 => x"15",
          5380 => x"c5",
          5381 => x"90",
          5382 => x"0b",
          5383 => x"ff",
          5384 => x"15",
          5385 => x"2e",
          5386 => x"81",
          5387 => x"e4",
          5388 => x"b7",
          5389 => x"cc",
          5390 => x"ff",
          5391 => x"81",
          5392 => x"06",
          5393 => x"81",
          5394 => x"51",
          5395 => x"82",
          5396 => x"80",
          5397 => x"87",
          5398 => x"15",
          5399 => x"14",
          5400 => x"3f",
          5401 => x"08",
          5402 => x"06",
          5403 => x"d4",
          5404 => x"81",
          5405 => x"38",
          5406 => x"d8",
          5407 => x"87",
          5408 => x"8b",
          5409 => x"2e",
          5410 => x"b3",
          5411 => x"14",
          5412 => x"3f",
          5413 => x"08",
          5414 => x"e4",
          5415 => x"81",
          5416 => x"84",
          5417 => x"d7",
          5418 => x"87",
          5419 => x"15",
          5420 => x"14",
          5421 => x"3f",
          5422 => x"08",
          5423 => x"76",
          5424 => x"9f",
          5425 => x"05",
          5426 => x"9f",
          5427 => x"86",
          5428 => x"0b",
          5429 => x"80",
          5430 => x"87",
          5431 => x"3d",
          5432 => x"3d",
          5433 => x"89",
          5434 => x"2e",
          5435 => x"08",
          5436 => x"2e",
          5437 => x"33",
          5438 => x"2e",
          5439 => x"13",
          5440 => x"22",
          5441 => x"76",
          5442 => x"06",
          5443 => x"13",
          5444 => x"c1",
          5445 => x"cc",
          5446 => x"52",
          5447 => x"71",
          5448 => x"55",
          5449 => x"53",
          5450 => x"0c",
          5451 => x"87",
          5452 => x"3d",
          5453 => x"3d",
          5454 => x"05",
          5455 => x"89",
          5456 => x"52",
          5457 => x"3f",
          5458 => x"0b",
          5459 => x"08",
          5460 => x"82",
          5461 => x"84",
          5462 => x"f0",
          5463 => x"55",
          5464 => x"2e",
          5465 => x"74",
          5466 => x"73",
          5467 => x"38",
          5468 => x"78",
          5469 => x"54",
          5470 => x"92",
          5471 => x"89",
          5472 => x"84",
          5473 => x"b1",
          5474 => x"cc",
          5475 => x"82",
          5476 => x"88",
          5477 => x"eb",
          5478 => x"02",
          5479 => x"e7",
          5480 => x"59",
          5481 => x"80",
          5482 => x"38",
          5483 => x"70",
          5484 => x"d0",
          5485 => x"3d",
          5486 => x"58",
          5487 => x"82",
          5488 => x"55",
          5489 => x"08",
          5490 => x"7a",
          5491 => x"8c",
          5492 => x"56",
          5493 => x"82",
          5494 => x"55",
          5495 => x"08",
          5496 => x"80",
          5497 => x"70",
          5498 => x"57",
          5499 => x"83",
          5500 => x"77",
          5501 => x"73",
          5502 => x"ab",
          5503 => x"2e",
          5504 => x"84",
          5505 => x"06",
          5506 => x"51",
          5507 => x"82",
          5508 => x"55",
          5509 => x"b2",
          5510 => x"06",
          5511 => x"b8",
          5512 => x"2a",
          5513 => x"51",
          5514 => x"2e",
          5515 => x"55",
          5516 => x"77",
          5517 => x"74",
          5518 => x"77",
          5519 => x"81",
          5520 => x"73",
          5521 => x"af",
          5522 => x"7a",
          5523 => x"3f",
          5524 => x"08",
          5525 => x"b2",
          5526 => x"8e",
          5527 => x"eb",
          5528 => x"a0",
          5529 => x"34",
          5530 => x"52",
          5531 => x"be",
          5532 => x"62",
          5533 => x"d4",
          5534 => x"54",
          5535 => x"15",
          5536 => x"2e",
          5537 => x"7a",
          5538 => x"51",
          5539 => x"75",
          5540 => x"d4",
          5541 => x"bf",
          5542 => x"cc",
          5543 => x"87",
          5544 => x"ca",
          5545 => x"74",
          5546 => x"02",
          5547 => x"70",
          5548 => x"81",
          5549 => x"56",
          5550 => x"86",
          5551 => x"82",
          5552 => x"81",
          5553 => x"06",
          5554 => x"80",
          5555 => x"75",
          5556 => x"73",
          5557 => x"38",
          5558 => x"92",
          5559 => x"7a",
          5560 => x"3f",
          5561 => x"08",
          5562 => x"8c",
          5563 => x"55",
          5564 => x"08",
          5565 => x"77",
          5566 => x"81",
          5567 => x"73",
          5568 => x"38",
          5569 => x"07",
          5570 => x"11",
          5571 => x"0c",
          5572 => x"0c",
          5573 => x"52",
          5574 => x"3f",
          5575 => x"08",
          5576 => x"08",
          5577 => x"63",
          5578 => x"5a",
          5579 => x"82",
          5580 => x"82",
          5581 => x"8c",
          5582 => x"7a",
          5583 => x"17",
          5584 => x"23",
          5585 => x"34",
          5586 => x"1a",
          5587 => x"9c",
          5588 => x"0b",
          5589 => x"77",
          5590 => x"81",
          5591 => x"73",
          5592 => x"8d",
          5593 => x"cc",
          5594 => x"81",
          5595 => x"87",
          5596 => x"1a",
          5597 => x"22",
          5598 => x"7b",
          5599 => x"a8",
          5600 => x"78",
          5601 => x"3f",
          5602 => x"08",
          5603 => x"cc",
          5604 => x"83",
          5605 => x"82",
          5606 => x"ff",
          5607 => x"06",
          5608 => x"55",
          5609 => x"56",
          5610 => x"76",
          5611 => x"51",
          5612 => x"27",
          5613 => x"70",
          5614 => x"5a",
          5615 => x"76",
          5616 => x"74",
          5617 => x"83",
          5618 => x"73",
          5619 => x"38",
          5620 => x"51",
          5621 => x"82",
          5622 => x"85",
          5623 => x"8e",
          5624 => x"2a",
          5625 => x"08",
          5626 => x"0c",
          5627 => x"79",
          5628 => x"73",
          5629 => x"0c",
          5630 => x"04",
          5631 => x"60",
          5632 => x"40",
          5633 => x"80",
          5634 => x"3d",
          5635 => x"78",
          5636 => x"3f",
          5637 => x"08",
          5638 => x"cc",
          5639 => x"91",
          5640 => x"74",
          5641 => x"38",
          5642 => x"c4",
          5643 => x"33",
          5644 => x"87",
          5645 => x"2e",
          5646 => x"95",
          5647 => x"91",
          5648 => x"56",
          5649 => x"81",
          5650 => x"34",
          5651 => x"a0",
          5652 => x"08",
          5653 => x"31",
          5654 => x"27",
          5655 => x"5c",
          5656 => x"82",
          5657 => x"19",
          5658 => x"ff",
          5659 => x"74",
          5660 => x"7e",
          5661 => x"ff",
          5662 => x"2a",
          5663 => x"79",
          5664 => x"87",
          5665 => x"08",
          5666 => x"98",
          5667 => x"78",
          5668 => x"3f",
          5669 => x"08",
          5670 => x"27",
          5671 => x"74",
          5672 => x"a3",
          5673 => x"1a",
          5674 => x"08",
          5675 => x"d4",
          5676 => x"87",
          5677 => x"2e",
          5678 => x"82",
          5679 => x"1a",
          5680 => x"59",
          5681 => x"2e",
          5682 => x"77",
          5683 => x"11",
          5684 => x"55",
          5685 => x"85",
          5686 => x"31",
          5687 => x"76",
          5688 => x"81",
          5689 => x"ca",
          5690 => x"87",
          5691 => x"d7",
          5692 => x"11",
          5693 => x"74",
          5694 => x"38",
          5695 => x"77",
          5696 => x"78",
          5697 => x"84",
          5698 => x"16",
          5699 => x"08",
          5700 => x"2b",
          5701 => x"cf",
          5702 => x"89",
          5703 => x"39",
          5704 => x"0c",
          5705 => x"83",
          5706 => x"80",
          5707 => x"55",
          5708 => x"83",
          5709 => x"9c",
          5710 => x"7e",
          5711 => x"3f",
          5712 => x"08",
          5713 => x"75",
          5714 => x"08",
          5715 => x"1f",
          5716 => x"7c",
          5717 => x"3f",
          5718 => x"7e",
          5719 => x"0c",
          5720 => x"1b",
          5721 => x"1c",
          5722 => x"fd",
          5723 => x"56",
          5724 => x"cc",
          5725 => x"0d",
          5726 => x"0d",
          5727 => x"64",
          5728 => x"58",
          5729 => x"90",
          5730 => x"52",
          5731 => x"d2",
          5732 => x"cc",
          5733 => x"87",
          5734 => x"38",
          5735 => x"55",
          5736 => x"86",
          5737 => x"83",
          5738 => x"18",
          5739 => x"2a",
          5740 => x"51",
          5741 => x"56",
          5742 => x"83",
          5743 => x"39",
          5744 => x"19",
          5745 => x"83",
          5746 => x"0b",
          5747 => x"81",
          5748 => x"39",
          5749 => x"7c",
          5750 => x"74",
          5751 => x"38",
          5752 => x"7b",
          5753 => x"ec",
          5754 => x"08",
          5755 => x"06",
          5756 => x"81",
          5757 => x"8a",
          5758 => x"05",
          5759 => x"06",
          5760 => x"bf",
          5761 => x"38",
          5762 => x"55",
          5763 => x"7a",
          5764 => x"98",
          5765 => x"77",
          5766 => x"3f",
          5767 => x"08",
          5768 => x"cc",
          5769 => x"82",
          5770 => x"81",
          5771 => x"38",
          5772 => x"ff",
          5773 => x"98",
          5774 => x"18",
          5775 => x"74",
          5776 => x"7e",
          5777 => x"08",
          5778 => x"2e",
          5779 => x"8d",
          5780 => x"ce",
          5781 => x"87",
          5782 => x"ee",
          5783 => x"08",
          5784 => x"d1",
          5785 => x"87",
          5786 => x"2e",
          5787 => x"82",
          5788 => x"1b",
          5789 => x"5a",
          5790 => x"2e",
          5791 => x"78",
          5792 => x"11",
          5793 => x"55",
          5794 => x"85",
          5795 => x"31",
          5796 => x"76",
          5797 => x"81",
          5798 => x"c8",
          5799 => x"87",
          5800 => x"a6",
          5801 => x"11",
          5802 => x"56",
          5803 => x"27",
          5804 => x"80",
          5805 => x"08",
          5806 => x"2b",
          5807 => x"b4",
          5808 => x"b6",
          5809 => x"80",
          5810 => x"34",
          5811 => x"56",
          5812 => x"8c",
          5813 => x"19",
          5814 => x"38",
          5815 => x"b7",
          5816 => x"cc",
          5817 => x"38",
          5818 => x"12",
          5819 => x"9c",
          5820 => x"18",
          5821 => x"06",
          5822 => x"31",
          5823 => x"76",
          5824 => x"7b",
          5825 => x"08",
          5826 => x"cd",
          5827 => x"87",
          5828 => x"b6",
          5829 => x"7c",
          5830 => x"08",
          5831 => x"1f",
          5832 => x"cb",
          5833 => x"55",
          5834 => x"16",
          5835 => x"31",
          5836 => x"7f",
          5837 => x"94",
          5838 => x"70",
          5839 => x"8c",
          5840 => x"58",
          5841 => x"76",
          5842 => x"75",
          5843 => x"19",
          5844 => x"39",
          5845 => x"80",
          5846 => x"74",
          5847 => x"80",
          5848 => x"87",
          5849 => x"3d",
          5850 => x"3d",
          5851 => x"3d",
          5852 => x"70",
          5853 => x"ea",
          5854 => x"cc",
          5855 => x"87",
          5856 => x"fb",
          5857 => x"33",
          5858 => x"70",
          5859 => x"55",
          5860 => x"2e",
          5861 => x"a0",
          5862 => x"78",
          5863 => x"3f",
          5864 => x"08",
          5865 => x"cc",
          5866 => x"38",
          5867 => x"8b",
          5868 => x"07",
          5869 => x"8b",
          5870 => x"16",
          5871 => x"52",
          5872 => x"dd",
          5873 => x"16",
          5874 => x"15",
          5875 => x"3f",
          5876 => x"0a",
          5877 => x"51",
          5878 => x"76",
          5879 => x"51",
          5880 => x"78",
          5881 => x"83",
          5882 => x"51",
          5883 => x"82",
          5884 => x"90",
          5885 => x"bf",
          5886 => x"73",
          5887 => x"76",
          5888 => x"0c",
          5889 => x"04",
          5890 => x"76",
          5891 => x"fe",
          5892 => x"87",
          5893 => x"82",
          5894 => x"9c",
          5895 => x"fc",
          5896 => x"51",
          5897 => x"82",
          5898 => x"53",
          5899 => x"08",
          5900 => x"87",
          5901 => x"0c",
          5902 => x"cc",
          5903 => x"0d",
          5904 => x"0d",
          5905 => x"e6",
          5906 => x"52",
          5907 => x"87",
          5908 => x"8b",
          5909 => x"cc",
          5910 => x"84",
          5911 => x"71",
          5912 => x"0c",
          5913 => x"04",
          5914 => x"80",
          5915 => x"d0",
          5916 => x"3d",
          5917 => x"3f",
          5918 => x"08",
          5919 => x"cc",
          5920 => x"38",
          5921 => x"52",
          5922 => x"05",
          5923 => x"3f",
          5924 => x"08",
          5925 => x"cc",
          5926 => x"02",
          5927 => x"33",
          5928 => x"55",
          5929 => x"25",
          5930 => x"7a",
          5931 => x"54",
          5932 => x"a2",
          5933 => x"84",
          5934 => x"06",
          5935 => x"73",
          5936 => x"38",
          5937 => x"70",
          5938 => x"a9",
          5939 => x"cc",
          5940 => x"0c",
          5941 => x"87",
          5942 => x"2e",
          5943 => x"83",
          5944 => x"74",
          5945 => x"0c",
          5946 => x"04",
          5947 => x"6f",
          5948 => x"80",
          5949 => x"53",
          5950 => x"b8",
          5951 => x"3d",
          5952 => x"3f",
          5953 => x"08",
          5954 => x"cc",
          5955 => x"38",
          5956 => x"7c",
          5957 => x"47",
          5958 => x"54",
          5959 => x"81",
          5960 => x"52",
          5961 => x"52",
          5962 => x"3f",
          5963 => x"08",
          5964 => x"cc",
          5965 => x"38",
          5966 => x"51",
          5967 => x"82",
          5968 => x"57",
          5969 => x"08",
          5970 => x"69",
          5971 => x"da",
          5972 => x"87",
          5973 => x"76",
          5974 => x"d5",
          5975 => x"87",
          5976 => x"82",
          5977 => x"82",
          5978 => x"52",
          5979 => x"ec",
          5980 => x"cc",
          5981 => x"87",
          5982 => x"38",
          5983 => x"51",
          5984 => x"73",
          5985 => x"08",
          5986 => x"76",
          5987 => x"d6",
          5988 => x"87",
          5989 => x"82",
          5990 => x"80",
          5991 => x"76",
          5992 => x"81",
          5993 => x"82",
          5994 => x"39",
          5995 => x"38",
          5996 => x"bc",
          5997 => x"51",
          5998 => x"76",
          5999 => x"11",
          6000 => x"51",
          6001 => x"73",
          6002 => x"38",
          6003 => x"55",
          6004 => x"16",
          6005 => x"56",
          6006 => x"38",
          6007 => x"73",
          6008 => x"90",
          6009 => x"2e",
          6010 => x"16",
          6011 => x"ff",
          6012 => x"ff",
          6013 => x"58",
          6014 => x"74",
          6015 => x"75",
          6016 => x"18",
          6017 => x"58",
          6018 => x"fe",
          6019 => x"7b",
          6020 => x"06",
          6021 => x"18",
          6022 => x"58",
          6023 => x"80",
          6024 => x"84",
          6025 => x"29",
          6026 => x"05",
          6027 => x"33",
          6028 => x"56",
          6029 => x"2e",
          6030 => x"16",
          6031 => x"33",
          6032 => x"73",
          6033 => x"16",
          6034 => x"26",
          6035 => x"55",
          6036 => x"91",
          6037 => x"54",
          6038 => x"70",
          6039 => x"34",
          6040 => x"ec",
          6041 => x"70",
          6042 => x"34",
          6043 => x"09",
          6044 => x"38",
          6045 => x"39",
          6046 => x"19",
          6047 => x"33",
          6048 => x"05",
          6049 => x"78",
          6050 => x"80",
          6051 => x"82",
          6052 => x"9e",
          6053 => x"f7",
          6054 => x"7d",
          6055 => x"05",
          6056 => x"57",
          6057 => x"3f",
          6058 => x"08",
          6059 => x"cc",
          6060 => x"38",
          6061 => x"53",
          6062 => x"38",
          6063 => x"54",
          6064 => x"92",
          6065 => x"33",
          6066 => x"70",
          6067 => x"54",
          6068 => x"38",
          6069 => x"15",
          6070 => x"70",
          6071 => x"58",
          6072 => x"82",
          6073 => x"8a",
          6074 => x"89",
          6075 => x"53",
          6076 => x"b7",
          6077 => x"ff",
          6078 => x"ad",
          6079 => x"87",
          6080 => x"15",
          6081 => x"53",
          6082 => x"ad",
          6083 => x"87",
          6084 => x"26",
          6085 => x"30",
          6086 => x"70",
          6087 => x"77",
          6088 => x"18",
          6089 => x"51",
          6090 => x"88",
          6091 => x"73",
          6092 => x"52",
          6093 => x"cb",
          6094 => x"cc",
          6095 => x"87",
          6096 => x"2e",
          6097 => x"82",
          6098 => x"ff",
          6099 => x"38",
          6100 => x"08",
          6101 => x"73",
          6102 => x"73",
          6103 => x"9c",
          6104 => x"27",
          6105 => x"75",
          6106 => x"16",
          6107 => x"17",
          6108 => x"33",
          6109 => x"70",
          6110 => x"55",
          6111 => x"80",
          6112 => x"73",
          6113 => x"cc",
          6114 => x"87",
          6115 => x"82",
          6116 => x"94",
          6117 => x"cc",
          6118 => x"39",
          6119 => x"51",
          6120 => x"82",
          6121 => x"54",
          6122 => x"be",
          6123 => x"27",
          6124 => x"53",
          6125 => x"08",
          6126 => x"73",
          6127 => x"ff",
          6128 => x"15",
          6129 => x"16",
          6130 => x"ff",
          6131 => x"80",
          6132 => x"73",
          6133 => x"c6",
          6134 => x"87",
          6135 => x"38",
          6136 => x"16",
          6137 => x"80",
          6138 => x"0b",
          6139 => x"81",
          6140 => x"75",
          6141 => x"87",
          6142 => x"58",
          6143 => x"54",
          6144 => x"74",
          6145 => x"73",
          6146 => x"90",
          6147 => x"c0",
          6148 => x"90",
          6149 => x"83",
          6150 => x"72",
          6151 => x"38",
          6152 => x"08",
          6153 => x"77",
          6154 => x"80",
          6155 => x"87",
          6156 => x"3d",
          6157 => x"3d",
          6158 => x"89",
          6159 => x"2e",
          6160 => x"80",
          6161 => x"fc",
          6162 => x"3d",
          6163 => x"e1",
          6164 => x"87",
          6165 => x"82",
          6166 => x"80",
          6167 => x"76",
          6168 => x"75",
          6169 => x"3f",
          6170 => x"08",
          6171 => x"cc",
          6172 => x"38",
          6173 => x"70",
          6174 => x"57",
          6175 => x"a2",
          6176 => x"33",
          6177 => x"70",
          6178 => x"55",
          6179 => x"2e",
          6180 => x"16",
          6181 => x"51",
          6182 => x"82",
          6183 => x"88",
          6184 => x"54",
          6185 => x"84",
          6186 => x"52",
          6187 => x"e6",
          6188 => x"cc",
          6189 => x"84",
          6190 => x"06",
          6191 => x"55",
          6192 => x"80",
          6193 => x"80",
          6194 => x"54",
          6195 => x"cc",
          6196 => x"0d",
          6197 => x"0d",
          6198 => x"fc",
          6199 => x"52",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"87",
          6203 => x"0c",
          6204 => x"04",
          6205 => x"77",
          6206 => x"fc",
          6207 => x"53",
          6208 => x"de",
          6209 => x"cc",
          6210 => x"87",
          6211 => x"df",
          6212 => x"38",
          6213 => x"08",
          6214 => x"cd",
          6215 => x"87",
          6216 => x"80",
          6217 => x"87",
          6218 => x"73",
          6219 => x"3f",
          6220 => x"08",
          6221 => x"cc",
          6222 => x"09",
          6223 => x"38",
          6224 => x"39",
          6225 => x"08",
          6226 => x"52",
          6227 => x"b4",
          6228 => x"73",
          6229 => x"3f",
          6230 => x"08",
          6231 => x"30",
          6232 => x"9f",
          6233 => x"87",
          6234 => x"51",
          6235 => x"72",
          6236 => x"0c",
          6237 => x"04",
          6238 => x"65",
          6239 => x"89",
          6240 => x"96",
          6241 => x"df",
          6242 => x"87",
          6243 => x"82",
          6244 => x"b2",
          6245 => x"75",
          6246 => x"3f",
          6247 => x"08",
          6248 => x"cc",
          6249 => x"02",
          6250 => x"33",
          6251 => x"55",
          6252 => x"25",
          6253 => x"55",
          6254 => x"80",
          6255 => x"76",
          6256 => x"d4",
          6257 => x"82",
          6258 => x"94",
          6259 => x"f0",
          6260 => x"65",
          6261 => x"53",
          6262 => x"05",
          6263 => x"51",
          6264 => x"82",
          6265 => x"5b",
          6266 => x"08",
          6267 => x"7c",
          6268 => x"08",
          6269 => x"fe",
          6270 => x"08",
          6271 => x"55",
          6272 => x"91",
          6273 => x"0c",
          6274 => x"81",
          6275 => x"39",
          6276 => x"c7",
          6277 => x"cc",
          6278 => x"55",
          6279 => x"2e",
          6280 => x"bf",
          6281 => x"5f",
          6282 => x"92",
          6283 => x"51",
          6284 => x"82",
          6285 => x"ff",
          6286 => x"82",
          6287 => x"81",
          6288 => x"82",
          6289 => x"30",
          6290 => x"cc",
          6291 => x"25",
          6292 => x"19",
          6293 => x"5a",
          6294 => x"08",
          6295 => x"38",
          6296 => x"a4",
          6297 => x"87",
          6298 => x"58",
          6299 => x"77",
          6300 => x"7d",
          6301 => x"bf",
          6302 => x"87",
          6303 => x"82",
          6304 => x"80",
          6305 => x"70",
          6306 => x"ff",
          6307 => x"56",
          6308 => x"2e",
          6309 => x"9e",
          6310 => x"51",
          6311 => x"3f",
          6312 => x"08",
          6313 => x"06",
          6314 => x"80",
          6315 => x"19",
          6316 => x"54",
          6317 => x"14",
          6318 => x"c6",
          6319 => x"cc",
          6320 => x"06",
          6321 => x"80",
          6322 => x"19",
          6323 => x"54",
          6324 => x"06",
          6325 => x"79",
          6326 => x"78",
          6327 => x"79",
          6328 => x"84",
          6329 => x"07",
          6330 => x"84",
          6331 => x"82",
          6332 => x"92",
          6333 => x"f9",
          6334 => x"8a",
          6335 => x"53",
          6336 => x"e3",
          6337 => x"87",
          6338 => x"82",
          6339 => x"81",
          6340 => x"17",
          6341 => x"81",
          6342 => x"17",
          6343 => x"2a",
          6344 => x"51",
          6345 => x"55",
          6346 => x"81",
          6347 => x"17",
          6348 => x"8c",
          6349 => x"81",
          6350 => x"9b",
          6351 => x"cc",
          6352 => x"17",
          6353 => x"51",
          6354 => x"82",
          6355 => x"74",
          6356 => x"56",
          6357 => x"98",
          6358 => x"76",
          6359 => x"c7",
          6360 => x"cc",
          6361 => x"09",
          6362 => x"38",
          6363 => x"87",
          6364 => x"2e",
          6365 => x"85",
          6366 => x"a3",
          6367 => x"38",
          6368 => x"87",
          6369 => x"15",
          6370 => x"38",
          6371 => x"53",
          6372 => x"08",
          6373 => x"c3",
          6374 => x"87",
          6375 => x"94",
          6376 => x"18",
          6377 => x"33",
          6378 => x"54",
          6379 => x"34",
          6380 => x"85",
          6381 => x"18",
          6382 => x"74",
          6383 => x"0c",
          6384 => x"04",
          6385 => x"82",
          6386 => x"ff",
          6387 => x"a1",
          6388 => x"e5",
          6389 => x"cc",
          6390 => x"87",
          6391 => x"f5",
          6392 => x"a1",
          6393 => x"95",
          6394 => x"58",
          6395 => x"82",
          6396 => x"55",
          6397 => x"08",
          6398 => x"02",
          6399 => x"33",
          6400 => x"70",
          6401 => x"55",
          6402 => x"73",
          6403 => x"75",
          6404 => x"80",
          6405 => x"bd",
          6406 => x"d6",
          6407 => x"81",
          6408 => x"87",
          6409 => x"ad",
          6410 => x"78",
          6411 => x"3f",
          6412 => x"08",
          6413 => x"70",
          6414 => x"55",
          6415 => x"2e",
          6416 => x"78",
          6417 => x"cc",
          6418 => x"08",
          6419 => x"38",
          6420 => x"87",
          6421 => x"76",
          6422 => x"70",
          6423 => x"b6",
          6424 => x"cc",
          6425 => x"87",
          6426 => x"e9",
          6427 => x"cc",
          6428 => x"51",
          6429 => x"82",
          6430 => x"55",
          6431 => x"08",
          6432 => x"55",
          6433 => x"82",
          6434 => x"84",
          6435 => x"82",
          6436 => x"80",
          6437 => x"51",
          6438 => x"82",
          6439 => x"82",
          6440 => x"30",
          6441 => x"cc",
          6442 => x"25",
          6443 => x"75",
          6444 => x"38",
          6445 => x"8f",
          6446 => x"75",
          6447 => x"c1",
          6448 => x"87",
          6449 => x"74",
          6450 => x"51",
          6451 => x"3f",
          6452 => x"08",
          6453 => x"87",
          6454 => x"3d",
          6455 => x"3d",
          6456 => x"99",
          6457 => x"52",
          6458 => x"d8",
          6459 => x"87",
          6460 => x"82",
          6461 => x"82",
          6462 => x"5e",
          6463 => x"3d",
          6464 => x"cf",
          6465 => x"87",
          6466 => x"82",
          6467 => x"86",
          6468 => x"82",
          6469 => x"87",
          6470 => x"2e",
          6471 => x"82",
          6472 => x"80",
          6473 => x"70",
          6474 => x"06",
          6475 => x"54",
          6476 => x"38",
          6477 => x"52",
          6478 => x"52",
          6479 => x"3f",
          6480 => x"08",
          6481 => x"82",
          6482 => x"83",
          6483 => x"82",
          6484 => x"81",
          6485 => x"06",
          6486 => x"54",
          6487 => x"08",
          6488 => x"81",
          6489 => x"81",
          6490 => x"39",
          6491 => x"38",
          6492 => x"08",
          6493 => x"c4",
          6494 => x"87",
          6495 => x"82",
          6496 => x"81",
          6497 => x"53",
          6498 => x"19",
          6499 => x"8d",
          6500 => x"ae",
          6501 => x"34",
          6502 => x"0b",
          6503 => x"82",
          6504 => x"52",
          6505 => x"51",
          6506 => x"3f",
          6507 => x"b4",
          6508 => x"c9",
          6509 => x"53",
          6510 => x"53",
          6511 => x"51",
          6512 => x"3f",
          6513 => x"0b",
          6514 => x"34",
          6515 => x"80",
          6516 => x"51",
          6517 => x"78",
          6518 => x"83",
          6519 => x"51",
          6520 => x"82",
          6521 => x"54",
          6522 => x"08",
          6523 => x"88",
          6524 => x"64",
          6525 => x"ff",
          6526 => x"75",
          6527 => x"78",
          6528 => x"3f",
          6529 => x"0b",
          6530 => x"78",
          6531 => x"83",
          6532 => x"51",
          6533 => x"3f",
          6534 => x"08",
          6535 => x"80",
          6536 => x"76",
          6537 => x"af",
          6538 => x"87",
          6539 => x"3d",
          6540 => x"3d",
          6541 => x"84",
          6542 => x"f2",
          6543 => x"a8",
          6544 => x"05",
          6545 => x"51",
          6546 => x"82",
          6547 => x"55",
          6548 => x"08",
          6549 => x"78",
          6550 => x"08",
          6551 => x"70",
          6552 => x"b9",
          6553 => x"cc",
          6554 => x"87",
          6555 => x"b9",
          6556 => x"9b",
          6557 => x"a0",
          6558 => x"55",
          6559 => x"38",
          6560 => x"3d",
          6561 => x"3d",
          6562 => x"51",
          6563 => x"3f",
          6564 => x"52",
          6565 => x"52",
          6566 => x"de",
          6567 => x"08",
          6568 => x"cb",
          6569 => x"87",
          6570 => x"82",
          6571 => x"95",
          6572 => x"2e",
          6573 => x"88",
          6574 => x"3d",
          6575 => x"38",
          6576 => x"e5",
          6577 => x"cc",
          6578 => x"09",
          6579 => x"b8",
          6580 => x"c9",
          6581 => x"87",
          6582 => x"82",
          6583 => x"81",
          6584 => x"56",
          6585 => x"3d",
          6586 => x"52",
          6587 => x"ff",
          6588 => x"02",
          6589 => x"8b",
          6590 => x"16",
          6591 => x"2a",
          6592 => x"51",
          6593 => x"89",
          6594 => x"07",
          6595 => x"17",
          6596 => x"81",
          6597 => x"34",
          6598 => x"70",
          6599 => x"81",
          6600 => x"55",
          6601 => x"80",
          6602 => x"64",
          6603 => x"38",
          6604 => x"51",
          6605 => x"82",
          6606 => x"52",
          6607 => x"b7",
          6608 => x"55",
          6609 => x"08",
          6610 => x"dd",
          6611 => x"cc",
          6612 => x"51",
          6613 => x"3f",
          6614 => x"08",
          6615 => x"11",
          6616 => x"82",
          6617 => x"80",
          6618 => x"16",
          6619 => x"ae",
          6620 => x"06",
          6621 => x"53",
          6622 => x"51",
          6623 => x"78",
          6624 => x"83",
          6625 => x"39",
          6626 => x"08",
          6627 => x"51",
          6628 => x"82",
          6629 => x"55",
          6630 => x"08",
          6631 => x"51",
          6632 => x"3f",
          6633 => x"08",
          6634 => x"87",
          6635 => x"3d",
          6636 => x"3d",
          6637 => x"db",
          6638 => x"84",
          6639 => x"05",
          6640 => x"82",
          6641 => x"d0",
          6642 => x"3d",
          6643 => x"3f",
          6644 => x"08",
          6645 => x"cc",
          6646 => x"38",
          6647 => x"52",
          6648 => x"05",
          6649 => x"3f",
          6650 => x"08",
          6651 => x"cc",
          6652 => x"02",
          6653 => x"33",
          6654 => x"54",
          6655 => x"aa",
          6656 => x"06",
          6657 => x"8b",
          6658 => x"06",
          6659 => x"07",
          6660 => x"56",
          6661 => x"34",
          6662 => x"0b",
          6663 => x"78",
          6664 => x"aa",
          6665 => x"cc",
          6666 => x"82",
          6667 => x"95",
          6668 => x"ef",
          6669 => x"56",
          6670 => x"3d",
          6671 => x"94",
          6672 => x"f5",
          6673 => x"cc",
          6674 => x"87",
          6675 => x"cb",
          6676 => x"63",
          6677 => x"d4",
          6678 => x"c1",
          6679 => x"cc",
          6680 => x"87",
          6681 => x"38",
          6682 => x"05",
          6683 => x"06",
          6684 => x"73",
          6685 => x"16",
          6686 => x"22",
          6687 => x"07",
          6688 => x"1f",
          6689 => x"c3",
          6690 => x"81",
          6691 => x"34",
          6692 => x"b3",
          6693 => x"87",
          6694 => x"74",
          6695 => x"0c",
          6696 => x"04",
          6697 => x"69",
          6698 => x"80",
          6699 => x"d0",
          6700 => x"3d",
          6701 => x"3f",
          6702 => x"08",
          6703 => x"08",
          6704 => x"87",
          6705 => x"80",
          6706 => x"57",
          6707 => x"81",
          6708 => x"70",
          6709 => x"55",
          6710 => x"80",
          6711 => x"5d",
          6712 => x"52",
          6713 => x"52",
          6714 => x"aa",
          6715 => x"cc",
          6716 => x"87",
          6717 => x"d1",
          6718 => x"73",
          6719 => x"3f",
          6720 => x"08",
          6721 => x"cc",
          6722 => x"82",
          6723 => x"82",
          6724 => x"65",
          6725 => x"78",
          6726 => x"7b",
          6727 => x"55",
          6728 => x"34",
          6729 => x"8a",
          6730 => x"38",
          6731 => x"1a",
          6732 => x"34",
          6733 => x"9e",
          6734 => x"70",
          6735 => x"51",
          6736 => x"a0",
          6737 => x"8e",
          6738 => x"2e",
          6739 => x"86",
          6740 => x"34",
          6741 => x"30",
          6742 => x"80",
          6743 => x"7a",
          6744 => x"c1",
          6745 => x"2e",
          6746 => x"a0",
          6747 => x"51",
          6748 => x"3f",
          6749 => x"08",
          6750 => x"cc",
          6751 => x"7b",
          6752 => x"55",
          6753 => x"73",
          6754 => x"38",
          6755 => x"73",
          6756 => x"38",
          6757 => x"15",
          6758 => x"ff",
          6759 => x"82",
          6760 => x"7b",
          6761 => x"87",
          6762 => x"3d",
          6763 => x"3d",
          6764 => x"9c",
          6765 => x"05",
          6766 => x"51",
          6767 => x"82",
          6768 => x"82",
          6769 => x"56",
          6770 => x"cc",
          6771 => x"38",
          6772 => x"52",
          6773 => x"52",
          6774 => x"c1",
          6775 => x"70",
          6776 => x"ff",
          6777 => x"55",
          6778 => x"27",
          6779 => x"78",
          6780 => x"ff",
          6781 => x"05",
          6782 => x"55",
          6783 => x"3f",
          6784 => x"08",
          6785 => x"38",
          6786 => x"70",
          6787 => x"ff",
          6788 => x"82",
          6789 => x"80",
          6790 => x"74",
          6791 => x"07",
          6792 => x"4e",
          6793 => x"82",
          6794 => x"55",
          6795 => x"70",
          6796 => x"06",
          6797 => x"99",
          6798 => x"e0",
          6799 => x"ff",
          6800 => x"54",
          6801 => x"27",
          6802 => x"80",
          6803 => x"55",
          6804 => x"a3",
          6805 => x"82",
          6806 => x"ff",
          6807 => x"82",
          6808 => x"93",
          6809 => x"75",
          6810 => x"76",
          6811 => x"38",
          6812 => x"77",
          6813 => x"86",
          6814 => x"39",
          6815 => x"27",
          6816 => x"88",
          6817 => x"78",
          6818 => x"5a",
          6819 => x"57",
          6820 => x"81",
          6821 => x"81",
          6822 => x"33",
          6823 => x"06",
          6824 => x"57",
          6825 => x"fe",
          6826 => x"3d",
          6827 => x"55",
          6828 => x"2e",
          6829 => x"76",
          6830 => x"38",
          6831 => x"55",
          6832 => x"33",
          6833 => x"a0",
          6834 => x"06",
          6835 => x"17",
          6836 => x"38",
          6837 => x"43",
          6838 => x"3d",
          6839 => x"ff",
          6840 => x"82",
          6841 => x"54",
          6842 => x"08",
          6843 => x"81",
          6844 => x"ff",
          6845 => x"82",
          6846 => x"54",
          6847 => x"08",
          6848 => x"80",
          6849 => x"54",
          6850 => x"80",
          6851 => x"87",
          6852 => x"2e",
          6853 => x"80",
          6854 => x"54",
          6855 => x"80",
          6856 => x"52",
          6857 => x"bd",
          6858 => x"87",
          6859 => x"82",
          6860 => x"b1",
          6861 => x"82",
          6862 => x"52",
          6863 => x"ab",
          6864 => x"54",
          6865 => x"15",
          6866 => x"78",
          6867 => x"ff",
          6868 => x"79",
          6869 => x"83",
          6870 => x"51",
          6871 => x"3f",
          6872 => x"08",
          6873 => x"74",
          6874 => x"0c",
          6875 => x"04",
          6876 => x"60",
          6877 => x"05",
          6878 => x"33",
          6879 => x"05",
          6880 => x"40",
          6881 => x"da",
          6882 => x"cc",
          6883 => x"87",
          6884 => x"bd",
          6885 => x"33",
          6886 => x"b5",
          6887 => x"2e",
          6888 => x"1a",
          6889 => x"90",
          6890 => x"33",
          6891 => x"70",
          6892 => x"55",
          6893 => x"38",
          6894 => x"97",
          6895 => x"82",
          6896 => x"58",
          6897 => x"7e",
          6898 => x"70",
          6899 => x"55",
          6900 => x"56",
          6901 => x"93",
          6902 => x"7d",
          6903 => x"70",
          6904 => x"2a",
          6905 => x"08",
          6906 => x"08",
          6907 => x"5d",
          6908 => x"77",
          6909 => x"98",
          6910 => x"26",
          6911 => x"57",
          6912 => x"59",
          6913 => x"52",
          6914 => x"ae",
          6915 => x"15",
          6916 => x"98",
          6917 => x"26",
          6918 => x"55",
          6919 => x"08",
          6920 => x"99",
          6921 => x"cc",
          6922 => x"ff",
          6923 => x"87",
          6924 => x"38",
          6925 => x"75",
          6926 => x"81",
          6927 => x"93",
          6928 => x"80",
          6929 => x"2e",
          6930 => x"ff",
          6931 => x"58",
          6932 => x"7d",
          6933 => x"38",
          6934 => x"55",
          6935 => x"b4",
          6936 => x"56",
          6937 => x"09",
          6938 => x"38",
          6939 => x"53",
          6940 => x"51",
          6941 => x"3f",
          6942 => x"08",
          6943 => x"cc",
          6944 => x"38",
          6945 => x"ff",
          6946 => x"5c",
          6947 => x"84",
          6948 => x"5c",
          6949 => x"12",
          6950 => x"80",
          6951 => x"78",
          6952 => x"7c",
          6953 => x"90",
          6954 => x"c0",
          6955 => x"90",
          6956 => x"15",
          6957 => x"90",
          6958 => x"54",
          6959 => x"91",
          6960 => x"31",
          6961 => x"84",
          6962 => x"07",
          6963 => x"16",
          6964 => x"73",
          6965 => x"0c",
          6966 => x"04",
          6967 => x"6b",
          6968 => x"05",
          6969 => x"33",
          6970 => x"5a",
          6971 => x"be",
          6972 => x"80",
          6973 => x"cc",
          6974 => x"f8",
          6975 => x"cc",
          6976 => x"82",
          6977 => x"70",
          6978 => x"74",
          6979 => x"38",
          6980 => x"82",
          6981 => x"81",
          6982 => x"81",
          6983 => x"ff",
          6984 => x"82",
          6985 => x"81",
          6986 => x"81",
          6987 => x"83",
          6988 => x"c0",
          6989 => x"2a",
          6990 => x"51",
          6991 => x"74",
          6992 => x"99",
          6993 => x"53",
          6994 => x"51",
          6995 => x"3f",
          6996 => x"08",
          6997 => x"55",
          6998 => x"92",
          6999 => x"80",
          7000 => x"38",
          7001 => x"06",
          7002 => x"2e",
          7003 => x"48",
          7004 => x"87",
          7005 => x"79",
          7006 => x"78",
          7007 => x"26",
          7008 => x"19",
          7009 => x"74",
          7010 => x"38",
          7011 => x"e4",
          7012 => x"2a",
          7013 => x"70",
          7014 => x"59",
          7015 => x"7a",
          7016 => x"56",
          7017 => x"80",
          7018 => x"51",
          7019 => x"74",
          7020 => x"99",
          7021 => x"53",
          7022 => x"51",
          7023 => x"3f",
          7024 => x"87",
          7025 => x"ac",
          7026 => x"2a",
          7027 => x"82",
          7028 => x"43",
          7029 => x"83",
          7030 => x"66",
          7031 => x"60",
          7032 => x"90",
          7033 => x"31",
          7034 => x"80",
          7035 => x"8a",
          7036 => x"56",
          7037 => x"26",
          7038 => x"77",
          7039 => x"81",
          7040 => x"74",
          7041 => x"38",
          7042 => x"55",
          7043 => x"83",
          7044 => x"81",
          7045 => x"80",
          7046 => x"38",
          7047 => x"55",
          7048 => x"5e",
          7049 => x"89",
          7050 => x"5a",
          7051 => x"09",
          7052 => x"e1",
          7053 => x"38",
          7054 => x"57",
          7055 => x"82",
          7056 => x"5a",
          7057 => x"9d",
          7058 => x"26",
          7059 => x"82",
          7060 => x"10",
          7061 => x"22",
          7062 => x"74",
          7063 => x"38",
          7064 => x"ee",
          7065 => x"66",
          7066 => x"ff",
          7067 => x"cc",
          7068 => x"84",
          7069 => x"89",
          7070 => x"a0",
          7071 => x"82",
          7072 => x"fc",
          7073 => x"56",
          7074 => x"f0",
          7075 => x"80",
          7076 => x"d3",
          7077 => x"38",
          7078 => x"57",
          7079 => x"82",
          7080 => x"5a",
          7081 => x"9d",
          7082 => x"26",
          7083 => x"82",
          7084 => x"10",
          7085 => x"22",
          7086 => x"74",
          7087 => x"38",
          7088 => x"ee",
          7089 => x"66",
          7090 => x"9f",
          7091 => x"cc",
          7092 => x"05",
          7093 => x"cc",
          7094 => x"26",
          7095 => x"0b",
          7096 => x"08",
          7097 => x"cc",
          7098 => x"11",
          7099 => x"05",
          7100 => x"83",
          7101 => x"2a",
          7102 => x"a0",
          7103 => x"7d",
          7104 => x"69",
          7105 => x"05",
          7106 => x"72",
          7107 => x"5c",
          7108 => x"59",
          7109 => x"2e",
          7110 => x"89",
          7111 => x"60",
          7112 => x"84",
          7113 => x"5d",
          7114 => x"18",
          7115 => x"68",
          7116 => x"74",
          7117 => x"af",
          7118 => x"31",
          7119 => x"53",
          7120 => x"52",
          7121 => x"a3",
          7122 => x"cc",
          7123 => x"83",
          7124 => x"06",
          7125 => x"87",
          7126 => x"ff",
          7127 => x"dd",
          7128 => x"83",
          7129 => x"2a",
          7130 => x"be",
          7131 => x"39",
          7132 => x"09",
          7133 => x"c5",
          7134 => x"f5",
          7135 => x"cc",
          7136 => x"38",
          7137 => x"79",
          7138 => x"80",
          7139 => x"38",
          7140 => x"96",
          7141 => x"06",
          7142 => x"2e",
          7143 => x"5e",
          7144 => x"82",
          7145 => x"9f",
          7146 => x"38",
          7147 => x"38",
          7148 => x"81",
          7149 => x"fc",
          7150 => x"ab",
          7151 => x"7d",
          7152 => x"81",
          7153 => x"7d",
          7154 => x"78",
          7155 => x"74",
          7156 => x"8e",
          7157 => x"9c",
          7158 => x"53",
          7159 => x"51",
          7160 => x"3f",
          7161 => x"80",
          7162 => x"51",
          7163 => x"3f",
          7164 => x"8b",
          7165 => x"a1",
          7166 => x"8d",
          7167 => x"83",
          7168 => x"52",
          7169 => x"ff",
          7170 => x"81",
          7171 => x"34",
          7172 => x"70",
          7173 => x"2a",
          7174 => x"54",
          7175 => x"1b",
          7176 => x"89",
          7177 => x"74",
          7178 => x"26",
          7179 => x"83",
          7180 => x"52",
          7181 => x"ff",
          7182 => x"8a",
          7183 => x"a0",
          7184 => x"a1",
          7185 => x"0b",
          7186 => x"bf",
          7187 => x"51",
          7188 => x"3f",
          7189 => x"9a",
          7190 => x"a0",
          7191 => x"52",
          7192 => x"ff",
          7193 => x"7d",
          7194 => x"81",
          7195 => x"38",
          7196 => x"0a",
          7197 => x"1b",
          7198 => x"cf",
          7199 => x"a4",
          7200 => x"a0",
          7201 => x"52",
          7202 => x"ff",
          7203 => x"81",
          7204 => x"51",
          7205 => x"3f",
          7206 => x"1b",
          7207 => x"8d",
          7208 => x"0b",
          7209 => x"34",
          7210 => x"c2",
          7211 => x"53",
          7212 => x"52",
          7213 => x"51",
          7214 => x"88",
          7215 => x"a7",
          7216 => x"a0",
          7217 => x"83",
          7218 => x"52",
          7219 => x"ff",
          7220 => x"ff",
          7221 => x"1c",
          7222 => x"a6",
          7223 => x"53",
          7224 => x"52",
          7225 => x"ff",
          7226 => x"82",
          7227 => x"83",
          7228 => x"52",
          7229 => x"b5",
          7230 => x"60",
          7231 => x"7e",
          7232 => x"d8",
          7233 => x"82",
          7234 => x"83",
          7235 => x"83",
          7236 => x"06",
          7237 => x"75",
          7238 => x"05",
          7239 => x"7e",
          7240 => x"b8",
          7241 => x"53",
          7242 => x"51",
          7243 => x"3f",
          7244 => x"a4",
          7245 => x"51",
          7246 => x"3f",
          7247 => x"e4",
          7248 => x"e4",
          7249 => x"9f",
          7250 => x"18",
          7251 => x"1b",
          7252 => x"f7",
          7253 => x"83",
          7254 => x"ff",
          7255 => x"82",
          7256 => x"78",
          7257 => x"c5",
          7258 => x"60",
          7259 => x"7a",
          7260 => x"ff",
          7261 => x"75",
          7262 => x"53",
          7263 => x"51",
          7264 => x"3f",
          7265 => x"52",
          7266 => x"9f",
          7267 => x"56",
          7268 => x"83",
          7269 => x"06",
          7270 => x"52",
          7271 => x"9e",
          7272 => x"52",
          7273 => x"ff",
          7274 => x"f0",
          7275 => x"1b",
          7276 => x"87",
          7277 => x"55",
          7278 => x"83",
          7279 => x"74",
          7280 => x"ff",
          7281 => x"7c",
          7282 => x"74",
          7283 => x"38",
          7284 => x"54",
          7285 => x"52",
          7286 => x"99",
          7287 => x"87",
          7288 => x"87",
          7289 => x"53",
          7290 => x"08",
          7291 => x"ff",
          7292 => x"76",
          7293 => x"31",
          7294 => x"cd",
          7295 => x"58",
          7296 => x"ff",
          7297 => x"55",
          7298 => x"83",
          7299 => x"61",
          7300 => x"26",
          7301 => x"57",
          7302 => x"53",
          7303 => x"51",
          7304 => x"3f",
          7305 => x"08",
          7306 => x"76",
          7307 => x"31",
          7308 => x"db",
          7309 => x"7d",
          7310 => x"38",
          7311 => x"83",
          7312 => x"8a",
          7313 => x"7d",
          7314 => x"38",
          7315 => x"81",
          7316 => x"80",
          7317 => x"80",
          7318 => x"7a",
          7319 => x"bd",
          7320 => x"d5",
          7321 => x"ff",
          7322 => x"83",
          7323 => x"77",
          7324 => x"0b",
          7325 => x"81",
          7326 => x"34",
          7327 => x"34",
          7328 => x"34",
          7329 => x"56",
          7330 => x"52",
          7331 => x"86",
          7332 => x"0b",
          7333 => x"82",
          7334 => x"82",
          7335 => x"56",
          7336 => x"34",
          7337 => x"08",
          7338 => x"60",
          7339 => x"1b",
          7340 => x"97",
          7341 => x"83",
          7342 => x"ff",
          7343 => x"81",
          7344 => x"7a",
          7345 => x"ff",
          7346 => x"81",
          7347 => x"cc",
          7348 => x"80",
          7349 => x"7e",
          7350 => x"e4",
          7351 => x"82",
          7352 => x"90",
          7353 => x"8e",
          7354 => x"81",
          7355 => x"82",
          7356 => x"56",
          7357 => x"cc",
          7358 => x"0d",
          7359 => x"0d",
          7360 => x"59",
          7361 => x"ff",
          7362 => x"57",
          7363 => x"b4",
          7364 => x"f8",
          7365 => x"81",
          7366 => x"52",
          7367 => x"dc",
          7368 => x"2e",
          7369 => x"9c",
          7370 => x"33",
          7371 => x"2e",
          7372 => x"76",
          7373 => x"58",
          7374 => x"57",
          7375 => x"09",
          7376 => x"38",
          7377 => x"78",
          7378 => x"38",
          7379 => x"82",
          7380 => x"8d",
          7381 => x"f7",
          7382 => x"02",
          7383 => x"05",
          7384 => x"77",
          7385 => x"81",
          7386 => x"8d",
          7387 => x"e7",
          7388 => x"08",
          7389 => x"24",
          7390 => x"17",
          7391 => x"8c",
          7392 => x"77",
          7393 => x"16",
          7394 => x"25",
          7395 => x"3d",
          7396 => x"75",
          7397 => x"52",
          7398 => x"cb",
          7399 => x"76",
          7400 => x"70",
          7401 => x"2a",
          7402 => x"51",
          7403 => x"84",
          7404 => x"19",
          7405 => x"8b",
          7406 => x"f9",
          7407 => x"84",
          7408 => x"56",
          7409 => x"a7",
          7410 => x"fc",
          7411 => x"53",
          7412 => x"75",
          7413 => x"a1",
          7414 => x"cc",
          7415 => x"84",
          7416 => x"2e",
          7417 => x"87",
          7418 => x"08",
          7419 => x"ff",
          7420 => x"87",
          7421 => x"3d",
          7422 => x"3d",
          7423 => x"80",
          7424 => x"52",
          7425 => x"9a",
          7426 => x"74",
          7427 => x"0d",
          7428 => x"0d",
          7429 => x"05",
          7430 => x"86",
          7431 => x"54",
          7432 => x"73",
          7433 => x"fe",
          7434 => x"51",
          7435 => x"98",
          7436 => x"00",
          7437 => x"ff",
          7438 => x"ff",
          7439 => x"ff",
          7440 => x"00",
          7441 => x"06",
          7442 => x"8a",
          7443 => x"91",
          7444 => x"98",
          7445 => x"9f",
          7446 => x"a6",
          7447 => x"ad",
          7448 => x"b4",
          7449 => x"bb",
          7450 => x"c2",
          7451 => x"c9",
          7452 => x"d0",
          7453 => x"d6",
          7454 => x"dc",
          7455 => x"e2",
          7456 => x"e8",
          7457 => x"ee",
          7458 => x"f4",
          7459 => x"fa",
          7460 => x"00",
          7461 => x"42",
          7462 => x"48",
          7463 => x"4e",
          7464 => x"54",
          7465 => x"5a",
          7466 => x"7c",
          7467 => x"70",
          7468 => x"63",
          7469 => x"97",
          7470 => x"58",
          7471 => x"51",
          7472 => x"13",
          7473 => x"6e",
          7474 => x"50",
          7475 => x"e6",
          7476 => x"6c",
          7477 => x"13",
          7478 => x"51",
          7479 => x"63",
          7480 => x"86",
          7481 => x"13",
          7482 => x"51",
          7483 => x"51",
          7484 => x"6c",
          7485 => x"e6",
          7486 => x"6e",
          7487 => x"97",
          7488 => x"69",
          7489 => x"00",
          7490 => x"63",
          7491 => x"00",
          7492 => x"69",
          7493 => x"00",
          7494 => x"61",
          7495 => x"00",
          7496 => x"65",
          7497 => x"00",
          7498 => x"65",
          7499 => x"00",
          7500 => x"70",
          7501 => x"00",
          7502 => x"66",
          7503 => x"00",
          7504 => x"6d",
          7505 => x"00",
          7506 => x"00",
          7507 => x"00",
          7508 => x"00",
          7509 => x"00",
          7510 => x"00",
          7511 => x"00",
          7512 => x"00",
          7513 => x"6c",
          7514 => x"00",
          7515 => x"00",
          7516 => x"74",
          7517 => x"00",
          7518 => x"65",
          7519 => x"00",
          7520 => x"6f",
          7521 => x"00",
          7522 => x"74",
          7523 => x"00",
          7524 => x"73",
          7525 => x"00",
          7526 => x"73",
          7527 => x"00",
          7528 => x"6f",
          7529 => x"00",
          7530 => x"00",
          7531 => x"6b",
          7532 => x"72",
          7533 => x"00",
          7534 => x"65",
          7535 => x"6c",
          7536 => x"72",
          7537 => x"0a",
          7538 => x"00",
          7539 => x"6b",
          7540 => x"74",
          7541 => x"61",
          7542 => x"0a",
          7543 => x"00",
          7544 => x"66",
          7545 => x"20",
          7546 => x"6e",
          7547 => x"00",
          7548 => x"70",
          7549 => x"20",
          7550 => x"6e",
          7551 => x"00",
          7552 => x"61",
          7553 => x"20",
          7554 => x"65",
          7555 => x"65",
          7556 => x"00",
          7557 => x"65",
          7558 => x"64",
          7559 => x"65",
          7560 => x"00",
          7561 => x"65",
          7562 => x"72",
          7563 => x"79",
          7564 => x"69",
          7565 => x"2e",
          7566 => x"00",
          7567 => x"65",
          7568 => x"6e",
          7569 => x"20",
          7570 => x"61",
          7571 => x"2e",
          7572 => x"00",
          7573 => x"69",
          7574 => x"72",
          7575 => x"20",
          7576 => x"74",
          7577 => x"65",
          7578 => x"00",
          7579 => x"76",
          7580 => x"75",
          7581 => x"72",
          7582 => x"20",
          7583 => x"61",
          7584 => x"2e",
          7585 => x"00",
          7586 => x"6b",
          7587 => x"74",
          7588 => x"61",
          7589 => x"64",
          7590 => x"00",
          7591 => x"63",
          7592 => x"61",
          7593 => x"6c",
          7594 => x"69",
          7595 => x"79",
          7596 => x"6d",
          7597 => x"75",
          7598 => x"6f",
          7599 => x"69",
          7600 => x"0a",
          7601 => x"00",
          7602 => x"6d",
          7603 => x"61",
          7604 => x"74",
          7605 => x"0a",
          7606 => x"00",
          7607 => x"65",
          7608 => x"2c",
          7609 => x"65",
          7610 => x"69",
          7611 => x"63",
          7612 => x"65",
          7613 => x"64",
          7614 => x"00",
          7615 => x"65",
          7616 => x"20",
          7617 => x"6b",
          7618 => x"0a",
          7619 => x"00",
          7620 => x"75",
          7621 => x"63",
          7622 => x"74",
          7623 => x"6d",
          7624 => x"2e",
          7625 => x"00",
          7626 => x"20",
          7627 => x"79",
          7628 => x"65",
          7629 => x"69",
          7630 => x"2e",
          7631 => x"00",
          7632 => x"61",
          7633 => x"65",
          7634 => x"69",
          7635 => x"72",
          7636 => x"74",
          7637 => x"00",
          7638 => x"63",
          7639 => x"2e",
          7640 => x"00",
          7641 => x"6e",
          7642 => x"20",
          7643 => x"6f",
          7644 => x"00",
          7645 => x"75",
          7646 => x"74",
          7647 => x"25",
          7648 => x"74",
          7649 => x"75",
          7650 => x"74",
          7651 => x"73",
          7652 => x"0a",
          7653 => x"00",
          7654 => x"64",
          7655 => x"00",
          7656 => x"58",
          7657 => x"00",
          7658 => x"00",
          7659 => x"58",
          7660 => x"00",
          7661 => x"20",
          7662 => x"20",
          7663 => x"00",
          7664 => x"58",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"54",
          7670 => x"00",
          7671 => x"20",
          7672 => x"28",
          7673 => x"00",
          7674 => x"30",
          7675 => x"30",
          7676 => x"00",
          7677 => x"35",
          7678 => x"00",
          7679 => x"55",
          7680 => x"65",
          7681 => x"30",
          7682 => x"20",
          7683 => x"25",
          7684 => x"2a",
          7685 => x"00",
          7686 => x"54",
          7687 => x"6e",
          7688 => x"72",
          7689 => x"20",
          7690 => x"64",
          7691 => x"0a",
          7692 => x"00",
          7693 => x"65",
          7694 => x"6e",
          7695 => x"72",
          7696 => x"0a",
          7697 => x"00",
          7698 => x"20",
          7699 => x"65",
          7700 => x"70",
          7701 => x"00",
          7702 => x"54",
          7703 => x"44",
          7704 => x"74",
          7705 => x"75",
          7706 => x"00",
          7707 => x"54",
          7708 => x"52",
          7709 => x"74",
          7710 => x"75",
          7711 => x"00",
          7712 => x"54",
          7713 => x"58",
          7714 => x"74",
          7715 => x"75",
          7716 => x"00",
          7717 => x"54",
          7718 => x"58",
          7719 => x"74",
          7720 => x"75",
          7721 => x"00",
          7722 => x"54",
          7723 => x"58",
          7724 => x"74",
          7725 => x"75",
          7726 => x"00",
          7727 => x"54",
          7728 => x"58",
          7729 => x"74",
          7730 => x"75",
          7731 => x"00",
          7732 => x"74",
          7733 => x"20",
          7734 => x"74",
          7735 => x"72",
          7736 => x"0a",
          7737 => x"00",
          7738 => x"62",
          7739 => x"67",
          7740 => x"6d",
          7741 => x"2e",
          7742 => x"00",
          7743 => x"6f",
          7744 => x"63",
          7745 => x"74",
          7746 => x"00",
          7747 => x"74",
          7748 => x"73",
          7749 => x"00",
          7750 => x"00",
          7751 => x"6c",
          7752 => x"74",
          7753 => x"6e",
          7754 => x"61",
          7755 => x"65",
          7756 => x"20",
          7757 => x"64",
          7758 => x"20",
          7759 => x"61",
          7760 => x"69",
          7761 => x"20",
          7762 => x"75",
          7763 => x"79",
          7764 => x"00",
          7765 => x"00",
          7766 => x"20",
          7767 => x"6b",
          7768 => x"21",
          7769 => x"00",
          7770 => x"74",
          7771 => x"69",
          7772 => x"2e",
          7773 => x"00",
          7774 => x"6c",
          7775 => x"74",
          7776 => x"6e",
          7777 => x"61",
          7778 => x"65",
          7779 => x"00",
          7780 => x"25",
          7781 => x"00",
          7782 => x"00",
          7783 => x"61",
          7784 => x"67",
          7785 => x"2e",
          7786 => x"00",
          7787 => x"79",
          7788 => x"2e",
          7789 => x"00",
          7790 => x"70",
          7791 => x"6e",
          7792 => x"2e",
          7793 => x"00",
          7794 => x"6c",
          7795 => x"30",
          7796 => x"2d",
          7797 => x"38",
          7798 => x"25",
          7799 => x"29",
          7800 => x"00",
          7801 => x"70",
          7802 => x"6d",
          7803 => x"0a",
          7804 => x"00",
          7805 => x"6d",
          7806 => x"74",
          7807 => x"00",
          7808 => x"58",
          7809 => x"32",
          7810 => x"00",
          7811 => x"0a",
          7812 => x"00",
          7813 => x"58",
          7814 => x"34",
          7815 => x"00",
          7816 => x"58",
          7817 => x"38",
          7818 => x"00",
          7819 => x"61",
          7820 => x"6e",
          7821 => x"6e",
          7822 => x"72",
          7823 => x"73",
          7824 => x"00",
          7825 => x"62",
          7826 => x"67",
          7827 => x"74",
          7828 => x"75",
          7829 => x"0a",
          7830 => x"00",
          7831 => x"61",
          7832 => x"64",
          7833 => x"72",
          7834 => x"69",
          7835 => x"00",
          7836 => x"62",
          7837 => x"67",
          7838 => x"72",
          7839 => x"69",
          7840 => x"00",
          7841 => x"63",
          7842 => x"6e",
          7843 => x"6f",
          7844 => x"40",
          7845 => x"38",
          7846 => x"2e",
          7847 => x"00",
          7848 => x"6c",
          7849 => x"20",
          7850 => x"65",
          7851 => x"25",
          7852 => x"20",
          7853 => x"0a",
          7854 => x"00",
          7855 => x"6c",
          7856 => x"74",
          7857 => x"65",
          7858 => x"6f",
          7859 => x"28",
          7860 => x"2e",
          7861 => x"00",
          7862 => x"74",
          7863 => x"69",
          7864 => x"61",
          7865 => x"69",
          7866 => x"69",
          7867 => x"2e",
          7868 => x"00",
          7869 => x"64",
          7870 => x"62",
          7871 => x"69",
          7872 => x"2e",
          7873 => x"00",
          7874 => x"00",
          7875 => x"00",
          7876 => x"5c",
          7877 => x"25",
          7878 => x"73",
          7879 => x"00",
          7880 => x"5c",
          7881 => x"25",
          7882 => x"00",
          7883 => x"5c",
          7884 => x"00",
          7885 => x"20",
          7886 => x"6d",
          7887 => x"2e",
          7888 => x"00",
          7889 => x"6e",
          7890 => x"2e",
          7891 => x"00",
          7892 => x"62",
          7893 => x"67",
          7894 => x"74",
          7895 => x"75",
          7896 => x"2e",
          7897 => x"00",
          7898 => x"25",
          7899 => x"64",
          7900 => x"3a",
          7901 => x"25",
          7902 => x"64",
          7903 => x"00",
          7904 => x"20",
          7905 => x"66",
          7906 => x"72",
          7907 => x"6f",
          7908 => x"00",
          7909 => x"72",
          7910 => x"53",
          7911 => x"63",
          7912 => x"69",
          7913 => x"00",
          7914 => x"65",
          7915 => x"65",
          7916 => x"6d",
          7917 => x"6d",
          7918 => x"65",
          7919 => x"00",
          7920 => x"20",
          7921 => x"53",
          7922 => x"4d",
          7923 => x"25",
          7924 => x"3a",
          7925 => x"58",
          7926 => x"00",
          7927 => x"20",
          7928 => x"41",
          7929 => x"20",
          7930 => x"25",
          7931 => x"3a",
          7932 => x"58",
          7933 => x"00",
          7934 => x"20",
          7935 => x"4e",
          7936 => x"41",
          7937 => x"25",
          7938 => x"3a",
          7939 => x"58",
          7940 => x"00",
          7941 => x"20",
          7942 => x"4d",
          7943 => x"20",
          7944 => x"25",
          7945 => x"3a",
          7946 => x"58",
          7947 => x"00",
          7948 => x"20",
          7949 => x"20",
          7950 => x"20",
          7951 => x"25",
          7952 => x"3a",
          7953 => x"58",
          7954 => x"00",
          7955 => x"20",
          7956 => x"43",
          7957 => x"20",
          7958 => x"44",
          7959 => x"63",
          7960 => x"3d",
          7961 => x"64",
          7962 => x"00",
          7963 => x"20",
          7964 => x"45",
          7965 => x"20",
          7966 => x"54",
          7967 => x"72",
          7968 => x"3d",
          7969 => x"64",
          7970 => x"00",
          7971 => x"20",
          7972 => x"52",
          7973 => x"52",
          7974 => x"43",
          7975 => x"6e",
          7976 => x"3d",
          7977 => x"64",
          7978 => x"00",
          7979 => x"20",
          7980 => x"48",
          7981 => x"45",
          7982 => x"53",
          7983 => x"00",
          7984 => x"20",
          7985 => x"49",
          7986 => x"00",
          7987 => x"20",
          7988 => x"54",
          7989 => x"00",
          7990 => x"20",
          7991 => x"0a",
          7992 => x"00",
          7993 => x"20",
          7994 => x"0a",
          7995 => x"00",
          7996 => x"72",
          7997 => x"65",
          7998 => x"00",
          7999 => x"20",
          8000 => x"20",
          8001 => x"65",
          8002 => x"65",
          8003 => x"72",
          8004 => x"64",
          8005 => x"73",
          8006 => x"25",
          8007 => x"0a",
          8008 => x"00",
          8009 => x"20",
          8010 => x"20",
          8011 => x"6f",
          8012 => x"53",
          8013 => x"74",
          8014 => x"64",
          8015 => x"73",
          8016 => x"25",
          8017 => x"0a",
          8018 => x"00",
          8019 => x"20",
          8020 => x"63",
          8021 => x"74",
          8022 => x"20",
          8023 => x"72",
          8024 => x"20",
          8025 => x"20",
          8026 => x"25",
          8027 => x"0a",
          8028 => x"00",
          8029 => x"63",
          8030 => x"00",
          8031 => x"20",
          8032 => x"20",
          8033 => x"20",
          8034 => x"20",
          8035 => x"20",
          8036 => x"20",
          8037 => x"20",
          8038 => x"25",
          8039 => x"0a",
          8040 => x"00",
          8041 => x"20",
          8042 => x"74",
          8043 => x"43",
          8044 => x"6b",
          8045 => x"65",
          8046 => x"20",
          8047 => x"20",
          8048 => x"25",
          8049 => x"30",
          8050 => x"48",
          8051 => x"00",
          8052 => x"20",
          8053 => x"41",
          8054 => x"6c",
          8055 => x"20",
          8056 => x"71",
          8057 => x"20",
          8058 => x"20",
          8059 => x"25",
          8060 => x"30",
          8061 => x"48",
          8062 => x"00",
          8063 => x"20",
          8064 => x"68",
          8065 => x"65",
          8066 => x"52",
          8067 => x"43",
          8068 => x"6b",
          8069 => x"65",
          8070 => x"25",
          8071 => x"30",
          8072 => x"48",
          8073 => x"00",
          8074 => x"6c",
          8075 => x"00",
          8076 => x"69",
          8077 => x"00",
          8078 => x"78",
          8079 => x"00",
          8080 => x"00",
          8081 => x"6d",
          8082 => x"00",
          8083 => x"6e",
          8084 => x"00",
          8085 => x"b0",
          8086 => x"00",
          8087 => x"02",
          8088 => x"ac",
          8089 => x"00",
          8090 => x"03",
          8091 => x"a8",
          8092 => x"00",
          8093 => x"04",
          8094 => x"a4",
          8095 => x"00",
          8096 => x"05",
          8097 => x"a0",
          8098 => x"00",
          8099 => x"06",
          8100 => x"9c",
          8101 => x"00",
          8102 => x"07",
          8103 => x"98",
          8104 => x"00",
          8105 => x"01",
          8106 => x"94",
          8107 => x"00",
          8108 => x"08",
          8109 => x"90",
          8110 => x"00",
          8111 => x"0b",
          8112 => x"8c",
          8113 => x"00",
          8114 => x"09",
          8115 => x"88",
          8116 => x"00",
          8117 => x"0a",
          8118 => x"84",
          8119 => x"00",
          8120 => x"0d",
          8121 => x"80",
          8122 => x"00",
          8123 => x"0c",
          8124 => x"7c",
          8125 => x"00",
          8126 => x"0e",
          8127 => x"78",
          8128 => x"00",
          8129 => x"0f",
          8130 => x"74",
          8131 => x"00",
          8132 => x"0f",
          8133 => x"70",
          8134 => x"00",
          8135 => x"10",
          8136 => x"6c",
          8137 => x"00",
          8138 => x"11",
          8139 => x"68",
          8140 => x"00",
          8141 => x"12",
          8142 => x"64",
          8143 => x"00",
          8144 => x"13",
          8145 => x"60",
          8146 => x"00",
          8147 => x"14",
          8148 => x"5c",
          8149 => x"00",
          8150 => x"15",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"7e",
          8156 => x"7e",
          8157 => x"7e",
          8158 => x"00",
          8159 => x"7e",
          8160 => x"7e",
          8161 => x"7e",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"74",
          8174 => x"00",
          8175 => x"74",
          8176 => x"00",
          8177 => x"00",
          8178 => x"64",
          8179 => x"73",
          8180 => x"00",
          8181 => x"6c",
          8182 => x"74",
          8183 => x"65",
          8184 => x"20",
          8185 => x"20",
          8186 => x"74",
          8187 => x"20",
          8188 => x"65",
          8189 => x"20",
          8190 => x"2e",
          8191 => x"00",
          8192 => x"6e",
          8193 => x"6f",
          8194 => x"2f",
          8195 => x"61",
          8196 => x"68",
          8197 => x"6f",
          8198 => x"66",
          8199 => x"2c",
          8200 => x"73",
          8201 => x"69",
          8202 => x"0a",
          8203 => x"00",
          8204 => x"00",
          8205 => x"2c",
          8206 => x"3d",
          8207 => x"5d",
          8208 => x"00",
          8209 => x"00",
          8210 => x"33",
          8211 => x"00",
          8212 => x"4d",
          8213 => x"53",
          8214 => x"00",
          8215 => x"4e",
          8216 => x"20",
          8217 => x"46",
          8218 => x"32",
          8219 => x"00",
          8220 => x"4e",
          8221 => x"20",
          8222 => x"46",
          8223 => x"20",
          8224 => x"00",
          8225 => x"30",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"41",
          8230 => x"80",
          8231 => x"49",
          8232 => x"8f",
          8233 => x"4f",
          8234 => x"55",
          8235 => x"9b",
          8236 => x"9f",
          8237 => x"55",
          8238 => x"a7",
          8239 => x"ab",
          8240 => x"af",
          8241 => x"b3",
          8242 => x"b7",
          8243 => x"bb",
          8244 => x"bf",
          8245 => x"c3",
          8246 => x"c7",
          8247 => x"cb",
          8248 => x"cf",
          8249 => x"d3",
          8250 => x"d7",
          8251 => x"db",
          8252 => x"df",
          8253 => x"e3",
          8254 => x"e7",
          8255 => x"eb",
          8256 => x"ef",
          8257 => x"f3",
          8258 => x"f7",
          8259 => x"fb",
          8260 => x"ff",
          8261 => x"3b",
          8262 => x"2f",
          8263 => x"3a",
          8264 => x"7c",
          8265 => x"00",
          8266 => x"04",
          8267 => x"40",
          8268 => x"00",
          8269 => x"00",
          8270 => x"02",
          8271 => x"08",
          8272 => x"20",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"08",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"10",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"18",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"20",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"28",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"30",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"38",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"40",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"48",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"4c",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"50",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"54",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"58",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"5c",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"60",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"64",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"6c",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"70",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"78",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"80",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"88",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"90",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"98",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"a0",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"a8",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"ff",
          8382 => x"00",
          8383 => x"ff",
          8384 => x"00",
          8385 => x"ff",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"ff",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"01",
          8399 => x"01",
          8400 => x"01",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"b4",
          8427 => x"00",
          8428 => x"bc",
          8429 => x"00",
          8430 => x"c4",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c4",
           273 => x"0b",
           274 => x"0b",
           275 => x"e4",
           276 => x"0b",
           277 => x"0b",
           278 => x"84",
           279 => x"0b",
           280 => x"0b",
           281 => x"a4",
           282 => x"0b",
           283 => x"0b",
           284 => x"c4",
           285 => x"0b",
           286 => x"0b",
           287 => x"e4",
           288 => x"0b",
           289 => x"0b",
           290 => x"83",
           291 => x"0b",
           292 => x"0b",
           293 => x"a1",
           294 => x"0b",
           295 => x"0b",
           296 => x"c1",
           297 => x"0b",
           298 => x"0b",
           299 => x"e1",
           300 => x"0b",
           301 => x"0b",
           302 => x"81",
           303 => x"0b",
           304 => x"0b",
           305 => x"a1",
           306 => x"0b",
           307 => x"0b",
           308 => x"c1",
           309 => x"0b",
           310 => x"0b",
           311 => x"e1",
           312 => x"0b",
           313 => x"0b",
           314 => x"81",
           315 => x"0b",
           316 => x"0b",
           317 => x"a1",
           318 => x"0b",
           319 => x"0b",
           320 => x"c1",
           321 => x"0b",
           322 => x"0b",
           323 => x"e1",
           324 => x"0b",
           325 => x"0b",
           326 => x"81",
           327 => x"0b",
           328 => x"0b",
           329 => x"a1",
           330 => x"0b",
           331 => x"0b",
           332 => x"c1",
           333 => x"0b",
           334 => x"0b",
           335 => x"e1",
           336 => x"0b",
           337 => x"0b",
           338 => x"81",
           339 => x"0b",
           340 => x"0b",
           341 => x"9f",
           342 => x"0b",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"87",
           386 => x"97",
           387 => x"d8",
           388 => x"90",
           389 => x"d8",
           390 => x"c3",
           391 => x"d8",
           392 => x"90",
           393 => x"d8",
           394 => x"82",
           395 => x"d8",
           396 => x"90",
           397 => x"d8",
           398 => x"a0",
           399 => x"d8",
           400 => x"90",
           401 => x"d8",
           402 => x"de",
           403 => x"d8",
           404 => x"90",
           405 => x"d8",
           406 => x"dc",
           407 => x"d8",
           408 => x"90",
           409 => x"d8",
           410 => x"c3",
           411 => x"d8",
           412 => x"90",
           413 => x"d8",
           414 => x"f9",
           415 => x"d8",
           416 => x"90",
           417 => x"d8",
           418 => x"eb",
           419 => x"d8",
           420 => x"90",
           421 => x"d8",
           422 => x"84",
           423 => x"d8",
           424 => x"90",
           425 => x"d8",
           426 => x"f5",
           427 => x"d8",
           428 => x"90",
           429 => x"d8",
           430 => x"9a",
           431 => x"d8",
           432 => x"90",
           433 => x"d8",
           434 => x"be",
           435 => x"d8",
           436 => x"90",
           437 => x"d8",
           438 => x"a0",
           439 => x"d8",
           440 => x"90",
           441 => x"d8",
           442 => x"ef",
           443 => x"d8",
           444 => x"90",
           445 => x"d8",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"82",
           451 => x"82",
           452 => x"82",
           453 => x"bb",
           454 => x"87",
           455 => x"a0",
           456 => x"87",
           457 => x"ab",
           458 => x"87",
           459 => x"a0",
           460 => x"87",
           461 => x"b8",
           462 => x"87",
           463 => x"a0",
           464 => x"87",
           465 => x"af",
           466 => x"87",
           467 => x"a0",
           468 => x"87",
           469 => x"b2",
           470 => x"87",
           471 => x"a0",
           472 => x"87",
           473 => x"bd",
           474 => x"87",
           475 => x"a0",
           476 => x"87",
           477 => x"c5",
           478 => x"87",
           479 => x"a0",
           480 => x"87",
           481 => x"b6",
           482 => x"87",
           483 => x"a0",
           484 => x"87",
           485 => x"c0",
           486 => x"87",
           487 => x"a0",
           488 => x"87",
           489 => x"c1",
           490 => x"87",
           491 => x"a0",
           492 => x"87",
           493 => x"c1",
           494 => x"87",
           495 => x"a0",
           496 => x"87",
           497 => x"c9",
           498 => x"87",
           499 => x"a0",
           500 => x"87",
           501 => x"c7",
           502 => x"87",
           503 => x"a0",
           504 => x"87",
           505 => x"cc",
           506 => x"87",
           507 => x"a0",
           508 => x"87",
           509 => x"c2",
           510 => x"87",
           511 => x"a0",
           512 => x"87",
           513 => x"cf",
           514 => x"87",
           515 => x"a0",
           516 => x"87",
           517 => x"d0",
           518 => x"87",
           519 => x"a0",
           520 => x"87",
           521 => x"b8",
           522 => x"87",
           523 => x"a0",
           524 => x"87",
           525 => x"b8",
           526 => x"87",
           527 => x"a0",
           528 => x"87",
           529 => x"b9",
           530 => x"87",
           531 => x"a0",
           532 => x"87",
           533 => x"c3",
           534 => x"87",
           535 => x"a0",
           536 => x"87",
           537 => x"d1",
           538 => x"87",
           539 => x"a0",
           540 => x"87",
           541 => x"d3",
           542 => x"87",
           543 => x"a0",
           544 => x"87",
           545 => x"d6",
           546 => x"87",
           547 => x"a0",
           548 => x"87",
           549 => x"aa",
           550 => x"87",
           551 => x"a0",
           552 => x"87",
           553 => x"d9",
           554 => x"87",
           555 => x"a0",
           556 => x"87",
           557 => x"e8",
           558 => x"87",
           559 => x"a0",
           560 => x"87",
           561 => x"e5",
           562 => x"87",
           563 => x"a0",
           564 => x"87",
           565 => x"fb",
           566 => x"87",
           567 => x"a0",
           568 => x"87",
           569 => x"fd",
           570 => x"87",
           571 => x"a0",
           572 => x"87",
           573 => x"ff",
           574 => x"87",
           575 => x"a0",
           576 => x"87",
           577 => x"fc",
           578 => x"d8",
           579 => x"90",
           580 => x"d8",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"82",
           586 => x"82",
           587 => x"82",
           588 => x"9a",
           589 => x"87",
           590 => x"a0",
           591 => x"04",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"04",
           601 => x"81",
           602 => x"83",
           603 => x"05",
           604 => x"10",
           605 => x"72",
           606 => x"51",
           607 => x"72",
           608 => x"06",
           609 => x"72",
           610 => x"10",
           611 => x"10",
           612 => x"ed",
           613 => x"53",
           614 => x"87",
           615 => x"9f",
           616 => x"38",
           617 => x"84",
           618 => x"0b",
           619 => x"9c",
           620 => x"51",
           621 => x"00",
           622 => x"08",
           623 => x"d8",
           624 => x"0d",
           625 => x"08",
           626 => x"82",
           627 => x"fc",
           628 => x"87",
           629 => x"05",
           630 => x"33",
           631 => x"08",
           632 => x"81",
           633 => x"d8",
           634 => x"0c",
           635 => x"06",
           636 => x"80",
           637 => x"da",
           638 => x"d8",
           639 => x"08",
           640 => x"87",
           641 => x"05",
           642 => x"d8",
           643 => x"08",
           644 => x"08",
           645 => x"31",
           646 => x"cc",
           647 => x"3d",
           648 => x"d8",
           649 => x"87",
           650 => x"82",
           651 => x"fe",
           652 => x"87",
           653 => x"05",
           654 => x"d8",
           655 => x"0c",
           656 => x"08",
           657 => x"52",
           658 => x"87",
           659 => x"05",
           660 => x"82",
           661 => x"8c",
           662 => x"87",
           663 => x"05",
           664 => x"70",
           665 => x"87",
           666 => x"05",
           667 => x"82",
           668 => x"fc",
           669 => x"81",
           670 => x"70",
           671 => x"38",
           672 => x"82",
           673 => x"88",
           674 => x"82",
           675 => x"51",
           676 => x"82",
           677 => x"04",
           678 => x"08",
           679 => x"d8",
           680 => x"0d",
           681 => x"08",
           682 => x"82",
           683 => x"fc",
           684 => x"87",
           685 => x"05",
           686 => x"d8",
           687 => x"0c",
           688 => x"08",
           689 => x"80",
           690 => x"38",
           691 => x"08",
           692 => x"81",
           693 => x"d8",
           694 => x"0c",
           695 => x"08",
           696 => x"ff",
           697 => x"d8",
           698 => x"0c",
           699 => x"08",
           700 => x"80",
           701 => x"82",
           702 => x"f8",
           703 => x"70",
           704 => x"d8",
           705 => x"08",
           706 => x"87",
           707 => x"05",
           708 => x"d8",
           709 => x"08",
           710 => x"71",
           711 => x"d8",
           712 => x"08",
           713 => x"87",
           714 => x"05",
           715 => x"39",
           716 => x"08",
           717 => x"70",
           718 => x"0c",
           719 => x"0d",
           720 => x"0c",
           721 => x"d8",
           722 => x"87",
           723 => x"3d",
           724 => x"d8",
           725 => x"08",
           726 => x"f4",
           727 => x"d8",
           728 => x"08",
           729 => x"82",
           730 => x"8c",
           731 => x"05",
           732 => x"08",
           733 => x"82",
           734 => x"88",
           735 => x"33",
           736 => x"06",
           737 => x"51",
           738 => x"84",
           739 => x"39",
           740 => x"08",
           741 => x"52",
           742 => x"87",
           743 => x"05",
           744 => x"82",
           745 => x"88",
           746 => x"81",
           747 => x"51",
           748 => x"80",
           749 => x"d8",
           750 => x"0c",
           751 => x"82",
           752 => x"90",
           753 => x"05",
           754 => x"08",
           755 => x"82",
           756 => x"90",
           757 => x"2e",
           758 => x"81",
           759 => x"d8",
           760 => x"08",
           761 => x"e8",
           762 => x"d8",
           763 => x"08",
           764 => x"53",
           765 => x"ff",
           766 => x"d8",
           767 => x"0c",
           768 => x"82",
           769 => x"8c",
           770 => x"05",
           771 => x"08",
           772 => x"82",
           773 => x"8c",
           774 => x"33",
           775 => x"8c",
           776 => x"82",
           777 => x"fc",
           778 => x"39",
           779 => x"08",
           780 => x"70",
           781 => x"d8",
           782 => x"08",
           783 => x"71",
           784 => x"87",
           785 => x"05",
           786 => x"52",
           787 => x"39",
           788 => x"87",
           789 => x"05",
           790 => x"d8",
           791 => x"08",
           792 => x"0c",
           793 => x"82",
           794 => x"04",
           795 => x"08",
           796 => x"d8",
           797 => x"0d",
           798 => x"08",
           799 => x"82",
           800 => x"fc",
           801 => x"87",
           802 => x"05",
           803 => x"80",
           804 => x"87",
           805 => x"05",
           806 => x"82",
           807 => x"90",
           808 => x"87",
           809 => x"05",
           810 => x"82",
           811 => x"90",
           812 => x"87",
           813 => x"05",
           814 => x"a9",
           815 => x"d8",
           816 => x"08",
           817 => x"87",
           818 => x"05",
           819 => x"71",
           820 => x"87",
           821 => x"05",
           822 => x"82",
           823 => x"fc",
           824 => x"be",
           825 => x"d8",
           826 => x"08",
           827 => x"cc",
           828 => x"3d",
           829 => x"d8",
           830 => x"3d",
           831 => x"08",
           832 => x"58",
           833 => x"80",
           834 => x"39",
           835 => x"f9",
           836 => x"87",
           837 => x"78",
           838 => x"33",
           839 => x"39",
           840 => x"73",
           841 => x"81",
           842 => x"81",
           843 => x"39",
           844 => x"90",
           845 => x"cc",
           846 => x"52",
           847 => x"3f",
           848 => x"08",
           849 => x"75",
           850 => x"f9",
           851 => x"cc",
           852 => x"84",
           853 => x"73",
           854 => x"b0",
           855 => x"70",
           856 => x"58",
           857 => x"27",
           858 => x"54",
           859 => x"cc",
           860 => x"0d",
           861 => x"0d",
           862 => x"93",
           863 => x"38",
           864 => x"81",
           865 => x"52",
           866 => x"81",
           867 => x"81",
           868 => x"eb",
           869 => x"f9",
           870 => x"cc",
           871 => x"39",
           872 => x"51",
           873 => x"81",
           874 => x"80",
           875 => x"ec",
           876 => x"dd",
           877 => x"94",
           878 => x"39",
           879 => x"51",
           880 => x"81",
           881 => x"80",
           882 => x"ec",
           883 => x"c1",
           884 => x"ec",
           885 => x"81",
           886 => x"b5",
           887 => x"9c",
           888 => x"81",
           889 => x"a9",
           890 => x"dc",
           891 => x"81",
           892 => x"9d",
           893 => x"90",
           894 => x"81",
           895 => x"91",
           896 => x"c0",
           897 => x"81",
           898 => x"85",
           899 => x"e4",
           900 => x"3f",
           901 => x"04",
           902 => x"77",
           903 => x"74",
           904 => x"8a",
           905 => x"75",
           906 => x"51",
           907 => x"e8",
           908 => x"80",
           909 => x"82",
           910 => x"52",
           911 => x"cf",
           912 => x"87",
           913 => x"79",
           914 => x"81",
           915 => x"b5",
           916 => x"3d",
           917 => x"3d",
           918 => x"84",
           919 => x"05",
           920 => x"80",
           921 => x"70",
           922 => x"25",
           923 => x"59",
           924 => x"87",
           925 => x"38",
           926 => x"76",
           927 => x"ff",
           928 => x"93",
           929 => x"82",
           930 => x"76",
           931 => x"70",
           932 => x"8e",
           933 => x"87",
           934 => x"82",
           935 => x"b9",
           936 => x"cc",
           937 => x"98",
           938 => x"87",
           939 => x"96",
           940 => x"54",
           941 => x"77",
           942 => x"81",
           943 => x"82",
           944 => x"57",
           945 => x"08",
           946 => x"55",
           947 => x"89",
           948 => x"75",
           949 => x"d7",
           950 => x"d8",
           951 => x"9a",
           952 => x"30",
           953 => x"80",
           954 => x"70",
           955 => x"06",
           956 => x"56",
           957 => x"90",
           958 => x"98",
           959 => x"98",
           960 => x"78",
           961 => x"3f",
           962 => x"82",
           963 => x"96",
           964 => x"f9",
           965 => x"02",
           966 => x"05",
           967 => x"ff",
           968 => x"7a",
           969 => x"fe",
           970 => x"87",
           971 => x"38",
           972 => x"88",
           973 => x"2e",
           974 => x"39",
           975 => x"54",
           976 => x"53",
           977 => x"51",
           978 => x"87",
           979 => x"83",
           980 => x"76",
           981 => x"0c",
           982 => x"04",
           983 => x"7f",
           984 => x"8c",
           985 => x"05",
           986 => x"15",
           987 => x"5c",
           988 => x"5e",
           989 => x"ef",
           990 => x"89",
           991 => x"a8",
           992 => x"3f",
           993 => x"79",
           994 => x"38",
           995 => x"89",
           996 => x"2e",
           997 => x"c1",
           998 => x"53",
           999 => x"8d",
          1000 => x"52",
          1001 => x"51",
          1002 => x"88",
          1003 => x"b8",
          1004 => x"3f",
          1005 => x"bf",
          1006 => x"53",
          1007 => x"8d",
          1008 => x"52",
          1009 => x"51",
          1010 => x"88",
          1011 => x"b4",
          1012 => x"3f",
          1013 => x"9f",
          1014 => x"53",
          1015 => x"8d",
          1016 => x"52",
          1017 => x"51",
          1018 => x"88",
          1019 => x"c8",
          1020 => x"3f",
          1021 => x"a0",
          1022 => x"3f",
          1023 => x"81",
          1024 => x"ac",
          1025 => x"55",
          1026 => x"bb",
          1027 => x"70",
          1028 => x"80",
          1029 => x"27",
          1030 => x"56",
          1031 => x"74",
          1032 => x"81",
          1033 => x"06",
          1034 => x"06",
          1035 => x"80",
          1036 => x"73",
          1037 => x"85",
          1038 => x"83",
          1039 => x"ab",
          1040 => x"15",
          1041 => x"81",
          1042 => x"ab",
          1043 => x"18",
          1044 => x"58",
          1045 => x"82",
          1046 => x"98",
          1047 => x"2c",
          1048 => x"a0",
          1049 => x"06",
          1050 => x"84",
          1051 => x"cc",
          1052 => x"70",
          1053 => x"a0",
          1054 => x"72",
          1055 => x"30",
          1056 => x"73",
          1057 => x"51",
          1058 => x"57",
          1059 => x"73",
          1060 => x"76",
          1061 => x"81",
          1062 => x"80",
          1063 => x"7c",
          1064 => x"78",
          1065 => x"38",
          1066 => x"82",
          1067 => x"8f",
          1068 => x"fc",
          1069 => x"9b",
          1070 => x"ef",
          1071 => x"ef",
          1072 => x"b0",
          1073 => x"86",
          1074 => x"a8",
          1075 => x"ef",
          1076 => x"ef",
          1077 => x"86",
          1078 => x"81",
          1079 => x"b0",
          1080 => x"80",
          1081 => x"a4",
          1082 => x"3d",
          1083 => x"3d",
          1084 => x"96",
          1085 => x"a9",
          1086 => x"51",
          1087 => x"81",
          1088 => x"9d",
          1089 => x"51",
          1090 => x"72",
          1091 => x"81",
          1092 => x"71",
          1093 => x"38",
          1094 => x"f2",
          1095 => x"b4",
          1096 => x"3f",
          1097 => x"e6",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"51",
          1102 => x"81",
          1103 => x"9c",
          1104 => x"51",
          1105 => x"72",
          1106 => x"81",
          1107 => x"71",
          1108 => x"38",
          1109 => x"b6",
          1110 => x"d8",
          1111 => x"3f",
          1112 => x"aa",
          1113 => x"2a",
          1114 => x"51",
          1115 => x"2e",
          1116 => x"51",
          1117 => x"81",
          1118 => x"9c",
          1119 => x"51",
          1120 => x"72",
          1121 => x"81",
          1122 => x"71",
          1123 => x"38",
          1124 => x"fa",
          1125 => x"80",
          1126 => x"3f",
          1127 => x"ee",
          1128 => x"2a",
          1129 => x"51",
          1130 => x"2e",
          1131 => x"51",
          1132 => x"81",
          1133 => x"9b",
          1134 => x"51",
          1135 => x"72",
          1136 => x"81",
          1137 => x"71",
          1138 => x"38",
          1139 => x"be",
          1140 => x"a8",
          1141 => x"3f",
          1142 => x"b2",
          1143 => x"2a",
          1144 => x"51",
          1145 => x"2e",
          1146 => x"51",
          1147 => x"81",
          1148 => x"9b",
          1149 => x"51",
          1150 => x"a7",
          1151 => x"3d",
          1152 => x"3d",
          1153 => x"84",
          1154 => x"33",
          1155 => x"56",
          1156 => x"51",
          1157 => x"0b",
          1158 => x"c8",
          1159 => x"a9",
          1160 => x"81",
          1161 => x"82",
          1162 => x"81",
          1163 => x"82",
          1164 => x"30",
          1165 => x"cc",
          1166 => x"25",
          1167 => x"51",
          1168 => x"0b",
          1169 => x"c8",
          1170 => x"82",
          1171 => x"54",
          1172 => x"09",
          1173 => x"38",
          1174 => x"53",
          1175 => x"51",
          1176 => x"3f",
          1177 => x"08",
          1178 => x"38",
          1179 => x"08",
          1180 => x"3f",
          1181 => x"9e",
          1182 => x"93",
          1183 => x"0b",
          1184 => x"82",
          1185 => x"0b",
          1186 => x"33",
          1187 => x"2e",
          1188 => x"8c",
          1189 => x"8c",
          1190 => x"75",
          1191 => x"3f",
          1192 => x"87",
          1193 => x"3d",
          1194 => x"3d",
          1195 => x"71",
          1196 => x"0c",
          1197 => x"52",
          1198 => x"d5",
          1199 => x"87",
          1200 => x"ff",
          1201 => x"7d",
          1202 => x"06",
          1203 => x"f2",
          1204 => x"3d",
          1205 => x"ac",
          1206 => x"53",
          1207 => x"88",
          1208 => x"84",
          1209 => x"87",
          1210 => x"2e",
          1211 => x"f2",
          1212 => x"b4",
          1213 => x"5f",
          1214 => x"d4",
          1215 => x"3f",
          1216 => x"46",
          1217 => x"52",
          1218 => x"f6",
          1219 => x"ff",
          1220 => x"f3",
          1221 => x"87",
          1222 => x"2b",
          1223 => x"51",
          1224 => x"c1",
          1225 => x"38",
          1226 => x"24",
          1227 => x"78",
          1228 => x"b8",
          1229 => x"24",
          1230 => x"82",
          1231 => x"38",
          1232 => x"8a",
          1233 => x"2e",
          1234 => x"8e",
          1235 => x"84",
          1236 => x"38",
          1237 => x"82",
          1238 => x"d2",
          1239 => x"2e",
          1240 => x"78",
          1241 => x"38",
          1242 => x"83",
          1243 => x"bc",
          1244 => x"38",
          1245 => x"78",
          1246 => x"c1",
          1247 => x"c0",
          1248 => x"38",
          1249 => x"78",
          1250 => x"8d",
          1251 => x"80",
          1252 => x"38",
          1253 => x"2e",
          1254 => x"78",
          1255 => x"92",
          1256 => x"c2",
          1257 => x"38",
          1258 => x"2e",
          1259 => x"8d",
          1260 => x"80",
          1261 => x"b2",
          1262 => x"d4",
          1263 => x"38",
          1264 => x"78",
          1265 => x"8d",
          1266 => x"81",
          1267 => x"38",
          1268 => x"2e",
          1269 => x"78",
          1270 => x"8c",
          1271 => x"ce",
          1272 => x"83",
          1273 => x"38",
          1274 => x"2e",
          1275 => x"8d",
          1276 => x"3d",
          1277 => x"53",
          1278 => x"51",
          1279 => x"82",
          1280 => x"88",
          1281 => x"d8",
          1282 => x"39",
          1283 => x"fc",
          1284 => x"84",
          1285 => x"e2",
          1286 => x"cc",
          1287 => x"88",
          1288 => x"25",
          1289 => x"43",
          1290 => x"05",
          1291 => x"80",
          1292 => x"51",
          1293 => x"3f",
          1294 => x"08",
          1295 => x"59",
          1296 => x"81",
          1297 => x"a3",
          1298 => x"5e",
          1299 => x"81",
          1300 => x"87",
          1301 => x"3d",
          1302 => x"53",
          1303 => x"51",
          1304 => x"82",
          1305 => x"80",
          1306 => x"38",
          1307 => x"52",
          1308 => x"05",
          1309 => x"d6",
          1310 => x"87",
          1311 => x"81",
          1312 => x"8c",
          1313 => x"3d",
          1314 => x"53",
          1315 => x"51",
          1316 => x"82",
          1317 => x"80",
          1318 => x"63",
          1319 => x"d9",
          1320 => x"fe",
          1321 => x"ff",
          1322 => x"aa",
          1323 => x"87",
          1324 => x"38",
          1325 => x"08",
          1326 => x"81",
          1327 => x"79",
          1328 => x"3f",
          1329 => x"05",
          1330 => x"52",
          1331 => x"29",
          1332 => x"05",
          1333 => x"df",
          1334 => x"cc",
          1335 => x"38",
          1336 => x"51",
          1337 => x"81",
          1338 => x"39",
          1339 => x"84",
          1340 => x"89",
          1341 => x"cc",
          1342 => x"ff",
          1343 => x"5b",
          1344 => x"81",
          1345 => x"cc",
          1346 => x"51",
          1347 => x"80",
          1348 => x"3d",
          1349 => x"51",
          1350 => x"82",
          1351 => x"b5",
          1352 => x"05",
          1353 => x"f9",
          1354 => x"cc",
          1355 => x"ff",
          1356 => x"5a",
          1357 => x"82",
          1358 => x"b5",
          1359 => x"05",
          1360 => x"dd",
          1361 => x"f0",
          1362 => x"dc",
          1363 => x"80",
          1364 => x"cc",
          1365 => x"06",
          1366 => x"79",
          1367 => x"f3",
          1368 => x"87",
          1369 => x"2e",
          1370 => x"82",
          1371 => x"51",
          1372 => x"fb",
          1373 => x"3d",
          1374 => x"53",
          1375 => x"51",
          1376 => x"82",
          1377 => x"80",
          1378 => x"38",
          1379 => x"fc",
          1380 => x"84",
          1381 => x"e2",
          1382 => x"cc",
          1383 => x"fa",
          1384 => x"3d",
          1385 => x"53",
          1386 => x"51",
          1387 => x"82",
          1388 => x"86",
          1389 => x"cc",
          1390 => x"f3",
          1391 => x"e1",
          1392 => x"5c",
          1393 => x"27",
          1394 => x"61",
          1395 => x"70",
          1396 => x"0c",
          1397 => x"f5",
          1398 => x"39",
          1399 => x"80",
          1400 => x"84",
          1401 => x"92",
          1402 => x"cc",
          1403 => x"fa",
          1404 => x"3d",
          1405 => x"53",
          1406 => x"51",
          1407 => x"82",
          1408 => x"80",
          1409 => x"38",
          1410 => x"f8",
          1411 => x"84",
          1412 => x"e6",
          1413 => x"cc",
          1414 => x"f9",
          1415 => x"f3",
          1416 => x"fd",
          1417 => x"79",
          1418 => x"87",
          1419 => x"79",
          1420 => x"5b",
          1421 => x"61",
          1422 => x"eb",
          1423 => x"ff",
          1424 => x"ff",
          1425 => x"a7",
          1426 => x"87",
          1427 => x"2e",
          1428 => x"b4",
          1429 => x"11",
          1430 => x"05",
          1431 => x"3f",
          1432 => x"08",
          1433 => x"91",
          1434 => x"fe",
          1435 => x"ff",
          1436 => x"a7",
          1437 => x"87",
          1438 => x"2e",
          1439 => x"81",
          1440 => x"9f",
          1441 => x"5a",
          1442 => x"a7",
          1443 => x"33",
          1444 => x"5a",
          1445 => x"2e",
          1446 => x"55",
          1447 => x"33",
          1448 => x"81",
          1449 => x"a4",
          1450 => x"1a",
          1451 => x"43",
          1452 => x"81",
          1453 => x"82",
          1454 => x"3d",
          1455 => x"53",
          1456 => x"51",
          1457 => x"82",
          1458 => x"80",
          1459 => x"86",
          1460 => x"78",
          1461 => x"38",
          1462 => x"08",
          1463 => x"39",
          1464 => x"33",
          1465 => x"2e",
          1466 => x"85",
          1467 => x"bc",
          1468 => x"ba",
          1469 => x"80",
          1470 => x"82",
          1471 => x"44",
          1472 => x"86",
          1473 => x"78",
          1474 => x"38",
          1475 => x"08",
          1476 => x"82",
          1477 => x"59",
          1478 => x"88",
          1479 => x"90",
          1480 => x"39",
          1481 => x"08",
          1482 => x"44",
          1483 => x"fc",
          1484 => x"84",
          1485 => x"c2",
          1486 => x"cc",
          1487 => x"38",
          1488 => x"33",
          1489 => x"2e",
          1490 => x"85",
          1491 => x"80",
          1492 => x"86",
          1493 => x"78",
          1494 => x"38",
          1495 => x"08",
          1496 => x"82",
          1497 => x"59",
          1498 => x"88",
          1499 => x"84",
          1500 => x"39",
          1501 => x"33",
          1502 => x"2e",
          1503 => x"86",
          1504 => x"99",
          1505 => x"b6",
          1506 => x"80",
          1507 => x"82",
          1508 => x"43",
          1509 => x"86",
          1510 => x"05",
          1511 => x"fe",
          1512 => x"ff",
          1513 => x"a4",
          1514 => x"87",
          1515 => x"2e",
          1516 => x"62",
          1517 => x"88",
          1518 => x"81",
          1519 => x"32",
          1520 => x"72",
          1521 => x"70",
          1522 => x"51",
          1523 => x"80",
          1524 => x"7a",
          1525 => x"38",
          1526 => x"f3",
          1527 => x"c1",
          1528 => x"63",
          1529 => x"62",
          1530 => x"ee",
          1531 => x"f3",
          1532 => x"ad",
          1533 => x"39",
          1534 => x"80",
          1535 => x"84",
          1536 => x"f6",
          1537 => x"cc",
          1538 => x"f5",
          1539 => x"3d",
          1540 => x"53",
          1541 => x"51",
          1542 => x"82",
          1543 => x"80",
          1544 => x"63",
          1545 => x"cb",
          1546 => x"34",
          1547 => x"44",
          1548 => x"fc",
          1549 => x"84",
          1550 => x"be",
          1551 => x"cc",
          1552 => x"f5",
          1553 => x"70",
          1554 => x"81",
          1555 => x"a1",
          1556 => x"f8",
          1557 => x"a2",
          1558 => x"45",
          1559 => x"78",
          1560 => x"95",
          1561 => x"27",
          1562 => x"3d",
          1563 => x"53",
          1564 => x"51",
          1565 => x"82",
          1566 => x"80",
          1567 => x"63",
          1568 => x"cb",
          1569 => x"34",
          1570 => x"44",
          1571 => x"81",
          1572 => x"9b",
          1573 => x"ae",
          1574 => x"fe",
          1575 => x"ff",
          1576 => x"a4",
          1577 => x"87",
          1578 => x"2e",
          1579 => x"b4",
          1580 => x"11",
          1581 => x"05",
          1582 => x"3f",
          1583 => x"08",
          1584 => x"38",
          1585 => x"be",
          1586 => x"70",
          1587 => x"23",
          1588 => x"3d",
          1589 => x"53",
          1590 => x"51",
          1591 => x"82",
          1592 => x"e0",
          1593 => x"39",
          1594 => x"54",
          1595 => x"94",
          1596 => x"3f",
          1597 => x"79",
          1598 => x"3f",
          1599 => x"33",
          1600 => x"2e",
          1601 => x"78",
          1602 => x"38",
          1603 => x"41",
          1604 => x"3d",
          1605 => x"53",
          1606 => x"51",
          1607 => x"82",
          1608 => x"80",
          1609 => x"60",
          1610 => x"05",
          1611 => x"82",
          1612 => x"78",
          1613 => x"39",
          1614 => x"51",
          1615 => x"ff",
          1616 => x"3d",
          1617 => x"53",
          1618 => x"51",
          1619 => x"82",
          1620 => x"80",
          1621 => x"38",
          1622 => x"f0",
          1623 => x"84",
          1624 => x"88",
          1625 => x"cc",
          1626 => x"a0",
          1627 => x"71",
          1628 => x"84",
          1629 => x"3d",
          1630 => x"53",
          1631 => x"51",
          1632 => x"82",
          1633 => x"e5",
          1634 => x"39",
          1635 => x"54",
          1636 => x"a0",
          1637 => x"3f",
          1638 => x"79",
          1639 => x"3f",
          1640 => x"33",
          1641 => x"2e",
          1642 => x"9f",
          1643 => x"38",
          1644 => x"f0",
          1645 => x"84",
          1646 => x"b0",
          1647 => x"cc",
          1648 => x"8d",
          1649 => x"71",
          1650 => x"84",
          1651 => x"bc",
          1652 => x"8c",
          1653 => x"3f",
          1654 => x"81",
          1655 => x"98",
          1656 => x"51",
          1657 => x"f2",
          1658 => x"f4",
          1659 => x"b1",
          1660 => x"96",
          1661 => x"81",
          1662 => x"dc",
          1663 => x"3f",
          1664 => x"0b",
          1665 => x"84",
          1666 => x"81",
          1667 => x"94",
          1668 => x"e5",
          1669 => x"f0",
          1670 => x"3f",
          1671 => x"0b",
          1672 => x"84",
          1673 => x"83",
          1674 => x"94",
          1675 => x"c9",
          1676 => x"ff",
          1677 => x"ff",
          1678 => x"9f",
          1679 => x"87",
          1680 => x"2e",
          1681 => x"63",
          1682 => x"84",
          1683 => x"3f",
          1684 => x"04",
          1685 => x"80",
          1686 => x"84",
          1687 => x"9a",
          1688 => x"cc",
          1689 => x"f1",
          1690 => x"52",
          1691 => x"51",
          1692 => x"63",
          1693 => x"82",
          1694 => x"80",
          1695 => x"38",
          1696 => x"08",
          1697 => x"bc",
          1698 => x"3f",
          1699 => x"81",
          1700 => x"97",
          1701 => x"82",
          1702 => x"39",
          1703 => x"51",
          1704 => x"80",
          1705 => x"39",
          1706 => x"f0",
          1707 => x"45",
          1708 => x"78",
          1709 => x"c1",
          1710 => x"06",
          1711 => x"2e",
          1712 => x"b4",
          1713 => x"05",
          1714 => x"3f",
          1715 => x"08",
          1716 => x"7b",
          1717 => x"38",
          1718 => x"89",
          1719 => x"2e",
          1720 => x"ca",
          1721 => x"2e",
          1722 => x"c2",
          1723 => x"88",
          1724 => x"81",
          1725 => x"80",
          1726 => x"90",
          1727 => x"ff",
          1728 => x"9c",
          1729 => x"39",
          1730 => x"52",
          1731 => x"b0",
          1732 => x"87",
          1733 => x"7a",
          1734 => x"8c",
          1735 => x"81",
          1736 => x"b4",
          1737 => x"05",
          1738 => x"3f",
          1739 => x"54",
          1740 => x"f6",
          1741 => x"3d",
          1742 => x"51",
          1743 => x"82",
          1744 => x"82",
          1745 => x"80",
          1746 => x"80",
          1747 => x"80",
          1748 => x"80",
          1749 => x"ff",
          1750 => x"e7",
          1751 => x"87",
          1752 => x"87",
          1753 => x"70",
          1754 => x"07",
          1755 => x"5b",
          1756 => x"5a",
          1757 => x"83",
          1758 => x"78",
          1759 => x"78",
          1760 => x"38",
          1761 => x"81",
          1762 => x"59",
          1763 => x"38",
          1764 => x"7d",
          1765 => x"59",
          1766 => x"7e",
          1767 => x"81",
          1768 => x"38",
          1769 => x"51",
          1770 => x"ee",
          1771 => x"3d",
          1772 => x"82",
          1773 => x"87",
          1774 => x"70",
          1775 => x"87",
          1776 => x"72",
          1777 => x"3f",
          1778 => x"08",
          1779 => x"08",
          1780 => x"84",
          1781 => x"51",
          1782 => x"72",
          1783 => x"08",
          1784 => x"87",
          1785 => x"70",
          1786 => x"87",
          1787 => x"72",
          1788 => x"3f",
          1789 => x"08",
          1790 => x"08",
          1791 => x"84",
          1792 => x"51",
          1793 => x"72",
          1794 => x"08",
          1795 => x"8c",
          1796 => x"87",
          1797 => x"0c",
          1798 => x"0b",
          1799 => x"94",
          1800 => x"0b",
          1801 => x"0c",
          1802 => x"0b",
          1803 => x"0c",
          1804 => x"92",
          1805 => x"f6",
          1806 => x"e5",
          1807 => x"d0",
          1808 => x"3f",
          1809 => x"92",
          1810 => x"51",
          1811 => x"ec",
          1812 => x"04",
          1813 => x"80",
          1814 => x"71",
          1815 => x"87",
          1816 => x"87",
          1817 => x"ff",
          1818 => x"ff",
          1819 => x"72",
          1820 => x"38",
          1821 => x"cc",
          1822 => x"0d",
          1823 => x"0d",
          1824 => x"54",
          1825 => x"52",
          1826 => x"2e",
          1827 => x"72",
          1828 => x"a0",
          1829 => x"06",
          1830 => x"13",
          1831 => x"72",
          1832 => x"a2",
          1833 => x"06",
          1834 => x"13",
          1835 => x"72",
          1836 => x"2e",
          1837 => x"9f",
          1838 => x"81",
          1839 => x"72",
          1840 => x"70",
          1841 => x"38",
          1842 => x"80",
          1843 => x"73",
          1844 => x"39",
          1845 => x"80",
          1846 => x"54",
          1847 => x"83",
          1848 => x"70",
          1849 => x"38",
          1850 => x"80",
          1851 => x"54",
          1852 => x"09",
          1853 => x"38",
          1854 => x"a2",
          1855 => x"70",
          1856 => x"07",
          1857 => x"70",
          1858 => x"38",
          1859 => x"81",
          1860 => x"71",
          1861 => x"51",
          1862 => x"cc",
          1863 => x"0d",
          1864 => x"0d",
          1865 => x"08",
          1866 => x"38",
          1867 => x"05",
          1868 => x"9b",
          1869 => x"87",
          1870 => x"38",
          1871 => x"39",
          1872 => x"82",
          1873 => x"86",
          1874 => x"fc",
          1875 => x"82",
          1876 => x"05",
          1877 => x"52",
          1878 => x"81",
          1879 => x"13",
          1880 => x"51",
          1881 => x"9e",
          1882 => x"38",
          1883 => x"51",
          1884 => x"97",
          1885 => x"38",
          1886 => x"51",
          1887 => x"bb",
          1888 => x"38",
          1889 => x"51",
          1890 => x"bb",
          1891 => x"38",
          1892 => x"55",
          1893 => x"87",
          1894 => x"d9",
          1895 => x"22",
          1896 => x"73",
          1897 => x"80",
          1898 => x"0b",
          1899 => x"9c",
          1900 => x"87",
          1901 => x"0c",
          1902 => x"87",
          1903 => x"0c",
          1904 => x"87",
          1905 => x"0c",
          1906 => x"87",
          1907 => x"0c",
          1908 => x"87",
          1909 => x"0c",
          1910 => x"87",
          1911 => x"0c",
          1912 => x"98",
          1913 => x"87",
          1914 => x"0c",
          1915 => x"c0",
          1916 => x"80",
          1917 => x"87",
          1918 => x"3d",
          1919 => x"3d",
          1920 => x"87",
          1921 => x"5d",
          1922 => x"87",
          1923 => x"08",
          1924 => x"23",
          1925 => x"b8",
          1926 => x"82",
          1927 => x"c0",
          1928 => x"5a",
          1929 => x"34",
          1930 => x"b0",
          1931 => x"84",
          1932 => x"c0",
          1933 => x"5a",
          1934 => x"34",
          1935 => x"a8",
          1936 => x"86",
          1937 => x"c0",
          1938 => x"5c",
          1939 => x"23",
          1940 => x"a0",
          1941 => x"8a",
          1942 => x"7d",
          1943 => x"ff",
          1944 => x"7b",
          1945 => x"06",
          1946 => x"33",
          1947 => x"33",
          1948 => x"33",
          1949 => x"33",
          1950 => x"33",
          1951 => x"ff",
          1952 => x"81",
          1953 => x"94",
          1954 => x"3d",
          1955 => x"3d",
          1956 => x"05",
          1957 => x"70",
          1958 => x"52",
          1959 => x"85",
          1960 => x"3d",
          1961 => x"3d",
          1962 => x"85",
          1963 => x"81",
          1964 => x"55",
          1965 => x"94",
          1966 => x"80",
          1967 => x"87",
          1968 => x"51",
          1969 => x"96",
          1970 => x"06",
          1971 => x"70",
          1972 => x"38",
          1973 => x"70",
          1974 => x"51",
          1975 => x"72",
          1976 => x"81",
          1977 => x"70",
          1978 => x"38",
          1979 => x"70",
          1980 => x"51",
          1981 => x"38",
          1982 => x"06",
          1983 => x"94",
          1984 => x"80",
          1985 => x"87",
          1986 => x"52",
          1987 => x"75",
          1988 => x"0c",
          1989 => x"04",
          1990 => x"02",
          1991 => x"82",
          1992 => x"70",
          1993 => x"57",
          1994 => x"c0",
          1995 => x"74",
          1996 => x"38",
          1997 => x"94",
          1998 => x"70",
          1999 => x"81",
          2000 => x"52",
          2001 => x"8c",
          2002 => x"2a",
          2003 => x"51",
          2004 => x"38",
          2005 => x"70",
          2006 => x"51",
          2007 => x"8d",
          2008 => x"2a",
          2009 => x"51",
          2010 => x"be",
          2011 => x"ff",
          2012 => x"c0",
          2013 => x"70",
          2014 => x"38",
          2015 => x"90",
          2016 => x"0c",
          2017 => x"04",
          2018 => x"79",
          2019 => x"33",
          2020 => x"06",
          2021 => x"70",
          2022 => x"fc",
          2023 => x"ff",
          2024 => x"82",
          2025 => x"70",
          2026 => x"59",
          2027 => x"87",
          2028 => x"51",
          2029 => x"86",
          2030 => x"94",
          2031 => x"08",
          2032 => x"70",
          2033 => x"54",
          2034 => x"2e",
          2035 => x"91",
          2036 => x"06",
          2037 => x"d7",
          2038 => x"32",
          2039 => x"51",
          2040 => x"2e",
          2041 => x"93",
          2042 => x"06",
          2043 => x"ff",
          2044 => x"81",
          2045 => x"87",
          2046 => x"52",
          2047 => x"86",
          2048 => x"94",
          2049 => x"72",
          2050 => x"74",
          2051 => x"ff",
          2052 => x"57",
          2053 => x"38",
          2054 => x"cc",
          2055 => x"0d",
          2056 => x"0d",
          2057 => x"33",
          2058 => x"06",
          2059 => x"c0",
          2060 => x"72",
          2061 => x"38",
          2062 => x"94",
          2063 => x"70",
          2064 => x"81",
          2065 => x"51",
          2066 => x"e2",
          2067 => x"ff",
          2068 => x"c0",
          2069 => x"70",
          2070 => x"38",
          2071 => x"90",
          2072 => x"70",
          2073 => x"82",
          2074 => x"51",
          2075 => x"04",
          2076 => x"82",
          2077 => x"70",
          2078 => x"52",
          2079 => x"94",
          2080 => x"80",
          2081 => x"87",
          2082 => x"52",
          2083 => x"82",
          2084 => x"06",
          2085 => x"ff",
          2086 => x"2e",
          2087 => x"81",
          2088 => x"87",
          2089 => x"52",
          2090 => x"86",
          2091 => x"94",
          2092 => x"08",
          2093 => x"70",
          2094 => x"53",
          2095 => x"87",
          2096 => x"3d",
          2097 => x"3d",
          2098 => x"9e",
          2099 => x"9c",
          2100 => x"51",
          2101 => x"2e",
          2102 => x"87",
          2103 => x"08",
          2104 => x"0c",
          2105 => x"a8",
          2106 => x"f4",
          2107 => x"9e",
          2108 => x"85",
          2109 => x"c0",
          2110 => x"82",
          2111 => x"87",
          2112 => x"08",
          2113 => x"0c",
          2114 => x"a0",
          2115 => x"84",
          2116 => x"9e",
          2117 => x"86",
          2118 => x"c0",
          2119 => x"82",
          2120 => x"87",
          2121 => x"08",
          2122 => x"0c",
          2123 => x"b8",
          2124 => x"94",
          2125 => x"9e",
          2126 => x"86",
          2127 => x"c0",
          2128 => x"82",
          2129 => x"87",
          2130 => x"08",
          2131 => x"0c",
          2132 => x"80",
          2133 => x"82",
          2134 => x"87",
          2135 => x"08",
          2136 => x"0c",
          2137 => x"88",
          2138 => x"ac",
          2139 => x"9e",
          2140 => x"86",
          2141 => x"0b",
          2142 => x"34",
          2143 => x"c0",
          2144 => x"70",
          2145 => x"06",
          2146 => x"70",
          2147 => x"38",
          2148 => x"82",
          2149 => x"80",
          2150 => x"9e",
          2151 => x"88",
          2152 => x"51",
          2153 => x"80",
          2154 => x"81",
          2155 => x"86",
          2156 => x"0b",
          2157 => x"90",
          2158 => x"80",
          2159 => x"52",
          2160 => x"2e",
          2161 => x"52",
          2162 => x"b7",
          2163 => x"87",
          2164 => x"08",
          2165 => x"80",
          2166 => x"52",
          2167 => x"83",
          2168 => x"71",
          2169 => x"34",
          2170 => x"c0",
          2171 => x"70",
          2172 => x"06",
          2173 => x"70",
          2174 => x"38",
          2175 => x"82",
          2176 => x"80",
          2177 => x"9e",
          2178 => x"90",
          2179 => x"51",
          2180 => x"80",
          2181 => x"81",
          2182 => x"86",
          2183 => x"0b",
          2184 => x"90",
          2185 => x"80",
          2186 => x"52",
          2187 => x"2e",
          2188 => x"52",
          2189 => x"bb",
          2190 => x"87",
          2191 => x"08",
          2192 => x"80",
          2193 => x"52",
          2194 => x"83",
          2195 => x"71",
          2196 => x"34",
          2197 => x"c0",
          2198 => x"70",
          2199 => x"06",
          2200 => x"70",
          2201 => x"38",
          2202 => x"82",
          2203 => x"80",
          2204 => x"9e",
          2205 => x"80",
          2206 => x"51",
          2207 => x"80",
          2208 => x"81",
          2209 => x"86",
          2210 => x"0b",
          2211 => x"90",
          2212 => x"80",
          2213 => x"52",
          2214 => x"83",
          2215 => x"71",
          2216 => x"34",
          2217 => x"90",
          2218 => x"80",
          2219 => x"2a",
          2220 => x"70",
          2221 => x"34",
          2222 => x"c0",
          2223 => x"70",
          2224 => x"51",
          2225 => x"80",
          2226 => x"81",
          2227 => x"86",
          2228 => x"c0",
          2229 => x"70",
          2230 => x"70",
          2231 => x"51",
          2232 => x"86",
          2233 => x"0b",
          2234 => x"90",
          2235 => x"06",
          2236 => x"70",
          2237 => x"38",
          2238 => x"82",
          2239 => x"87",
          2240 => x"08",
          2241 => x"51",
          2242 => x"86",
          2243 => x"3d",
          2244 => x"3d",
          2245 => x"80",
          2246 => x"3f",
          2247 => x"33",
          2248 => x"2e",
          2249 => x"f7",
          2250 => x"f5",
          2251 => x"a8",
          2252 => x"3f",
          2253 => x"33",
          2254 => x"2e",
          2255 => x"86",
          2256 => x"86",
          2257 => x"54",
          2258 => x"c0",
          2259 => x"3f",
          2260 => x"33",
          2261 => x"2e",
          2262 => x"86",
          2263 => x"86",
          2264 => x"54",
          2265 => x"dc",
          2266 => x"3f",
          2267 => x"33",
          2268 => x"2e",
          2269 => x"85",
          2270 => x"85",
          2271 => x"54",
          2272 => x"f8",
          2273 => x"3f",
          2274 => x"33",
          2275 => x"2e",
          2276 => x"85",
          2277 => x"85",
          2278 => x"54",
          2279 => x"94",
          2280 => x"3f",
          2281 => x"33",
          2282 => x"2e",
          2283 => x"86",
          2284 => x"86",
          2285 => x"54",
          2286 => x"b0",
          2287 => x"3f",
          2288 => x"33",
          2289 => x"2e",
          2290 => x"86",
          2291 => x"81",
          2292 => x"8a",
          2293 => x"86",
          2294 => x"73",
          2295 => x"38",
          2296 => x"33",
          2297 => x"ec",
          2298 => x"3f",
          2299 => x"33",
          2300 => x"2e",
          2301 => x"86",
          2302 => x"81",
          2303 => x"8a",
          2304 => x"86",
          2305 => x"73",
          2306 => x"38",
          2307 => x"51",
          2308 => x"82",
          2309 => x"54",
          2310 => x"88",
          2311 => x"c0",
          2312 => x"3f",
          2313 => x"33",
          2314 => x"2e",
          2315 => x"f9",
          2316 => x"ed",
          2317 => x"bd",
          2318 => x"80",
          2319 => x"81",
          2320 => x"83",
          2321 => x"86",
          2322 => x"73",
          2323 => x"38",
          2324 => x"51",
          2325 => x"81",
          2326 => x"83",
          2327 => x"86",
          2328 => x"81",
          2329 => x"89",
          2330 => x"86",
          2331 => x"81",
          2332 => x"89",
          2333 => x"86",
          2334 => x"81",
          2335 => x"89",
          2336 => x"fa",
          2337 => x"99",
          2338 => x"a4",
          2339 => x"fa",
          2340 => x"f1",
          2341 => x"a8",
          2342 => x"84",
          2343 => x"51",
          2344 => x"82",
          2345 => x"bd",
          2346 => x"76",
          2347 => x"54",
          2348 => x"08",
          2349 => x"a4",
          2350 => x"3f",
          2351 => x"33",
          2352 => x"2e",
          2353 => x"86",
          2354 => x"bd",
          2355 => x"75",
          2356 => x"3f",
          2357 => x"08",
          2358 => x"29",
          2359 => x"54",
          2360 => x"cc",
          2361 => x"fb",
          2362 => x"99",
          2363 => x"b6",
          2364 => x"80",
          2365 => x"82",
          2366 => x"56",
          2367 => x"52",
          2368 => x"e8",
          2369 => x"cc",
          2370 => x"c0",
          2371 => x"31",
          2372 => x"87",
          2373 => x"81",
          2374 => x"87",
          2375 => x"f2",
          2376 => x"fd",
          2377 => x"0d",
          2378 => x"0d",
          2379 => x"33",
          2380 => x"71",
          2381 => x"38",
          2382 => x"81",
          2383 => x"52",
          2384 => x"81",
          2385 => x"9d",
          2386 => x"b0",
          2387 => x"81",
          2388 => x"91",
          2389 => x"c0",
          2390 => x"81",
          2391 => x"85",
          2392 => x"cc",
          2393 => x"3f",
          2394 => x"04",
          2395 => x"0c",
          2396 => x"0d",
          2397 => x"84",
          2398 => x"52",
          2399 => x"70",
          2400 => x"82",
          2401 => x"72",
          2402 => x"0d",
          2403 => x"0d",
          2404 => x"84",
          2405 => x"86",
          2406 => x"80",
          2407 => x"09",
          2408 => x"c8",
          2409 => x"82",
          2410 => x"73",
          2411 => x"3d",
          2412 => x"0b",
          2413 => x"84",
          2414 => x"86",
          2415 => x"c0",
          2416 => x"04",
          2417 => x"02",
          2418 => x"53",
          2419 => x"09",
          2420 => x"38",
          2421 => x"3f",
          2422 => x"08",
          2423 => x"2e",
          2424 => x"72",
          2425 => x"dc",
          2426 => x"82",
          2427 => x"8f",
          2428 => x"d4",
          2429 => x"80",
          2430 => x"72",
          2431 => x"84",
          2432 => x"fe",
          2433 => x"97",
          2434 => x"9e",
          2435 => x"82",
          2436 => x"54",
          2437 => x"3f",
          2438 => x"d4",
          2439 => x"0d",
          2440 => x"0d",
          2441 => x"33",
          2442 => x"06",
          2443 => x"80",
          2444 => x"72",
          2445 => x"51",
          2446 => x"ff",
          2447 => x"39",
          2448 => x"04",
          2449 => x"77",
          2450 => x"08",
          2451 => x"d4",
          2452 => x"73",
          2453 => x"ff",
          2454 => x"71",
          2455 => x"38",
          2456 => x"06",
          2457 => x"54",
          2458 => x"e7",
          2459 => x"9e",
          2460 => x"3d",
          2461 => x"3d",
          2462 => x"59",
          2463 => x"81",
          2464 => x"56",
          2465 => x"84",
          2466 => x"a5",
          2467 => x"06",
          2468 => x"80",
          2469 => x"81",
          2470 => x"58",
          2471 => x"b0",
          2472 => x"06",
          2473 => x"5a",
          2474 => x"ad",
          2475 => x"06",
          2476 => x"5a",
          2477 => x"05",
          2478 => x"75",
          2479 => x"81",
          2480 => x"77",
          2481 => x"08",
          2482 => x"05",
          2483 => x"5d",
          2484 => x"39",
          2485 => x"72",
          2486 => x"38",
          2487 => x"7b",
          2488 => x"05",
          2489 => x"70",
          2490 => x"33",
          2491 => x"39",
          2492 => x"32",
          2493 => x"72",
          2494 => x"78",
          2495 => x"70",
          2496 => x"07",
          2497 => x"07",
          2498 => x"51",
          2499 => x"80",
          2500 => x"79",
          2501 => x"70",
          2502 => x"33",
          2503 => x"80",
          2504 => x"38",
          2505 => x"e0",
          2506 => x"38",
          2507 => x"81",
          2508 => x"53",
          2509 => x"2e",
          2510 => x"73",
          2511 => x"a2",
          2512 => x"c3",
          2513 => x"38",
          2514 => x"24",
          2515 => x"80",
          2516 => x"8c",
          2517 => x"39",
          2518 => x"2e",
          2519 => x"81",
          2520 => x"80",
          2521 => x"80",
          2522 => x"d5",
          2523 => x"73",
          2524 => x"8e",
          2525 => x"39",
          2526 => x"2e",
          2527 => x"80",
          2528 => x"84",
          2529 => x"56",
          2530 => x"74",
          2531 => x"72",
          2532 => x"38",
          2533 => x"15",
          2534 => x"54",
          2535 => x"38",
          2536 => x"56",
          2537 => x"81",
          2538 => x"72",
          2539 => x"38",
          2540 => x"90",
          2541 => x"06",
          2542 => x"2e",
          2543 => x"51",
          2544 => x"74",
          2545 => x"53",
          2546 => x"fd",
          2547 => x"51",
          2548 => x"ef",
          2549 => x"19",
          2550 => x"53",
          2551 => x"39",
          2552 => x"39",
          2553 => x"39",
          2554 => x"39",
          2555 => x"39",
          2556 => x"d0",
          2557 => x"39",
          2558 => x"70",
          2559 => x"53",
          2560 => x"88",
          2561 => x"19",
          2562 => x"39",
          2563 => x"54",
          2564 => x"74",
          2565 => x"70",
          2566 => x"07",
          2567 => x"55",
          2568 => x"80",
          2569 => x"72",
          2570 => x"38",
          2571 => x"90",
          2572 => x"80",
          2573 => x"5e",
          2574 => x"74",
          2575 => x"3f",
          2576 => x"08",
          2577 => x"7c",
          2578 => x"54",
          2579 => x"82",
          2580 => x"55",
          2581 => x"92",
          2582 => x"53",
          2583 => x"2e",
          2584 => x"14",
          2585 => x"ff",
          2586 => x"14",
          2587 => x"70",
          2588 => x"34",
          2589 => x"30",
          2590 => x"9f",
          2591 => x"57",
          2592 => x"85",
          2593 => x"b1",
          2594 => x"2a",
          2595 => x"51",
          2596 => x"2e",
          2597 => x"3d",
          2598 => x"05",
          2599 => x"34",
          2600 => x"76",
          2601 => x"54",
          2602 => x"72",
          2603 => x"54",
          2604 => x"70",
          2605 => x"56",
          2606 => x"81",
          2607 => x"7b",
          2608 => x"73",
          2609 => x"3f",
          2610 => x"53",
          2611 => x"74",
          2612 => x"53",
          2613 => x"eb",
          2614 => x"77",
          2615 => x"53",
          2616 => x"14",
          2617 => x"54",
          2618 => x"3f",
          2619 => x"74",
          2620 => x"53",
          2621 => x"fb",
          2622 => x"51",
          2623 => x"ef",
          2624 => x"0d",
          2625 => x"0d",
          2626 => x"70",
          2627 => x"08",
          2628 => x"51",
          2629 => x"85",
          2630 => x"fe",
          2631 => x"82",
          2632 => x"85",
          2633 => x"52",
          2634 => x"ca",
          2635 => x"dc",
          2636 => x"73",
          2637 => x"82",
          2638 => x"84",
          2639 => x"fd",
          2640 => x"9e",
          2641 => x"82",
          2642 => x"87",
          2643 => x"53",
          2644 => x"fa",
          2645 => x"82",
          2646 => x"85",
          2647 => x"fb",
          2648 => x"79",
          2649 => x"08",
          2650 => x"57",
          2651 => x"71",
          2652 => x"e0",
          2653 => x"d8",
          2654 => x"2d",
          2655 => x"08",
          2656 => x"53",
          2657 => x"80",
          2658 => x"8d",
          2659 => x"72",
          2660 => x"30",
          2661 => x"51",
          2662 => x"80",
          2663 => x"71",
          2664 => x"38",
          2665 => x"97",
          2666 => x"25",
          2667 => x"16",
          2668 => x"25",
          2669 => x"14",
          2670 => x"34",
          2671 => x"72",
          2672 => x"3f",
          2673 => x"73",
          2674 => x"72",
          2675 => x"f7",
          2676 => x"53",
          2677 => x"cc",
          2678 => x"0d",
          2679 => x"0d",
          2680 => x"08",
          2681 => x"d8",
          2682 => x"76",
          2683 => x"ef",
          2684 => x"9e",
          2685 => x"3d",
          2686 => x"3d",
          2687 => x"5a",
          2688 => x"7a",
          2689 => x"08",
          2690 => x"53",
          2691 => x"09",
          2692 => x"38",
          2693 => x"0c",
          2694 => x"ad",
          2695 => x"06",
          2696 => x"76",
          2697 => x"0c",
          2698 => x"33",
          2699 => x"73",
          2700 => x"81",
          2701 => x"38",
          2702 => x"05",
          2703 => x"08",
          2704 => x"53",
          2705 => x"2e",
          2706 => x"57",
          2707 => x"2e",
          2708 => x"39",
          2709 => x"13",
          2710 => x"08",
          2711 => x"53",
          2712 => x"55",
          2713 => x"80",
          2714 => x"14",
          2715 => x"88",
          2716 => x"27",
          2717 => x"eb",
          2718 => x"53",
          2719 => x"89",
          2720 => x"38",
          2721 => x"55",
          2722 => x"8a",
          2723 => x"a0",
          2724 => x"c2",
          2725 => x"74",
          2726 => x"e0",
          2727 => x"ff",
          2728 => x"d0",
          2729 => x"ff",
          2730 => x"90",
          2731 => x"38",
          2732 => x"81",
          2733 => x"53",
          2734 => x"ca",
          2735 => x"27",
          2736 => x"77",
          2737 => x"08",
          2738 => x"0c",
          2739 => x"33",
          2740 => x"ff",
          2741 => x"80",
          2742 => x"74",
          2743 => x"79",
          2744 => x"74",
          2745 => x"0c",
          2746 => x"04",
          2747 => x"7a",
          2748 => x"80",
          2749 => x"58",
          2750 => x"33",
          2751 => x"a0",
          2752 => x"06",
          2753 => x"13",
          2754 => x"39",
          2755 => x"09",
          2756 => x"38",
          2757 => x"11",
          2758 => x"08",
          2759 => x"54",
          2760 => x"2e",
          2761 => x"80",
          2762 => x"08",
          2763 => x"0c",
          2764 => x"33",
          2765 => x"80",
          2766 => x"38",
          2767 => x"80",
          2768 => x"38",
          2769 => x"57",
          2770 => x"0c",
          2771 => x"33",
          2772 => x"39",
          2773 => x"74",
          2774 => x"38",
          2775 => x"80",
          2776 => x"89",
          2777 => x"38",
          2778 => x"d0",
          2779 => x"55",
          2780 => x"80",
          2781 => x"39",
          2782 => x"d9",
          2783 => x"80",
          2784 => x"27",
          2785 => x"80",
          2786 => x"89",
          2787 => x"70",
          2788 => x"55",
          2789 => x"70",
          2790 => x"55",
          2791 => x"27",
          2792 => x"14",
          2793 => x"06",
          2794 => x"74",
          2795 => x"73",
          2796 => x"38",
          2797 => x"14",
          2798 => x"05",
          2799 => x"08",
          2800 => x"54",
          2801 => x"39",
          2802 => x"84",
          2803 => x"55",
          2804 => x"81",
          2805 => x"87",
          2806 => x"3d",
          2807 => x"3d",
          2808 => x"2b",
          2809 => x"79",
          2810 => x"98",
          2811 => x"13",
          2812 => x"51",
          2813 => x"51",
          2814 => x"81",
          2815 => x"33",
          2816 => x"74",
          2817 => x"81",
          2818 => x"08",
          2819 => x"05",
          2820 => x"71",
          2821 => x"52",
          2822 => x"09",
          2823 => x"38",
          2824 => x"82",
          2825 => x"85",
          2826 => x"fc",
          2827 => x"02",
          2828 => x"05",
          2829 => x"54",
          2830 => x"80",
          2831 => x"88",
          2832 => x"3f",
          2833 => x"fc",
          2834 => x"f2",
          2835 => x"33",
          2836 => x"71",
          2837 => x"81",
          2838 => x"de",
          2839 => x"f3",
          2840 => x"73",
          2841 => x"0d",
          2842 => x"0d",
          2843 => x"05",
          2844 => x"02",
          2845 => x"05",
          2846 => x"a4",
          2847 => x"29",
          2848 => x"05",
          2849 => x"59",
          2850 => x"59",
          2851 => x"86",
          2852 => x"9e",
          2853 => x"87",
          2854 => x"84",
          2855 => x"cc",
          2856 => x"70",
          2857 => x"5a",
          2858 => x"82",
          2859 => x"75",
          2860 => x"a4",
          2861 => x"29",
          2862 => x"05",
          2863 => x"56",
          2864 => x"2e",
          2865 => x"53",
          2866 => x"51",
          2867 => x"3f",
          2868 => x"33",
          2869 => x"74",
          2870 => x"34",
          2871 => x"06",
          2872 => x"27",
          2873 => x"0b",
          2874 => x"34",
          2875 => x"b6",
          2876 => x"a0",
          2877 => x"80",
          2878 => x"82",
          2879 => x"55",
          2880 => x"8c",
          2881 => x"54",
          2882 => x"52",
          2883 => x"d8",
          2884 => x"87",
          2885 => x"8a",
          2886 => x"f6",
          2887 => x"a0",
          2888 => x"dc",
          2889 => x"3d",
          2890 => x"3d",
          2891 => x"cc",
          2892 => x"72",
          2893 => x"80",
          2894 => x"71",
          2895 => x"3f",
          2896 => x"ff",
          2897 => x"54",
          2898 => x"25",
          2899 => x"0b",
          2900 => x"34",
          2901 => x"08",
          2902 => x"2e",
          2903 => x"51",
          2904 => x"3f",
          2905 => x"08",
          2906 => x"3f",
          2907 => x"87",
          2908 => x"3d",
          2909 => x"3d",
          2910 => x"80",
          2911 => x"a0",
          2912 => x"e2",
          2913 => x"87",
          2914 => x"d2",
          2915 => x"a0",
          2916 => x"f8",
          2917 => x"70",
          2918 => x"8a",
          2919 => x"87",
          2920 => x"2e",
          2921 => x"51",
          2922 => x"3f",
          2923 => x"08",
          2924 => x"82",
          2925 => x"25",
          2926 => x"87",
          2927 => x"05",
          2928 => x"55",
          2929 => x"75",
          2930 => x"81",
          2931 => x"c8",
          2932 => x"b1",
          2933 => x"2e",
          2934 => x"ff",
          2935 => x"3d",
          2936 => x"3d",
          2937 => x"08",
          2938 => x"5a",
          2939 => x"58",
          2940 => x"82",
          2941 => x"51",
          2942 => x"3f",
          2943 => x"08",
          2944 => x"ff",
          2945 => x"a0",
          2946 => x"80",
          2947 => x"3d",
          2948 => x"81",
          2949 => x"82",
          2950 => x"80",
          2951 => x"75",
          2952 => x"94",
          2953 => x"cc",
          2954 => x"58",
          2955 => x"82",
          2956 => x"25",
          2957 => x"87",
          2958 => x"05",
          2959 => x"55",
          2960 => x"74",
          2961 => x"70",
          2962 => x"2a",
          2963 => x"78",
          2964 => x"38",
          2965 => x"38",
          2966 => x"08",
          2967 => x"53",
          2968 => x"b4",
          2969 => x"cc",
          2970 => x"88",
          2971 => x"d4",
          2972 => x"3f",
          2973 => x"09",
          2974 => x"38",
          2975 => x"51",
          2976 => x"3f",
          2977 => x"b6",
          2978 => x"3d",
          2979 => x"87",
          2980 => x"34",
          2981 => x"82",
          2982 => x"a9",
          2983 => x"f6",
          2984 => x"7e",
          2985 => x"72",
          2986 => x"5a",
          2987 => x"2e",
          2988 => x"a2",
          2989 => x"78",
          2990 => x"76",
          2991 => x"81",
          2992 => x"70",
          2993 => x"58",
          2994 => x"2e",
          2995 => x"86",
          2996 => x"26",
          2997 => x"54",
          2998 => x"82",
          2999 => x"70",
          3000 => x"ff",
          3001 => x"82",
          3002 => x"53",
          3003 => x"08",
          3004 => x"d1",
          3005 => x"cc",
          3006 => x"38",
          3007 => x"55",
          3008 => x"88",
          3009 => x"2e",
          3010 => x"39",
          3011 => x"ac",
          3012 => x"5a",
          3013 => x"11",
          3014 => x"51",
          3015 => x"82",
          3016 => x"80",
          3017 => x"ff",
          3018 => x"52",
          3019 => x"b2",
          3020 => x"cc",
          3021 => x"06",
          3022 => x"38",
          3023 => x"39",
          3024 => x"81",
          3025 => x"54",
          3026 => x"ff",
          3027 => x"54",
          3028 => x"cc",
          3029 => x"0d",
          3030 => x"0d",
          3031 => x"b2",
          3032 => x"3d",
          3033 => x"5a",
          3034 => x"3d",
          3035 => x"a4",
          3036 => x"a0",
          3037 => x"73",
          3038 => x"73",
          3039 => x"33",
          3040 => x"83",
          3041 => x"76",
          3042 => x"bb",
          3043 => x"76",
          3044 => x"73",
          3045 => x"ac",
          3046 => x"9b",
          3047 => x"87",
          3048 => x"87",
          3049 => x"87",
          3050 => x"2e",
          3051 => x"93",
          3052 => x"82",
          3053 => x"51",
          3054 => x"3f",
          3055 => x"08",
          3056 => x"38",
          3057 => x"51",
          3058 => x"80",
          3059 => x"87",
          3060 => x"82",
          3061 => x"53",
          3062 => x"90",
          3063 => x"54",
          3064 => x"3f",
          3065 => x"08",
          3066 => x"cc",
          3067 => x"09",
          3068 => x"d0",
          3069 => x"cc",
          3070 => x"b3",
          3071 => x"87",
          3072 => x"80",
          3073 => x"cc",
          3074 => x"38",
          3075 => x"08",
          3076 => x"17",
          3077 => x"74",
          3078 => x"74",
          3079 => x"52",
          3080 => x"c5",
          3081 => x"70",
          3082 => x"5c",
          3083 => x"27",
          3084 => x"5b",
          3085 => x"09",
          3086 => x"97",
          3087 => x"75",
          3088 => x"34",
          3089 => x"82",
          3090 => x"80",
          3091 => x"f9",
          3092 => x"3d",
          3093 => x"3f",
          3094 => x"08",
          3095 => x"98",
          3096 => x"78",
          3097 => x"38",
          3098 => x"06",
          3099 => x"33",
          3100 => x"70",
          3101 => x"9e",
          3102 => x"98",
          3103 => x"2c",
          3104 => x"05",
          3105 => x"81",
          3106 => x"70",
          3107 => x"33",
          3108 => x"51",
          3109 => x"59",
          3110 => x"56",
          3111 => x"80",
          3112 => x"74",
          3113 => x"74",
          3114 => x"29",
          3115 => x"05",
          3116 => x"51",
          3117 => x"24",
          3118 => x"76",
          3119 => x"77",
          3120 => x"3f",
          3121 => x"08",
          3122 => x"54",
          3123 => x"d7",
          3124 => x"9e",
          3125 => x"56",
          3126 => x"81",
          3127 => x"81",
          3128 => x"70",
          3129 => x"81",
          3130 => x"51",
          3131 => x"26",
          3132 => x"53",
          3133 => x"51",
          3134 => x"82",
          3135 => x"81",
          3136 => x"73",
          3137 => x"39",
          3138 => x"80",
          3139 => x"38",
          3140 => x"74",
          3141 => x"34",
          3142 => x"70",
          3143 => x"9e",
          3144 => x"98",
          3145 => x"2c",
          3146 => x"70",
          3147 => x"fc",
          3148 => x"5e",
          3149 => x"57",
          3150 => x"74",
          3151 => x"81",
          3152 => x"38",
          3153 => x"14",
          3154 => x"80",
          3155 => x"e4",
          3156 => x"82",
          3157 => x"92",
          3158 => x"9e",
          3159 => x"82",
          3160 => x"78",
          3161 => x"75",
          3162 => x"54",
          3163 => x"fd",
          3164 => x"84",
          3165 => x"a8",
          3166 => x"08",
          3167 => x"ec",
          3168 => x"7e",
          3169 => x"38",
          3170 => x"33",
          3171 => x"27",
          3172 => x"98",
          3173 => x"2c",
          3174 => x"75",
          3175 => x"74",
          3176 => x"33",
          3177 => x"74",
          3178 => x"29",
          3179 => x"05",
          3180 => x"82",
          3181 => x"56",
          3182 => x"39",
          3183 => x"33",
          3184 => x"54",
          3185 => x"ec",
          3186 => x"54",
          3187 => x"74",
          3188 => x"e8",
          3189 => x"7e",
          3190 => x"81",
          3191 => x"82",
          3192 => x"82",
          3193 => x"70",
          3194 => x"29",
          3195 => x"05",
          3196 => x"82",
          3197 => x"5a",
          3198 => x"74",
          3199 => x"38",
          3200 => x"33",
          3201 => x"bc",
          3202 => x"80",
          3203 => x"80",
          3204 => x"98",
          3205 => x"e8",
          3206 => x"55",
          3207 => x"e0",
          3208 => x"ec",
          3209 => x"2b",
          3210 => x"82",
          3211 => x"5a",
          3212 => x"74",
          3213 => x"9a",
          3214 => x"e7",
          3215 => x"81",
          3216 => x"81",
          3217 => x"70",
          3218 => x"9e",
          3219 => x"51",
          3220 => x"24",
          3221 => x"fa",
          3222 => x"34",
          3223 => x"1b",
          3224 => x"ec",
          3225 => x"81",
          3226 => x"f3",
          3227 => x"df",
          3228 => x"ec",
          3229 => x"ff",
          3230 => x"73",
          3231 => x"d2",
          3232 => x"e8",
          3233 => x"54",
          3234 => x"e8",
          3235 => x"54",
          3236 => x"ec",
          3237 => x"e6",
          3238 => x"9e",
          3239 => x"98",
          3240 => x"2c",
          3241 => x"33",
          3242 => x"57",
          3243 => x"a7",
          3244 => x"54",
          3245 => x"74",
          3246 => x"51",
          3247 => x"74",
          3248 => x"29",
          3249 => x"05",
          3250 => x"82",
          3251 => x"58",
          3252 => x"75",
          3253 => x"a0",
          3254 => x"3f",
          3255 => x"33",
          3256 => x"70",
          3257 => x"9e",
          3258 => x"51",
          3259 => x"74",
          3260 => x"38",
          3261 => x"cc",
          3262 => x"80",
          3263 => x"80",
          3264 => x"98",
          3265 => x"e8",
          3266 => x"55",
          3267 => x"e4",
          3268 => x"39",
          3269 => x"33",
          3270 => x"80",
          3271 => x"51",
          3272 => x"82",
          3273 => x"79",
          3274 => x"3f",
          3275 => x"08",
          3276 => x"54",
          3277 => x"82",
          3278 => x"54",
          3279 => x"8f",
          3280 => x"73",
          3281 => x"f2",
          3282 => x"39",
          3283 => x"80",
          3284 => x"ec",
          3285 => x"82",
          3286 => x"79",
          3287 => x"0c",
          3288 => x"04",
          3289 => x"33",
          3290 => x"2e",
          3291 => x"88",
          3292 => x"3f",
          3293 => x"33",
          3294 => x"73",
          3295 => x"34",
          3296 => x"06",
          3297 => x"82",
          3298 => x"82",
          3299 => x"55",
          3300 => x"2e",
          3301 => x"ff",
          3302 => x"82",
          3303 => x"74",
          3304 => x"98",
          3305 => x"ff",
          3306 => x"55",
          3307 => x"a7",
          3308 => x"54",
          3309 => x"74",
          3310 => x"51",
          3311 => x"74",
          3312 => x"29",
          3313 => x"05",
          3314 => x"82",
          3315 => x"58",
          3316 => x"75",
          3317 => x"a0",
          3318 => x"3f",
          3319 => x"33",
          3320 => x"70",
          3321 => x"9e",
          3322 => x"51",
          3323 => x"74",
          3324 => x"38",
          3325 => x"cc",
          3326 => x"80",
          3327 => x"80",
          3328 => x"98",
          3329 => x"e8",
          3330 => x"55",
          3331 => x"e4",
          3332 => x"39",
          3333 => x"33",
          3334 => x"06",
          3335 => x"33",
          3336 => x"74",
          3337 => x"aa",
          3338 => x"54",
          3339 => x"ec",
          3340 => x"70",
          3341 => x"e3",
          3342 => x"9e",
          3343 => x"81",
          3344 => x"9e",
          3345 => x"56",
          3346 => x"26",
          3347 => x"82",
          3348 => x"ec",
          3349 => x"81",
          3350 => x"ef",
          3351 => x"0b",
          3352 => x"34",
          3353 => x"9e",
          3354 => x"e6",
          3355 => x"38",
          3356 => x"08",
          3357 => x"2e",
          3358 => x"51",
          3359 => x"3f",
          3360 => x"08",
          3361 => x"34",
          3362 => x"08",
          3363 => x"81",
          3364 => x"52",
          3365 => x"ab",
          3366 => x"5b",
          3367 => x"7a",
          3368 => x"86",
          3369 => x"11",
          3370 => x"74",
          3371 => x"38",
          3372 => x"aa",
          3373 => x"87",
          3374 => x"9e",
          3375 => x"87",
          3376 => x"ff",
          3377 => x"53",
          3378 => x"51",
          3379 => x"3f",
          3380 => x"80",
          3381 => x"08",
          3382 => x"2e",
          3383 => x"74",
          3384 => x"d4",
          3385 => x"7a",
          3386 => x"81",
          3387 => x"82",
          3388 => x"55",
          3389 => x"a4",
          3390 => x"ff",
          3391 => x"82",
          3392 => x"82",
          3393 => x"82",
          3394 => x"81",
          3395 => x"05",
          3396 => x"79",
          3397 => x"80",
          3398 => x"39",
          3399 => x"82",
          3400 => x"70",
          3401 => x"74",
          3402 => x"38",
          3403 => x"a9",
          3404 => x"87",
          3405 => x"9e",
          3406 => x"87",
          3407 => x"ff",
          3408 => x"53",
          3409 => x"51",
          3410 => x"3f",
          3411 => x"73",
          3412 => x"5b",
          3413 => x"82",
          3414 => x"74",
          3415 => x"9e",
          3416 => x"9e",
          3417 => x"79",
          3418 => x"3f",
          3419 => x"82",
          3420 => x"70",
          3421 => x"82",
          3422 => x"59",
          3423 => x"77",
          3424 => x"38",
          3425 => x"73",
          3426 => x"34",
          3427 => x"33",
          3428 => x"b0",
          3429 => x"39",
          3430 => x"33",
          3431 => x"2e",
          3432 => x"88",
          3433 => x"3f",
          3434 => x"33",
          3435 => x"73",
          3436 => x"34",
          3437 => x"fb",
          3438 => x"9f",
          3439 => x"2c",
          3440 => x"7a",
          3441 => x"31",
          3442 => x"7d",
          3443 => x"32",
          3444 => x"58",
          3445 => x"55",
          3446 => x"3f",
          3447 => x"08",
          3448 => x"31",
          3449 => x"0c",
          3450 => x"04",
          3451 => x"78",
          3452 => x"a0",
          3453 => x"2e",
          3454 => x"51",
          3455 => x"82",
          3456 => x"52",
          3457 => x"74",
          3458 => x"38",
          3459 => x"e3",
          3460 => x"87",
          3461 => x"53",
          3462 => x"9f",
          3463 => x"38",
          3464 => x"9f",
          3465 => x"38",
          3466 => x"71",
          3467 => x"31",
          3468 => x"58",
          3469 => x"80",
          3470 => x"2e",
          3471 => x"10",
          3472 => x"07",
          3473 => x"07",
          3474 => x"ff",
          3475 => x"70",
          3476 => x"72",
          3477 => x"31",
          3478 => x"56",
          3479 => x"54",
          3480 => x"da",
          3481 => x"76",
          3482 => x"82",
          3483 => x"88",
          3484 => x"fd",
          3485 => x"70",
          3486 => x"06",
          3487 => x"72",
          3488 => x"70",
          3489 => x"71",
          3490 => x"2a",
          3491 => x"83",
          3492 => x"70",
          3493 => x"25",
          3494 => x"71",
          3495 => x"2a",
          3496 => x"05",
          3497 => x"06",
          3498 => x"80",
          3499 => x"84",
          3500 => x"71",
          3501 => x"73",
          3502 => x"06",
          3503 => x"80",
          3504 => x"71",
          3505 => x"2a",
          3506 => x"81",
          3507 => x"06",
          3508 => x"74",
          3509 => x"19",
          3510 => x"cc",
          3511 => x"5f",
          3512 => x"52",
          3513 => x"53",
          3514 => x"51",
          3515 => x"85",
          3516 => x"fd",
          3517 => x"77",
          3518 => x"53",
          3519 => x"b7",
          3520 => x"cc",
          3521 => x"74",
          3522 => x"87",
          3523 => x"85",
          3524 => x"fa",
          3525 => x"7a",
          3526 => x"52",
          3527 => x"8b",
          3528 => x"fe",
          3529 => x"87",
          3530 => x"e0",
          3531 => x"80",
          3532 => x"74",
          3533 => x"3f",
          3534 => x"cc",
          3535 => x"74",
          3536 => x"26",
          3537 => x"80",
          3538 => x"2e",
          3539 => x"81",
          3540 => x"2a",
          3541 => x"77",
          3542 => x"54",
          3543 => x"57",
          3544 => x"a8",
          3545 => x"75",
          3546 => x"75",
          3547 => x"77",
          3548 => x"11",
          3549 => x"81",
          3550 => x"06",
          3551 => x"ff",
          3552 => x"52",
          3553 => x"56",
          3554 => x"38",
          3555 => x"82",
          3556 => x"88",
          3557 => x"f9",
          3558 => x"c0",
          3559 => x"87",
          3560 => x"80",
          3561 => x"c0",
          3562 => x"53",
          3563 => x"c0",
          3564 => x"a9",
          3565 => x"87",
          3566 => x"80",
          3567 => x"34",
          3568 => x"81",
          3569 => x"87",
          3570 => x"77",
          3571 => x"76",
          3572 => x"82",
          3573 => x"54",
          3574 => x"34",
          3575 => x"34",
          3576 => x"08",
          3577 => x"22",
          3578 => x"80",
          3579 => x"83",
          3580 => x"70",
          3581 => x"51",
          3582 => x"88",
          3583 => x"89",
          3584 => x"87",
          3585 => x"88",
          3586 => x"c4",
          3587 => x"11",
          3588 => x"77",
          3589 => x"76",
          3590 => x"89",
          3591 => x"ff",
          3592 => x"52",
          3593 => x"72",
          3594 => x"fb",
          3595 => x"82",
          3596 => x"ff",
          3597 => x"51",
          3598 => x"87",
          3599 => x"3d",
          3600 => x"3d",
          3601 => x"05",
          3602 => x"05",
          3603 => x"71",
          3604 => x"c4",
          3605 => x"2b",
          3606 => x"83",
          3607 => x"70",
          3608 => x"33",
          3609 => x"07",
          3610 => x"ae",
          3611 => x"81",
          3612 => x"07",
          3613 => x"53",
          3614 => x"54",
          3615 => x"53",
          3616 => x"77",
          3617 => x"18",
          3618 => x"c4",
          3619 => x"88",
          3620 => x"70",
          3621 => x"74",
          3622 => x"82",
          3623 => x"70",
          3624 => x"81",
          3625 => x"88",
          3626 => x"83",
          3627 => x"f8",
          3628 => x"56",
          3629 => x"73",
          3630 => x"06",
          3631 => x"54",
          3632 => x"82",
          3633 => x"81",
          3634 => x"72",
          3635 => x"82",
          3636 => x"16",
          3637 => x"34",
          3638 => x"34",
          3639 => x"04",
          3640 => x"82",
          3641 => x"02",
          3642 => x"05",
          3643 => x"2b",
          3644 => x"11",
          3645 => x"33",
          3646 => x"71",
          3647 => x"58",
          3648 => x"55",
          3649 => x"84",
          3650 => x"13",
          3651 => x"2b",
          3652 => x"2a",
          3653 => x"52",
          3654 => x"34",
          3655 => x"34",
          3656 => x"08",
          3657 => x"11",
          3658 => x"33",
          3659 => x"71",
          3660 => x"56",
          3661 => x"72",
          3662 => x"33",
          3663 => x"71",
          3664 => x"70",
          3665 => x"56",
          3666 => x"86",
          3667 => x"87",
          3668 => x"87",
          3669 => x"70",
          3670 => x"33",
          3671 => x"07",
          3672 => x"ff",
          3673 => x"2a",
          3674 => x"53",
          3675 => x"34",
          3676 => x"34",
          3677 => x"04",
          3678 => x"02",
          3679 => x"82",
          3680 => x"71",
          3681 => x"11",
          3682 => x"12",
          3683 => x"2b",
          3684 => x"29",
          3685 => x"81",
          3686 => x"98",
          3687 => x"2b",
          3688 => x"53",
          3689 => x"56",
          3690 => x"71",
          3691 => x"f6",
          3692 => x"fe",
          3693 => x"87",
          3694 => x"16",
          3695 => x"12",
          3696 => x"2b",
          3697 => x"07",
          3698 => x"33",
          3699 => x"71",
          3700 => x"70",
          3701 => x"ff",
          3702 => x"52",
          3703 => x"5a",
          3704 => x"05",
          3705 => x"54",
          3706 => x"13",
          3707 => x"13",
          3708 => x"c4",
          3709 => x"70",
          3710 => x"33",
          3711 => x"71",
          3712 => x"56",
          3713 => x"72",
          3714 => x"81",
          3715 => x"88",
          3716 => x"81",
          3717 => x"70",
          3718 => x"51",
          3719 => x"72",
          3720 => x"81",
          3721 => x"3d",
          3722 => x"3d",
          3723 => x"c4",
          3724 => x"05",
          3725 => x"70",
          3726 => x"11",
          3727 => x"83",
          3728 => x"8b",
          3729 => x"2b",
          3730 => x"59",
          3731 => x"73",
          3732 => x"81",
          3733 => x"88",
          3734 => x"8c",
          3735 => x"22",
          3736 => x"88",
          3737 => x"53",
          3738 => x"73",
          3739 => x"14",
          3740 => x"c4",
          3741 => x"70",
          3742 => x"33",
          3743 => x"71",
          3744 => x"56",
          3745 => x"72",
          3746 => x"33",
          3747 => x"71",
          3748 => x"70",
          3749 => x"55",
          3750 => x"82",
          3751 => x"83",
          3752 => x"87",
          3753 => x"82",
          3754 => x"12",
          3755 => x"2b",
          3756 => x"cc",
          3757 => x"87",
          3758 => x"f7",
          3759 => x"82",
          3760 => x"31",
          3761 => x"83",
          3762 => x"70",
          3763 => x"fd",
          3764 => x"87",
          3765 => x"83",
          3766 => x"82",
          3767 => x"12",
          3768 => x"2b",
          3769 => x"07",
          3770 => x"33",
          3771 => x"71",
          3772 => x"90",
          3773 => x"42",
          3774 => x"5b",
          3775 => x"54",
          3776 => x"8d",
          3777 => x"80",
          3778 => x"fe",
          3779 => x"84",
          3780 => x"33",
          3781 => x"71",
          3782 => x"83",
          3783 => x"11",
          3784 => x"53",
          3785 => x"55",
          3786 => x"34",
          3787 => x"06",
          3788 => x"14",
          3789 => x"c4",
          3790 => x"84",
          3791 => x"13",
          3792 => x"2b",
          3793 => x"2a",
          3794 => x"56",
          3795 => x"16",
          3796 => x"16",
          3797 => x"c4",
          3798 => x"80",
          3799 => x"34",
          3800 => x"14",
          3801 => x"c4",
          3802 => x"84",
          3803 => x"85",
          3804 => x"87",
          3805 => x"70",
          3806 => x"33",
          3807 => x"07",
          3808 => x"80",
          3809 => x"2a",
          3810 => x"56",
          3811 => x"34",
          3812 => x"34",
          3813 => x"04",
          3814 => x"73",
          3815 => x"c4",
          3816 => x"f7",
          3817 => x"80",
          3818 => x"71",
          3819 => x"3f",
          3820 => x"04",
          3821 => x"80",
          3822 => x"f8",
          3823 => x"87",
          3824 => x"ff",
          3825 => x"87",
          3826 => x"11",
          3827 => x"33",
          3828 => x"07",
          3829 => x"56",
          3830 => x"ff",
          3831 => x"78",
          3832 => x"38",
          3833 => x"17",
          3834 => x"12",
          3835 => x"2b",
          3836 => x"ff",
          3837 => x"31",
          3838 => x"ff",
          3839 => x"27",
          3840 => x"56",
          3841 => x"79",
          3842 => x"73",
          3843 => x"38",
          3844 => x"5b",
          3845 => x"85",
          3846 => x"88",
          3847 => x"54",
          3848 => x"78",
          3849 => x"2e",
          3850 => x"79",
          3851 => x"76",
          3852 => x"87",
          3853 => x"70",
          3854 => x"33",
          3855 => x"07",
          3856 => x"ff",
          3857 => x"5a",
          3858 => x"73",
          3859 => x"38",
          3860 => x"54",
          3861 => x"81",
          3862 => x"54",
          3863 => x"81",
          3864 => x"7a",
          3865 => x"06",
          3866 => x"51",
          3867 => x"81",
          3868 => x"80",
          3869 => x"52",
          3870 => x"c6",
          3871 => x"c4",
          3872 => x"86",
          3873 => x"12",
          3874 => x"2b",
          3875 => x"07",
          3876 => x"55",
          3877 => x"17",
          3878 => x"ff",
          3879 => x"2a",
          3880 => x"54",
          3881 => x"34",
          3882 => x"06",
          3883 => x"15",
          3884 => x"c4",
          3885 => x"2b",
          3886 => x"1e",
          3887 => x"87",
          3888 => x"88",
          3889 => x"88",
          3890 => x"5e",
          3891 => x"54",
          3892 => x"34",
          3893 => x"34",
          3894 => x"08",
          3895 => x"11",
          3896 => x"33",
          3897 => x"71",
          3898 => x"53",
          3899 => x"74",
          3900 => x"86",
          3901 => x"87",
          3902 => x"87",
          3903 => x"16",
          3904 => x"11",
          3905 => x"33",
          3906 => x"07",
          3907 => x"53",
          3908 => x"56",
          3909 => x"16",
          3910 => x"16",
          3911 => x"c4",
          3912 => x"05",
          3913 => x"87",
          3914 => x"3d",
          3915 => x"3d",
          3916 => x"82",
          3917 => x"84",
          3918 => x"3f",
          3919 => x"80",
          3920 => x"71",
          3921 => x"3f",
          3922 => x"08",
          3923 => x"87",
          3924 => x"3d",
          3925 => x"3d",
          3926 => x"05",
          3927 => x"52",
          3928 => x"87",
          3929 => x"c8",
          3930 => x"71",
          3931 => x"0c",
          3932 => x"04",
          3933 => x"02",
          3934 => x"02",
          3935 => x"05",
          3936 => x"83",
          3937 => x"26",
          3938 => x"72",
          3939 => x"c0",
          3940 => x"53",
          3941 => x"74",
          3942 => x"38",
          3943 => x"73",
          3944 => x"c0",
          3945 => x"51",
          3946 => x"85",
          3947 => x"98",
          3948 => x"52",
          3949 => x"82",
          3950 => x"70",
          3951 => x"38",
          3952 => x"8c",
          3953 => x"ec",
          3954 => x"fc",
          3955 => x"52",
          3956 => x"87",
          3957 => x"08",
          3958 => x"2e",
          3959 => x"82",
          3960 => x"34",
          3961 => x"13",
          3962 => x"82",
          3963 => x"86",
          3964 => x"f3",
          3965 => x"62",
          3966 => x"05",
          3967 => x"57",
          3968 => x"83",
          3969 => x"fe",
          3970 => x"87",
          3971 => x"06",
          3972 => x"71",
          3973 => x"71",
          3974 => x"2b",
          3975 => x"80",
          3976 => x"92",
          3977 => x"c0",
          3978 => x"41",
          3979 => x"5a",
          3980 => x"87",
          3981 => x"0c",
          3982 => x"84",
          3983 => x"08",
          3984 => x"70",
          3985 => x"53",
          3986 => x"2e",
          3987 => x"08",
          3988 => x"70",
          3989 => x"34",
          3990 => x"80",
          3991 => x"53",
          3992 => x"2e",
          3993 => x"53",
          3994 => x"26",
          3995 => x"80",
          3996 => x"87",
          3997 => x"08",
          3998 => x"38",
          3999 => x"8c",
          4000 => x"80",
          4001 => x"78",
          4002 => x"99",
          4003 => x"0c",
          4004 => x"8c",
          4005 => x"08",
          4006 => x"51",
          4007 => x"38",
          4008 => x"8d",
          4009 => x"17",
          4010 => x"81",
          4011 => x"53",
          4012 => x"2e",
          4013 => x"fc",
          4014 => x"52",
          4015 => x"7d",
          4016 => x"ed",
          4017 => x"80",
          4018 => x"71",
          4019 => x"38",
          4020 => x"53",
          4021 => x"cc",
          4022 => x"0d",
          4023 => x"0d",
          4024 => x"02",
          4025 => x"05",
          4026 => x"58",
          4027 => x"80",
          4028 => x"fc",
          4029 => x"87",
          4030 => x"06",
          4031 => x"71",
          4032 => x"81",
          4033 => x"38",
          4034 => x"2b",
          4035 => x"80",
          4036 => x"92",
          4037 => x"c0",
          4038 => x"40",
          4039 => x"5a",
          4040 => x"c0",
          4041 => x"76",
          4042 => x"76",
          4043 => x"75",
          4044 => x"2a",
          4045 => x"51",
          4046 => x"80",
          4047 => x"7a",
          4048 => x"5c",
          4049 => x"81",
          4050 => x"81",
          4051 => x"06",
          4052 => x"80",
          4053 => x"87",
          4054 => x"08",
          4055 => x"38",
          4056 => x"8c",
          4057 => x"80",
          4058 => x"77",
          4059 => x"99",
          4060 => x"0c",
          4061 => x"8c",
          4062 => x"08",
          4063 => x"51",
          4064 => x"38",
          4065 => x"8d",
          4066 => x"70",
          4067 => x"84",
          4068 => x"5b",
          4069 => x"2e",
          4070 => x"fc",
          4071 => x"52",
          4072 => x"7d",
          4073 => x"f8",
          4074 => x"80",
          4075 => x"71",
          4076 => x"38",
          4077 => x"53",
          4078 => x"cc",
          4079 => x"0d",
          4080 => x"0d",
          4081 => x"05",
          4082 => x"02",
          4083 => x"05",
          4084 => x"54",
          4085 => x"fe",
          4086 => x"cc",
          4087 => x"53",
          4088 => x"80",
          4089 => x"0b",
          4090 => x"8c",
          4091 => x"71",
          4092 => x"dc",
          4093 => x"24",
          4094 => x"84",
          4095 => x"92",
          4096 => x"54",
          4097 => x"8d",
          4098 => x"39",
          4099 => x"80",
          4100 => x"cb",
          4101 => x"70",
          4102 => x"81",
          4103 => x"52",
          4104 => x"8a",
          4105 => x"98",
          4106 => x"71",
          4107 => x"c0",
          4108 => x"52",
          4109 => x"81",
          4110 => x"c0",
          4111 => x"53",
          4112 => x"82",
          4113 => x"71",
          4114 => x"39",
          4115 => x"39",
          4116 => x"77",
          4117 => x"81",
          4118 => x"72",
          4119 => x"84",
          4120 => x"73",
          4121 => x"0c",
          4122 => x"04",
          4123 => x"74",
          4124 => x"71",
          4125 => x"2b",
          4126 => x"cc",
          4127 => x"84",
          4128 => x"fd",
          4129 => x"83",
          4130 => x"12",
          4131 => x"2b",
          4132 => x"07",
          4133 => x"70",
          4134 => x"2b",
          4135 => x"07",
          4136 => x"0c",
          4137 => x"56",
          4138 => x"3d",
          4139 => x"3d",
          4140 => x"84",
          4141 => x"22",
          4142 => x"72",
          4143 => x"54",
          4144 => x"2a",
          4145 => x"34",
          4146 => x"04",
          4147 => x"73",
          4148 => x"70",
          4149 => x"05",
          4150 => x"88",
          4151 => x"72",
          4152 => x"54",
          4153 => x"2a",
          4154 => x"70",
          4155 => x"34",
          4156 => x"51",
          4157 => x"83",
          4158 => x"fe",
          4159 => x"75",
          4160 => x"51",
          4161 => x"92",
          4162 => x"81",
          4163 => x"73",
          4164 => x"55",
          4165 => x"51",
          4166 => x"3d",
          4167 => x"3d",
          4168 => x"76",
          4169 => x"72",
          4170 => x"05",
          4171 => x"11",
          4172 => x"38",
          4173 => x"04",
          4174 => x"78",
          4175 => x"56",
          4176 => x"81",
          4177 => x"74",
          4178 => x"56",
          4179 => x"31",
          4180 => x"52",
          4181 => x"80",
          4182 => x"71",
          4183 => x"38",
          4184 => x"cc",
          4185 => x"0d",
          4186 => x"0d",
          4187 => x"51",
          4188 => x"73",
          4189 => x"81",
          4190 => x"33",
          4191 => x"38",
          4192 => x"87",
          4193 => x"3d",
          4194 => x"0b",
          4195 => x"0c",
          4196 => x"82",
          4197 => x"04",
          4198 => x"7b",
          4199 => x"83",
          4200 => x"5a",
          4201 => x"80",
          4202 => x"54",
          4203 => x"53",
          4204 => x"53",
          4205 => x"52",
          4206 => x"3f",
          4207 => x"08",
          4208 => x"81",
          4209 => x"82",
          4210 => x"83",
          4211 => x"16",
          4212 => x"18",
          4213 => x"18",
          4214 => x"58",
          4215 => x"9f",
          4216 => x"33",
          4217 => x"2e",
          4218 => x"93",
          4219 => x"76",
          4220 => x"52",
          4221 => x"51",
          4222 => x"83",
          4223 => x"79",
          4224 => x"0c",
          4225 => x"04",
          4226 => x"78",
          4227 => x"80",
          4228 => x"17",
          4229 => x"38",
          4230 => x"fc",
          4231 => x"cc",
          4232 => x"87",
          4233 => x"38",
          4234 => x"53",
          4235 => x"81",
          4236 => x"f7",
          4237 => x"87",
          4238 => x"2e",
          4239 => x"55",
          4240 => x"b0",
          4241 => x"82",
          4242 => x"88",
          4243 => x"f8",
          4244 => x"70",
          4245 => x"c0",
          4246 => x"cc",
          4247 => x"87",
          4248 => x"91",
          4249 => x"55",
          4250 => x"09",
          4251 => x"f0",
          4252 => x"33",
          4253 => x"2e",
          4254 => x"80",
          4255 => x"80",
          4256 => x"cc",
          4257 => x"17",
          4258 => x"fd",
          4259 => x"d4",
          4260 => x"b2",
          4261 => x"96",
          4262 => x"85",
          4263 => x"75",
          4264 => x"3f",
          4265 => x"e4",
          4266 => x"98",
          4267 => x"9c",
          4268 => x"08",
          4269 => x"17",
          4270 => x"3f",
          4271 => x"52",
          4272 => x"51",
          4273 => x"a0",
          4274 => x"05",
          4275 => x"0c",
          4276 => x"75",
          4277 => x"33",
          4278 => x"3f",
          4279 => x"34",
          4280 => x"52",
          4281 => x"51",
          4282 => x"82",
          4283 => x"80",
          4284 => x"81",
          4285 => x"87",
          4286 => x"3d",
          4287 => x"3d",
          4288 => x"1a",
          4289 => x"fe",
          4290 => x"54",
          4291 => x"73",
          4292 => x"8a",
          4293 => x"71",
          4294 => x"08",
          4295 => x"75",
          4296 => x"0c",
          4297 => x"04",
          4298 => x"7a",
          4299 => x"56",
          4300 => x"77",
          4301 => x"38",
          4302 => x"08",
          4303 => x"38",
          4304 => x"54",
          4305 => x"2e",
          4306 => x"72",
          4307 => x"38",
          4308 => x"8d",
          4309 => x"39",
          4310 => x"81",
          4311 => x"b6",
          4312 => x"2a",
          4313 => x"2a",
          4314 => x"05",
          4315 => x"55",
          4316 => x"82",
          4317 => x"81",
          4318 => x"83",
          4319 => x"b4",
          4320 => x"17",
          4321 => x"a4",
          4322 => x"55",
          4323 => x"57",
          4324 => x"3f",
          4325 => x"08",
          4326 => x"74",
          4327 => x"14",
          4328 => x"70",
          4329 => x"07",
          4330 => x"71",
          4331 => x"52",
          4332 => x"72",
          4333 => x"75",
          4334 => x"58",
          4335 => x"76",
          4336 => x"15",
          4337 => x"73",
          4338 => x"3f",
          4339 => x"08",
          4340 => x"76",
          4341 => x"06",
          4342 => x"05",
          4343 => x"3f",
          4344 => x"08",
          4345 => x"06",
          4346 => x"76",
          4347 => x"15",
          4348 => x"73",
          4349 => x"3f",
          4350 => x"08",
          4351 => x"82",
          4352 => x"06",
          4353 => x"05",
          4354 => x"3f",
          4355 => x"08",
          4356 => x"58",
          4357 => x"58",
          4358 => x"cc",
          4359 => x"0d",
          4360 => x"0d",
          4361 => x"5a",
          4362 => x"59",
          4363 => x"82",
          4364 => x"98",
          4365 => x"82",
          4366 => x"33",
          4367 => x"2e",
          4368 => x"72",
          4369 => x"38",
          4370 => x"8d",
          4371 => x"39",
          4372 => x"81",
          4373 => x"f7",
          4374 => x"2a",
          4375 => x"2a",
          4376 => x"05",
          4377 => x"55",
          4378 => x"82",
          4379 => x"59",
          4380 => x"08",
          4381 => x"74",
          4382 => x"16",
          4383 => x"16",
          4384 => x"59",
          4385 => x"53",
          4386 => x"8f",
          4387 => x"2b",
          4388 => x"74",
          4389 => x"71",
          4390 => x"72",
          4391 => x"0b",
          4392 => x"74",
          4393 => x"17",
          4394 => x"75",
          4395 => x"3f",
          4396 => x"08",
          4397 => x"cc",
          4398 => x"38",
          4399 => x"06",
          4400 => x"78",
          4401 => x"54",
          4402 => x"77",
          4403 => x"33",
          4404 => x"71",
          4405 => x"51",
          4406 => x"34",
          4407 => x"76",
          4408 => x"17",
          4409 => x"75",
          4410 => x"3f",
          4411 => x"08",
          4412 => x"cc",
          4413 => x"38",
          4414 => x"ff",
          4415 => x"10",
          4416 => x"76",
          4417 => x"51",
          4418 => x"be",
          4419 => x"2a",
          4420 => x"05",
          4421 => x"f9",
          4422 => x"87",
          4423 => x"82",
          4424 => x"ab",
          4425 => x"0a",
          4426 => x"2b",
          4427 => x"70",
          4428 => x"70",
          4429 => x"54",
          4430 => x"82",
          4431 => x"8f",
          4432 => x"07",
          4433 => x"f7",
          4434 => x"0b",
          4435 => x"78",
          4436 => x"0c",
          4437 => x"04",
          4438 => x"7a",
          4439 => x"08",
          4440 => x"59",
          4441 => x"a4",
          4442 => x"17",
          4443 => x"38",
          4444 => x"aa",
          4445 => x"73",
          4446 => x"fd",
          4447 => x"87",
          4448 => x"82",
          4449 => x"80",
          4450 => x"39",
          4451 => x"eb",
          4452 => x"80",
          4453 => x"87",
          4454 => x"80",
          4455 => x"52",
          4456 => x"84",
          4457 => x"cc",
          4458 => x"87",
          4459 => x"2e",
          4460 => x"82",
          4461 => x"81",
          4462 => x"82",
          4463 => x"ff",
          4464 => x"80",
          4465 => x"75",
          4466 => x"3f",
          4467 => x"08",
          4468 => x"16",
          4469 => x"90",
          4470 => x"55",
          4471 => x"27",
          4472 => x"15",
          4473 => x"84",
          4474 => x"07",
          4475 => x"17",
          4476 => x"76",
          4477 => x"a6",
          4478 => x"73",
          4479 => x"0c",
          4480 => x"04",
          4481 => x"7c",
          4482 => x"59",
          4483 => x"95",
          4484 => x"08",
          4485 => x"2e",
          4486 => x"17",
          4487 => x"b2",
          4488 => x"ae",
          4489 => x"7a",
          4490 => x"3f",
          4491 => x"82",
          4492 => x"27",
          4493 => x"82",
          4494 => x"55",
          4495 => x"08",
          4496 => x"d2",
          4497 => x"08",
          4498 => x"08",
          4499 => x"38",
          4500 => x"17",
          4501 => x"54",
          4502 => x"82",
          4503 => x"7a",
          4504 => x"06",
          4505 => x"81",
          4506 => x"17",
          4507 => x"83",
          4508 => x"75",
          4509 => x"f9",
          4510 => x"59",
          4511 => x"08",
          4512 => x"81",
          4513 => x"82",
          4514 => x"59",
          4515 => x"08",
          4516 => x"70",
          4517 => x"25",
          4518 => x"82",
          4519 => x"54",
          4520 => x"55",
          4521 => x"38",
          4522 => x"08",
          4523 => x"38",
          4524 => x"54",
          4525 => x"90",
          4526 => x"18",
          4527 => x"38",
          4528 => x"39",
          4529 => x"38",
          4530 => x"16",
          4531 => x"08",
          4532 => x"38",
          4533 => x"78",
          4534 => x"38",
          4535 => x"51",
          4536 => x"82",
          4537 => x"80",
          4538 => x"80",
          4539 => x"cc",
          4540 => x"09",
          4541 => x"38",
          4542 => x"08",
          4543 => x"cc",
          4544 => x"30",
          4545 => x"80",
          4546 => x"07",
          4547 => x"55",
          4548 => x"38",
          4549 => x"09",
          4550 => x"ae",
          4551 => x"80",
          4552 => x"53",
          4553 => x"51",
          4554 => x"82",
          4555 => x"82",
          4556 => x"30",
          4557 => x"cc",
          4558 => x"25",
          4559 => x"79",
          4560 => x"38",
          4561 => x"8f",
          4562 => x"79",
          4563 => x"f9",
          4564 => x"87",
          4565 => x"74",
          4566 => x"8c",
          4567 => x"17",
          4568 => x"90",
          4569 => x"54",
          4570 => x"86",
          4571 => x"90",
          4572 => x"17",
          4573 => x"54",
          4574 => x"34",
          4575 => x"56",
          4576 => x"90",
          4577 => x"80",
          4578 => x"82",
          4579 => x"55",
          4580 => x"56",
          4581 => x"82",
          4582 => x"8c",
          4583 => x"f8",
          4584 => x"70",
          4585 => x"f0",
          4586 => x"cc",
          4587 => x"56",
          4588 => x"08",
          4589 => x"7b",
          4590 => x"f6",
          4591 => x"87",
          4592 => x"87",
          4593 => x"17",
          4594 => x"80",
          4595 => x"b4",
          4596 => x"57",
          4597 => x"77",
          4598 => x"81",
          4599 => x"15",
          4600 => x"78",
          4601 => x"81",
          4602 => x"53",
          4603 => x"15",
          4604 => x"e9",
          4605 => x"cc",
          4606 => x"df",
          4607 => x"22",
          4608 => x"30",
          4609 => x"70",
          4610 => x"51",
          4611 => x"82",
          4612 => x"8a",
          4613 => x"f8",
          4614 => x"7c",
          4615 => x"56",
          4616 => x"80",
          4617 => x"f1",
          4618 => x"06",
          4619 => x"e9",
          4620 => x"18",
          4621 => x"08",
          4622 => x"38",
          4623 => x"82",
          4624 => x"38",
          4625 => x"54",
          4626 => x"74",
          4627 => x"82",
          4628 => x"22",
          4629 => x"79",
          4630 => x"38",
          4631 => x"98",
          4632 => x"cd",
          4633 => x"22",
          4634 => x"54",
          4635 => x"26",
          4636 => x"52",
          4637 => x"b0",
          4638 => x"cc",
          4639 => x"87",
          4640 => x"2e",
          4641 => x"0b",
          4642 => x"08",
          4643 => x"98",
          4644 => x"87",
          4645 => x"85",
          4646 => x"bd",
          4647 => x"31",
          4648 => x"73",
          4649 => x"f4",
          4650 => x"87",
          4651 => x"18",
          4652 => x"18",
          4653 => x"08",
          4654 => x"72",
          4655 => x"38",
          4656 => x"58",
          4657 => x"89",
          4658 => x"18",
          4659 => x"ff",
          4660 => x"05",
          4661 => x"80",
          4662 => x"87",
          4663 => x"3d",
          4664 => x"3d",
          4665 => x"08",
          4666 => x"a0",
          4667 => x"54",
          4668 => x"77",
          4669 => x"80",
          4670 => x"0c",
          4671 => x"53",
          4672 => x"80",
          4673 => x"38",
          4674 => x"06",
          4675 => x"b5",
          4676 => x"98",
          4677 => x"14",
          4678 => x"92",
          4679 => x"2a",
          4680 => x"56",
          4681 => x"26",
          4682 => x"80",
          4683 => x"16",
          4684 => x"77",
          4685 => x"53",
          4686 => x"38",
          4687 => x"51",
          4688 => x"82",
          4689 => x"53",
          4690 => x"0b",
          4691 => x"08",
          4692 => x"38",
          4693 => x"87",
          4694 => x"2e",
          4695 => x"98",
          4696 => x"87",
          4697 => x"80",
          4698 => x"8a",
          4699 => x"15",
          4700 => x"80",
          4701 => x"14",
          4702 => x"51",
          4703 => x"82",
          4704 => x"53",
          4705 => x"87",
          4706 => x"2e",
          4707 => x"82",
          4708 => x"cc",
          4709 => x"ba",
          4710 => x"82",
          4711 => x"ff",
          4712 => x"82",
          4713 => x"52",
          4714 => x"f3",
          4715 => x"cc",
          4716 => x"72",
          4717 => x"72",
          4718 => x"f2",
          4719 => x"87",
          4720 => x"15",
          4721 => x"15",
          4722 => x"b4",
          4723 => x"0c",
          4724 => x"82",
          4725 => x"8a",
          4726 => x"f7",
          4727 => x"7d",
          4728 => x"5b",
          4729 => x"76",
          4730 => x"3f",
          4731 => x"08",
          4732 => x"cc",
          4733 => x"38",
          4734 => x"08",
          4735 => x"08",
          4736 => x"f0",
          4737 => x"87",
          4738 => x"82",
          4739 => x"80",
          4740 => x"87",
          4741 => x"18",
          4742 => x"51",
          4743 => x"81",
          4744 => x"81",
          4745 => x"81",
          4746 => x"cc",
          4747 => x"83",
          4748 => x"77",
          4749 => x"72",
          4750 => x"38",
          4751 => x"75",
          4752 => x"81",
          4753 => x"a5",
          4754 => x"cc",
          4755 => x"52",
          4756 => x"8e",
          4757 => x"cc",
          4758 => x"87",
          4759 => x"2e",
          4760 => x"73",
          4761 => x"81",
          4762 => x"87",
          4763 => x"87",
          4764 => x"3d",
          4765 => x"3d",
          4766 => x"11",
          4767 => x"ec",
          4768 => x"cc",
          4769 => x"ff",
          4770 => x"33",
          4771 => x"71",
          4772 => x"81",
          4773 => x"94",
          4774 => x"d0",
          4775 => x"cc",
          4776 => x"73",
          4777 => x"82",
          4778 => x"85",
          4779 => x"fc",
          4780 => x"79",
          4781 => x"ff",
          4782 => x"12",
          4783 => x"eb",
          4784 => x"70",
          4785 => x"72",
          4786 => x"81",
          4787 => x"73",
          4788 => x"94",
          4789 => x"d6",
          4790 => x"0d",
          4791 => x"0d",
          4792 => x"55",
          4793 => x"5a",
          4794 => x"08",
          4795 => x"8a",
          4796 => x"08",
          4797 => x"ee",
          4798 => x"87",
          4799 => x"82",
          4800 => x"80",
          4801 => x"15",
          4802 => x"55",
          4803 => x"38",
          4804 => x"e6",
          4805 => x"33",
          4806 => x"70",
          4807 => x"58",
          4808 => x"86",
          4809 => x"87",
          4810 => x"73",
          4811 => x"83",
          4812 => x"73",
          4813 => x"38",
          4814 => x"06",
          4815 => x"80",
          4816 => x"75",
          4817 => x"38",
          4818 => x"08",
          4819 => x"54",
          4820 => x"2e",
          4821 => x"83",
          4822 => x"73",
          4823 => x"38",
          4824 => x"51",
          4825 => x"82",
          4826 => x"58",
          4827 => x"08",
          4828 => x"15",
          4829 => x"38",
          4830 => x"0b",
          4831 => x"77",
          4832 => x"0c",
          4833 => x"04",
          4834 => x"77",
          4835 => x"54",
          4836 => x"51",
          4837 => x"82",
          4838 => x"55",
          4839 => x"08",
          4840 => x"14",
          4841 => x"51",
          4842 => x"82",
          4843 => x"55",
          4844 => x"08",
          4845 => x"53",
          4846 => x"08",
          4847 => x"08",
          4848 => x"3f",
          4849 => x"14",
          4850 => x"08",
          4851 => x"3f",
          4852 => x"17",
          4853 => x"87",
          4854 => x"3d",
          4855 => x"3d",
          4856 => x"08",
          4857 => x"54",
          4858 => x"53",
          4859 => x"82",
          4860 => x"8d",
          4861 => x"08",
          4862 => x"34",
          4863 => x"15",
          4864 => x"0d",
          4865 => x"0d",
          4866 => x"57",
          4867 => x"17",
          4868 => x"08",
          4869 => x"82",
          4870 => x"89",
          4871 => x"55",
          4872 => x"14",
          4873 => x"16",
          4874 => x"71",
          4875 => x"38",
          4876 => x"09",
          4877 => x"38",
          4878 => x"73",
          4879 => x"81",
          4880 => x"ae",
          4881 => x"05",
          4882 => x"15",
          4883 => x"70",
          4884 => x"34",
          4885 => x"8a",
          4886 => x"38",
          4887 => x"05",
          4888 => x"81",
          4889 => x"17",
          4890 => x"12",
          4891 => x"34",
          4892 => x"9c",
          4893 => x"e8",
          4894 => x"87",
          4895 => x"0c",
          4896 => x"e7",
          4897 => x"87",
          4898 => x"17",
          4899 => x"51",
          4900 => x"82",
          4901 => x"84",
          4902 => x"3d",
          4903 => x"3d",
          4904 => x"08",
          4905 => x"61",
          4906 => x"55",
          4907 => x"2e",
          4908 => x"55",
          4909 => x"2e",
          4910 => x"80",
          4911 => x"94",
          4912 => x"1c",
          4913 => x"81",
          4914 => x"61",
          4915 => x"56",
          4916 => x"2e",
          4917 => x"83",
          4918 => x"73",
          4919 => x"70",
          4920 => x"25",
          4921 => x"51",
          4922 => x"38",
          4923 => x"0c",
          4924 => x"51",
          4925 => x"26",
          4926 => x"80",
          4927 => x"34",
          4928 => x"51",
          4929 => x"82",
          4930 => x"55",
          4931 => x"91",
          4932 => x"1d",
          4933 => x"8b",
          4934 => x"79",
          4935 => x"3f",
          4936 => x"57",
          4937 => x"55",
          4938 => x"2e",
          4939 => x"80",
          4940 => x"18",
          4941 => x"1a",
          4942 => x"70",
          4943 => x"2a",
          4944 => x"07",
          4945 => x"5a",
          4946 => x"8c",
          4947 => x"54",
          4948 => x"81",
          4949 => x"39",
          4950 => x"70",
          4951 => x"2a",
          4952 => x"75",
          4953 => x"8c",
          4954 => x"2e",
          4955 => x"a0",
          4956 => x"38",
          4957 => x"0c",
          4958 => x"76",
          4959 => x"38",
          4960 => x"b8",
          4961 => x"70",
          4962 => x"5a",
          4963 => x"76",
          4964 => x"38",
          4965 => x"70",
          4966 => x"dc",
          4967 => x"72",
          4968 => x"80",
          4969 => x"51",
          4970 => x"73",
          4971 => x"38",
          4972 => x"18",
          4973 => x"1a",
          4974 => x"55",
          4975 => x"2e",
          4976 => x"83",
          4977 => x"73",
          4978 => x"70",
          4979 => x"25",
          4980 => x"51",
          4981 => x"38",
          4982 => x"75",
          4983 => x"81",
          4984 => x"81",
          4985 => x"27",
          4986 => x"73",
          4987 => x"38",
          4988 => x"70",
          4989 => x"32",
          4990 => x"80",
          4991 => x"2a",
          4992 => x"56",
          4993 => x"81",
          4994 => x"57",
          4995 => x"f5",
          4996 => x"2b",
          4997 => x"25",
          4998 => x"80",
          4999 => x"81",
          5000 => x"57",
          5001 => x"e6",
          5002 => x"87",
          5003 => x"2e",
          5004 => x"18",
          5005 => x"1a",
          5006 => x"56",
          5007 => x"3f",
          5008 => x"08",
          5009 => x"e8",
          5010 => x"54",
          5011 => x"80",
          5012 => x"17",
          5013 => x"34",
          5014 => x"11",
          5015 => x"74",
          5016 => x"75",
          5017 => x"b4",
          5018 => x"3f",
          5019 => x"08",
          5020 => x"9f",
          5021 => x"99",
          5022 => x"e0",
          5023 => x"ff",
          5024 => x"79",
          5025 => x"74",
          5026 => x"57",
          5027 => x"77",
          5028 => x"76",
          5029 => x"38",
          5030 => x"73",
          5031 => x"09",
          5032 => x"38",
          5033 => x"84",
          5034 => x"27",
          5035 => x"39",
          5036 => x"f2",
          5037 => x"80",
          5038 => x"54",
          5039 => x"34",
          5040 => x"58",
          5041 => x"f2",
          5042 => x"87",
          5043 => x"82",
          5044 => x"80",
          5045 => x"1b",
          5046 => x"51",
          5047 => x"82",
          5048 => x"56",
          5049 => x"08",
          5050 => x"9c",
          5051 => x"33",
          5052 => x"80",
          5053 => x"38",
          5054 => x"bf",
          5055 => x"86",
          5056 => x"15",
          5057 => x"2a",
          5058 => x"51",
          5059 => x"92",
          5060 => x"79",
          5061 => x"e4",
          5062 => x"87",
          5063 => x"2e",
          5064 => x"52",
          5065 => x"ba",
          5066 => x"39",
          5067 => x"33",
          5068 => x"80",
          5069 => x"74",
          5070 => x"81",
          5071 => x"38",
          5072 => x"70",
          5073 => x"82",
          5074 => x"54",
          5075 => x"96",
          5076 => x"06",
          5077 => x"2e",
          5078 => x"ff",
          5079 => x"1c",
          5080 => x"80",
          5081 => x"81",
          5082 => x"ba",
          5083 => x"b6",
          5084 => x"2a",
          5085 => x"51",
          5086 => x"38",
          5087 => x"70",
          5088 => x"81",
          5089 => x"55",
          5090 => x"e1",
          5091 => x"08",
          5092 => x"1d",
          5093 => x"7c",
          5094 => x"3f",
          5095 => x"08",
          5096 => x"fa",
          5097 => x"82",
          5098 => x"8f",
          5099 => x"f6",
          5100 => x"5b",
          5101 => x"70",
          5102 => x"59",
          5103 => x"73",
          5104 => x"c6",
          5105 => x"81",
          5106 => x"70",
          5107 => x"52",
          5108 => x"8d",
          5109 => x"38",
          5110 => x"09",
          5111 => x"a5",
          5112 => x"d0",
          5113 => x"ff",
          5114 => x"53",
          5115 => x"91",
          5116 => x"73",
          5117 => x"d0",
          5118 => x"71",
          5119 => x"f7",
          5120 => x"82",
          5121 => x"55",
          5122 => x"55",
          5123 => x"81",
          5124 => x"74",
          5125 => x"56",
          5126 => x"12",
          5127 => x"70",
          5128 => x"38",
          5129 => x"81",
          5130 => x"51",
          5131 => x"51",
          5132 => x"89",
          5133 => x"70",
          5134 => x"53",
          5135 => x"70",
          5136 => x"51",
          5137 => x"09",
          5138 => x"38",
          5139 => x"38",
          5140 => x"77",
          5141 => x"70",
          5142 => x"2a",
          5143 => x"07",
          5144 => x"51",
          5145 => x"8f",
          5146 => x"84",
          5147 => x"83",
          5148 => x"94",
          5149 => x"74",
          5150 => x"38",
          5151 => x"0c",
          5152 => x"86",
          5153 => x"84",
          5154 => x"82",
          5155 => x"8c",
          5156 => x"fa",
          5157 => x"56",
          5158 => x"17",
          5159 => x"b0",
          5160 => x"52",
          5161 => x"e0",
          5162 => x"82",
          5163 => x"81",
          5164 => x"b2",
          5165 => x"b4",
          5166 => x"cc",
          5167 => x"ff",
          5168 => x"55",
          5169 => x"d5",
          5170 => x"06",
          5171 => x"80",
          5172 => x"33",
          5173 => x"81",
          5174 => x"81",
          5175 => x"81",
          5176 => x"eb",
          5177 => x"70",
          5178 => x"07",
          5179 => x"73",
          5180 => x"81",
          5181 => x"81",
          5182 => x"83",
          5183 => x"c4",
          5184 => x"16",
          5185 => x"3f",
          5186 => x"08",
          5187 => x"cc",
          5188 => x"9d",
          5189 => x"82",
          5190 => x"81",
          5191 => x"e0",
          5192 => x"87",
          5193 => x"82",
          5194 => x"80",
          5195 => x"82",
          5196 => x"87",
          5197 => x"3d",
          5198 => x"3d",
          5199 => x"84",
          5200 => x"05",
          5201 => x"80",
          5202 => x"51",
          5203 => x"82",
          5204 => x"58",
          5205 => x"0b",
          5206 => x"08",
          5207 => x"38",
          5208 => x"08",
          5209 => x"9e",
          5210 => x"08",
          5211 => x"56",
          5212 => x"86",
          5213 => x"75",
          5214 => x"fe",
          5215 => x"54",
          5216 => x"2e",
          5217 => x"14",
          5218 => x"ca",
          5219 => x"cc",
          5220 => x"06",
          5221 => x"54",
          5222 => x"38",
          5223 => x"86",
          5224 => x"82",
          5225 => x"06",
          5226 => x"56",
          5227 => x"38",
          5228 => x"80",
          5229 => x"81",
          5230 => x"52",
          5231 => x"51",
          5232 => x"82",
          5233 => x"81",
          5234 => x"81",
          5235 => x"83",
          5236 => x"86",
          5237 => x"2e",
          5238 => x"82",
          5239 => x"06",
          5240 => x"56",
          5241 => x"38",
          5242 => x"74",
          5243 => x"a3",
          5244 => x"cc",
          5245 => x"06",
          5246 => x"2e",
          5247 => x"80",
          5248 => x"3d",
          5249 => x"83",
          5250 => x"15",
          5251 => x"53",
          5252 => x"8d",
          5253 => x"15",
          5254 => x"3f",
          5255 => x"08",
          5256 => x"70",
          5257 => x"0c",
          5258 => x"16",
          5259 => x"80",
          5260 => x"80",
          5261 => x"54",
          5262 => x"84",
          5263 => x"5b",
          5264 => x"80",
          5265 => x"7a",
          5266 => x"fc",
          5267 => x"87",
          5268 => x"ff",
          5269 => x"77",
          5270 => x"81",
          5271 => x"76",
          5272 => x"81",
          5273 => x"2e",
          5274 => x"8d",
          5275 => x"26",
          5276 => x"bf",
          5277 => x"f4",
          5278 => x"cc",
          5279 => x"ff",
          5280 => x"84",
          5281 => x"81",
          5282 => x"38",
          5283 => x"51",
          5284 => x"82",
          5285 => x"83",
          5286 => x"58",
          5287 => x"80",
          5288 => x"db",
          5289 => x"87",
          5290 => x"77",
          5291 => x"80",
          5292 => x"82",
          5293 => x"c4",
          5294 => x"11",
          5295 => x"06",
          5296 => x"8d",
          5297 => x"26",
          5298 => x"74",
          5299 => x"78",
          5300 => x"c1",
          5301 => x"59",
          5302 => x"15",
          5303 => x"2e",
          5304 => x"13",
          5305 => x"72",
          5306 => x"38",
          5307 => x"ea",
          5308 => x"14",
          5309 => x"3f",
          5310 => x"08",
          5311 => x"cc",
          5312 => x"23",
          5313 => x"57",
          5314 => x"83",
          5315 => x"c7",
          5316 => x"d8",
          5317 => x"cc",
          5318 => x"ff",
          5319 => x"8d",
          5320 => x"14",
          5321 => x"3f",
          5322 => x"08",
          5323 => x"14",
          5324 => x"3f",
          5325 => x"08",
          5326 => x"06",
          5327 => x"72",
          5328 => x"96",
          5329 => x"22",
          5330 => x"84",
          5331 => x"5a",
          5332 => x"83",
          5333 => x"14",
          5334 => x"79",
          5335 => x"8c",
          5336 => x"cc",
          5337 => x"87",
          5338 => x"2e",
          5339 => x"82",
          5340 => x"80",
          5341 => x"f5",
          5342 => x"83",
          5343 => x"ff",
          5344 => x"38",
          5345 => x"9f",
          5346 => x"38",
          5347 => x"39",
          5348 => x"80",
          5349 => x"38",
          5350 => x"98",
          5351 => x"a0",
          5352 => x"1c",
          5353 => x"0c",
          5354 => x"17",
          5355 => x"76",
          5356 => x"81",
          5357 => x"80",
          5358 => x"d9",
          5359 => x"87",
          5360 => x"ff",
          5361 => x"8d",
          5362 => x"8e",
          5363 => x"8a",
          5364 => x"14",
          5365 => x"3f",
          5366 => x"08",
          5367 => x"74",
          5368 => x"a2",
          5369 => x"79",
          5370 => x"ee",
          5371 => x"a8",
          5372 => x"15",
          5373 => x"2e",
          5374 => x"10",
          5375 => x"2a",
          5376 => x"05",
          5377 => x"ff",
          5378 => x"53",
          5379 => x"9c",
          5380 => x"81",
          5381 => x"0b",
          5382 => x"ff",
          5383 => x"0c",
          5384 => x"84",
          5385 => x"83",
          5386 => x"06",
          5387 => x"80",
          5388 => x"d8",
          5389 => x"87",
          5390 => x"ff",
          5391 => x"72",
          5392 => x"81",
          5393 => x"38",
          5394 => x"73",
          5395 => x"3f",
          5396 => x"08",
          5397 => x"82",
          5398 => x"84",
          5399 => x"b2",
          5400 => x"88",
          5401 => x"cc",
          5402 => x"ff",
          5403 => x"82",
          5404 => x"09",
          5405 => x"c8",
          5406 => x"51",
          5407 => x"82",
          5408 => x"84",
          5409 => x"d2",
          5410 => x"06",
          5411 => x"98",
          5412 => x"ef",
          5413 => x"cc",
          5414 => x"85",
          5415 => x"09",
          5416 => x"38",
          5417 => x"51",
          5418 => x"82",
          5419 => x"90",
          5420 => x"a0",
          5421 => x"cb",
          5422 => x"cc",
          5423 => x"0c",
          5424 => x"82",
          5425 => x"81",
          5426 => x"82",
          5427 => x"72",
          5428 => x"80",
          5429 => x"0c",
          5430 => x"82",
          5431 => x"90",
          5432 => x"fb",
          5433 => x"54",
          5434 => x"80",
          5435 => x"73",
          5436 => x"80",
          5437 => x"72",
          5438 => x"80",
          5439 => x"86",
          5440 => x"15",
          5441 => x"71",
          5442 => x"81",
          5443 => x"81",
          5444 => x"d0",
          5445 => x"87",
          5446 => x"06",
          5447 => x"38",
          5448 => x"54",
          5449 => x"80",
          5450 => x"71",
          5451 => x"82",
          5452 => x"87",
          5453 => x"fa",
          5454 => x"ab",
          5455 => x"58",
          5456 => x"05",
          5457 => x"e7",
          5458 => x"80",
          5459 => x"cc",
          5460 => x"38",
          5461 => x"08",
          5462 => x"9e",
          5463 => x"08",
          5464 => x"80",
          5465 => x"80",
          5466 => x"54",
          5467 => x"84",
          5468 => x"34",
          5469 => x"75",
          5470 => x"2e",
          5471 => x"53",
          5472 => x"53",
          5473 => x"f7",
          5474 => x"87",
          5475 => x"73",
          5476 => x"0c",
          5477 => x"04",
          5478 => x"67",
          5479 => x"80",
          5480 => x"59",
          5481 => x"78",
          5482 => x"c8",
          5483 => x"06",
          5484 => x"3d",
          5485 => x"99",
          5486 => x"52",
          5487 => x"3f",
          5488 => x"08",
          5489 => x"cc",
          5490 => x"38",
          5491 => x"52",
          5492 => x"52",
          5493 => x"3f",
          5494 => x"08",
          5495 => x"cc",
          5496 => x"02",
          5497 => x"33",
          5498 => x"55",
          5499 => x"25",
          5500 => x"55",
          5501 => x"54",
          5502 => x"81",
          5503 => x"80",
          5504 => x"74",
          5505 => x"81",
          5506 => x"75",
          5507 => x"3f",
          5508 => x"08",
          5509 => x"02",
          5510 => x"91",
          5511 => x"81",
          5512 => x"82",
          5513 => x"06",
          5514 => x"80",
          5515 => x"88",
          5516 => x"39",
          5517 => x"58",
          5518 => x"38",
          5519 => x"70",
          5520 => x"54",
          5521 => x"81",
          5522 => x"52",
          5523 => x"a6",
          5524 => x"cc",
          5525 => x"88",
          5526 => x"62",
          5527 => x"d4",
          5528 => x"54",
          5529 => x"15",
          5530 => x"62",
          5531 => x"e8",
          5532 => x"52",
          5533 => x"51",
          5534 => x"7a",
          5535 => x"83",
          5536 => x"80",
          5537 => x"38",
          5538 => x"08",
          5539 => x"53",
          5540 => x"3d",
          5541 => x"dd",
          5542 => x"87",
          5543 => x"82",
          5544 => x"82",
          5545 => x"39",
          5546 => x"38",
          5547 => x"33",
          5548 => x"70",
          5549 => x"55",
          5550 => x"2e",
          5551 => x"55",
          5552 => x"77",
          5553 => x"81",
          5554 => x"73",
          5555 => x"38",
          5556 => x"54",
          5557 => x"a0",
          5558 => x"82",
          5559 => x"52",
          5560 => x"a4",
          5561 => x"cc",
          5562 => x"18",
          5563 => x"55",
          5564 => x"cc",
          5565 => x"38",
          5566 => x"70",
          5567 => x"54",
          5568 => x"86",
          5569 => x"c0",
          5570 => x"b0",
          5571 => x"1b",
          5572 => x"1b",
          5573 => x"70",
          5574 => x"da",
          5575 => x"cc",
          5576 => x"cc",
          5577 => x"0c",
          5578 => x"52",
          5579 => x"3f",
          5580 => x"08",
          5581 => x"08",
          5582 => x"77",
          5583 => x"86",
          5584 => x"1a",
          5585 => x"1a",
          5586 => x"91",
          5587 => x"0b",
          5588 => x"80",
          5589 => x"0c",
          5590 => x"70",
          5591 => x"54",
          5592 => x"81",
          5593 => x"87",
          5594 => x"2e",
          5595 => x"82",
          5596 => x"94",
          5597 => x"17",
          5598 => x"2b",
          5599 => x"57",
          5600 => x"52",
          5601 => x"a0",
          5602 => x"cc",
          5603 => x"87",
          5604 => x"26",
          5605 => x"55",
          5606 => x"08",
          5607 => x"81",
          5608 => x"79",
          5609 => x"31",
          5610 => x"70",
          5611 => x"25",
          5612 => x"76",
          5613 => x"81",
          5614 => x"55",
          5615 => x"38",
          5616 => x"0c",
          5617 => x"75",
          5618 => x"54",
          5619 => x"a2",
          5620 => x"7a",
          5621 => x"3f",
          5622 => x"08",
          5623 => x"55",
          5624 => x"89",
          5625 => x"cc",
          5626 => x"1a",
          5627 => x"80",
          5628 => x"54",
          5629 => x"cc",
          5630 => x"0d",
          5631 => x"0d",
          5632 => x"64",
          5633 => x"59",
          5634 => x"90",
          5635 => x"52",
          5636 => x"cf",
          5637 => x"cc",
          5638 => x"87",
          5639 => x"38",
          5640 => x"55",
          5641 => x"86",
          5642 => x"82",
          5643 => x"19",
          5644 => x"55",
          5645 => x"80",
          5646 => x"38",
          5647 => x"0b",
          5648 => x"82",
          5649 => x"39",
          5650 => x"1a",
          5651 => x"82",
          5652 => x"19",
          5653 => x"08",
          5654 => x"7c",
          5655 => x"74",
          5656 => x"2e",
          5657 => x"94",
          5658 => x"83",
          5659 => x"56",
          5660 => x"38",
          5661 => x"22",
          5662 => x"89",
          5663 => x"55",
          5664 => x"75",
          5665 => x"19",
          5666 => x"39",
          5667 => x"52",
          5668 => x"94",
          5669 => x"cc",
          5670 => x"75",
          5671 => x"38",
          5672 => x"ff",
          5673 => x"98",
          5674 => x"19",
          5675 => x"51",
          5676 => x"82",
          5677 => x"80",
          5678 => x"38",
          5679 => x"08",
          5680 => x"2a",
          5681 => x"80",
          5682 => x"38",
          5683 => x"8a",
          5684 => x"5c",
          5685 => x"27",
          5686 => x"7a",
          5687 => x"54",
          5688 => x"52",
          5689 => x"51",
          5690 => x"82",
          5691 => x"fe",
          5692 => x"83",
          5693 => x"56",
          5694 => x"9f",
          5695 => x"08",
          5696 => x"74",
          5697 => x"38",
          5698 => x"b4",
          5699 => x"16",
          5700 => x"89",
          5701 => x"51",
          5702 => x"77",
          5703 => x"b9",
          5704 => x"1a",
          5705 => x"08",
          5706 => x"84",
          5707 => x"57",
          5708 => x"27",
          5709 => x"56",
          5710 => x"52",
          5711 => x"c8",
          5712 => x"cc",
          5713 => x"38",
          5714 => x"19",
          5715 => x"06",
          5716 => x"52",
          5717 => x"a3",
          5718 => x"31",
          5719 => x"7f",
          5720 => x"94",
          5721 => x"94",
          5722 => x"5c",
          5723 => x"80",
          5724 => x"87",
          5725 => x"3d",
          5726 => x"3d",
          5727 => x"65",
          5728 => x"5d",
          5729 => x"0c",
          5730 => x"05",
          5731 => x"f6",
          5732 => x"87",
          5733 => x"82",
          5734 => x"8a",
          5735 => x"33",
          5736 => x"2e",
          5737 => x"56",
          5738 => x"90",
          5739 => x"81",
          5740 => x"06",
          5741 => x"87",
          5742 => x"2e",
          5743 => x"95",
          5744 => x"91",
          5745 => x"56",
          5746 => x"81",
          5747 => x"34",
          5748 => x"8e",
          5749 => x"08",
          5750 => x"56",
          5751 => x"84",
          5752 => x"5c",
          5753 => x"82",
          5754 => x"18",
          5755 => x"ff",
          5756 => x"74",
          5757 => x"7e",
          5758 => x"ff",
          5759 => x"2a",
          5760 => x"7a",
          5761 => x"8c",
          5762 => x"08",
          5763 => x"38",
          5764 => x"39",
          5765 => x"52",
          5766 => x"e8",
          5767 => x"cc",
          5768 => x"87",
          5769 => x"2e",
          5770 => x"74",
          5771 => x"91",
          5772 => x"2e",
          5773 => x"74",
          5774 => x"88",
          5775 => x"38",
          5776 => x"0c",
          5777 => x"15",
          5778 => x"08",
          5779 => x"06",
          5780 => x"51",
          5781 => x"82",
          5782 => x"fe",
          5783 => x"18",
          5784 => x"51",
          5785 => x"82",
          5786 => x"80",
          5787 => x"38",
          5788 => x"08",
          5789 => x"2a",
          5790 => x"80",
          5791 => x"38",
          5792 => x"8a",
          5793 => x"5b",
          5794 => x"27",
          5795 => x"7b",
          5796 => x"54",
          5797 => x"52",
          5798 => x"51",
          5799 => x"82",
          5800 => x"fe",
          5801 => x"b0",
          5802 => x"31",
          5803 => x"79",
          5804 => x"84",
          5805 => x"16",
          5806 => x"89",
          5807 => x"52",
          5808 => x"cc",
          5809 => x"55",
          5810 => x"16",
          5811 => x"2b",
          5812 => x"39",
          5813 => x"94",
          5814 => x"93",
          5815 => x"cd",
          5816 => x"87",
          5817 => x"e3",
          5818 => x"b0",
          5819 => x"76",
          5820 => x"94",
          5821 => x"ff",
          5822 => x"71",
          5823 => x"7b",
          5824 => x"38",
          5825 => x"18",
          5826 => x"51",
          5827 => x"82",
          5828 => x"fd",
          5829 => x"53",
          5830 => x"18",
          5831 => x"06",
          5832 => x"51",
          5833 => x"7e",
          5834 => x"83",
          5835 => x"76",
          5836 => x"17",
          5837 => x"1e",
          5838 => x"18",
          5839 => x"0c",
          5840 => x"58",
          5841 => x"74",
          5842 => x"38",
          5843 => x"8c",
          5844 => x"90",
          5845 => x"33",
          5846 => x"55",
          5847 => x"34",
          5848 => x"82",
          5849 => x"90",
          5850 => x"f8",
          5851 => x"8b",
          5852 => x"53",
          5853 => x"f2",
          5854 => x"87",
          5855 => x"82",
          5856 => x"80",
          5857 => x"16",
          5858 => x"2a",
          5859 => x"51",
          5860 => x"80",
          5861 => x"38",
          5862 => x"52",
          5863 => x"e8",
          5864 => x"cc",
          5865 => x"87",
          5866 => x"d4",
          5867 => x"08",
          5868 => x"a0",
          5869 => x"73",
          5870 => x"88",
          5871 => x"74",
          5872 => x"51",
          5873 => x"8c",
          5874 => x"9c",
          5875 => x"fc",
          5876 => x"b2",
          5877 => x"15",
          5878 => x"3f",
          5879 => x"15",
          5880 => x"3f",
          5881 => x"0b",
          5882 => x"78",
          5883 => x"3f",
          5884 => x"08",
          5885 => x"81",
          5886 => x"57",
          5887 => x"34",
          5888 => x"cc",
          5889 => x"0d",
          5890 => x"0d",
          5891 => x"54",
          5892 => x"82",
          5893 => x"53",
          5894 => x"08",
          5895 => x"3d",
          5896 => x"73",
          5897 => x"3f",
          5898 => x"08",
          5899 => x"cc",
          5900 => x"82",
          5901 => x"74",
          5902 => x"87",
          5903 => x"3d",
          5904 => x"3d",
          5905 => x"51",
          5906 => x"8b",
          5907 => x"82",
          5908 => x"24",
          5909 => x"87",
          5910 => x"9f",
          5911 => x"52",
          5912 => x"cc",
          5913 => x"0d",
          5914 => x"0d",
          5915 => x"3d",
          5916 => x"94",
          5917 => x"c2",
          5918 => x"cc",
          5919 => x"87",
          5920 => x"e0",
          5921 => x"63",
          5922 => x"d4",
          5923 => x"8e",
          5924 => x"cc",
          5925 => x"87",
          5926 => x"38",
          5927 => x"05",
          5928 => x"2b",
          5929 => x"80",
          5930 => x"76",
          5931 => x"0c",
          5932 => x"02",
          5933 => x"70",
          5934 => x"81",
          5935 => x"56",
          5936 => x"9e",
          5937 => x"53",
          5938 => x"db",
          5939 => x"87",
          5940 => x"15",
          5941 => x"82",
          5942 => x"84",
          5943 => x"06",
          5944 => x"55",
          5945 => x"cc",
          5946 => x"0d",
          5947 => x"0d",
          5948 => x"5b",
          5949 => x"80",
          5950 => x"ff",
          5951 => x"9f",
          5952 => x"b6",
          5953 => x"cc",
          5954 => x"87",
          5955 => x"fc",
          5956 => x"7a",
          5957 => x"08",
          5958 => x"64",
          5959 => x"2e",
          5960 => x"a0",
          5961 => x"70",
          5962 => x"eb",
          5963 => x"cc",
          5964 => x"87",
          5965 => x"d4",
          5966 => x"7b",
          5967 => x"3f",
          5968 => x"08",
          5969 => x"cc",
          5970 => x"38",
          5971 => x"51",
          5972 => x"82",
          5973 => x"45",
          5974 => x"51",
          5975 => x"82",
          5976 => x"57",
          5977 => x"08",
          5978 => x"80",
          5979 => x"da",
          5980 => x"87",
          5981 => x"82",
          5982 => x"a4",
          5983 => x"7b",
          5984 => x"3f",
          5985 => x"cc",
          5986 => x"38",
          5987 => x"51",
          5988 => x"82",
          5989 => x"57",
          5990 => x"08",
          5991 => x"38",
          5992 => x"09",
          5993 => x"38",
          5994 => x"e0",
          5995 => x"dc",
          5996 => x"ff",
          5997 => x"74",
          5998 => x"3f",
          5999 => x"78",
          6000 => x"33",
          6001 => x"56",
          6002 => x"91",
          6003 => x"05",
          6004 => x"81",
          6005 => x"56",
          6006 => x"f5",
          6007 => x"54",
          6008 => x"81",
          6009 => x"80",
          6010 => x"78",
          6011 => x"55",
          6012 => x"11",
          6013 => x"18",
          6014 => x"58",
          6015 => x"34",
          6016 => x"ff",
          6017 => x"55",
          6018 => x"34",
          6019 => x"77",
          6020 => x"81",
          6021 => x"ff",
          6022 => x"55",
          6023 => x"34",
          6024 => x"9f",
          6025 => x"84",
          6026 => x"84",
          6027 => x"70",
          6028 => x"56",
          6029 => x"76",
          6030 => x"81",
          6031 => x"70",
          6032 => x"56",
          6033 => x"82",
          6034 => x"78",
          6035 => x"80",
          6036 => x"27",
          6037 => x"19",
          6038 => x"7a",
          6039 => x"5c",
          6040 => x"55",
          6041 => x"7a",
          6042 => x"5c",
          6043 => x"2e",
          6044 => x"85",
          6045 => x"94",
          6046 => x"81",
          6047 => x"73",
          6048 => x"81",
          6049 => x"7a",
          6050 => x"38",
          6051 => x"76",
          6052 => x"0c",
          6053 => x"04",
          6054 => x"7b",
          6055 => x"fc",
          6056 => x"53",
          6057 => x"bb",
          6058 => x"cc",
          6059 => x"87",
          6060 => x"fa",
          6061 => x"33",
          6062 => x"f2",
          6063 => x"08",
          6064 => x"27",
          6065 => x"15",
          6066 => x"2a",
          6067 => x"51",
          6068 => x"83",
          6069 => x"94",
          6070 => x"80",
          6071 => x"0c",
          6072 => x"2e",
          6073 => x"79",
          6074 => x"70",
          6075 => x"51",
          6076 => x"2e",
          6077 => x"52",
          6078 => x"ff",
          6079 => x"82",
          6080 => x"ff",
          6081 => x"70",
          6082 => x"ff",
          6083 => x"82",
          6084 => x"73",
          6085 => x"76",
          6086 => x"06",
          6087 => x"0c",
          6088 => x"98",
          6089 => x"58",
          6090 => x"39",
          6091 => x"54",
          6092 => x"73",
          6093 => x"cd",
          6094 => x"87",
          6095 => x"82",
          6096 => x"81",
          6097 => x"38",
          6098 => x"08",
          6099 => x"9b",
          6100 => x"cc",
          6101 => x"0c",
          6102 => x"0c",
          6103 => x"81",
          6104 => x"76",
          6105 => x"38",
          6106 => x"94",
          6107 => x"94",
          6108 => x"16",
          6109 => x"2a",
          6110 => x"51",
          6111 => x"72",
          6112 => x"38",
          6113 => x"51",
          6114 => x"82",
          6115 => x"54",
          6116 => x"08",
          6117 => x"87",
          6118 => x"a7",
          6119 => x"74",
          6120 => x"3f",
          6121 => x"08",
          6122 => x"2e",
          6123 => x"74",
          6124 => x"79",
          6125 => x"14",
          6126 => x"38",
          6127 => x"0c",
          6128 => x"94",
          6129 => x"94",
          6130 => x"83",
          6131 => x"72",
          6132 => x"38",
          6133 => x"51",
          6134 => x"82",
          6135 => x"94",
          6136 => x"91",
          6137 => x"53",
          6138 => x"81",
          6139 => x"34",
          6140 => x"39",
          6141 => x"82",
          6142 => x"05",
          6143 => x"08",
          6144 => x"08",
          6145 => x"38",
          6146 => x"0c",
          6147 => x"80",
          6148 => x"72",
          6149 => x"73",
          6150 => x"53",
          6151 => x"8c",
          6152 => x"16",
          6153 => x"38",
          6154 => x"0c",
          6155 => x"82",
          6156 => x"8b",
          6157 => x"f9",
          6158 => x"56",
          6159 => x"80",
          6160 => x"38",
          6161 => x"3d",
          6162 => x"8a",
          6163 => x"51",
          6164 => x"82",
          6165 => x"55",
          6166 => x"08",
          6167 => x"77",
          6168 => x"52",
          6169 => x"b6",
          6170 => x"cc",
          6171 => x"87",
          6172 => x"c3",
          6173 => x"33",
          6174 => x"55",
          6175 => x"24",
          6176 => x"16",
          6177 => x"2a",
          6178 => x"51",
          6179 => x"80",
          6180 => x"9c",
          6181 => x"77",
          6182 => x"3f",
          6183 => x"08",
          6184 => x"77",
          6185 => x"22",
          6186 => x"74",
          6187 => x"ce",
          6188 => x"87",
          6189 => x"74",
          6190 => x"81",
          6191 => x"85",
          6192 => x"74",
          6193 => x"38",
          6194 => x"74",
          6195 => x"87",
          6196 => x"3d",
          6197 => x"3d",
          6198 => x"3d",
          6199 => x"70",
          6200 => x"ff",
          6201 => x"cc",
          6202 => x"82",
          6203 => x"73",
          6204 => x"0d",
          6205 => x"0d",
          6206 => x"3d",
          6207 => x"71",
          6208 => x"e7",
          6209 => x"87",
          6210 => x"82",
          6211 => x"80",
          6212 => x"93",
          6213 => x"cc",
          6214 => x"51",
          6215 => x"82",
          6216 => x"53",
          6217 => x"82",
          6218 => x"52",
          6219 => x"ad",
          6220 => x"cc",
          6221 => x"87",
          6222 => x"2e",
          6223 => x"85",
          6224 => x"87",
          6225 => x"cc",
          6226 => x"74",
          6227 => x"d5",
          6228 => x"52",
          6229 => x"8a",
          6230 => x"cc",
          6231 => x"70",
          6232 => x"07",
          6233 => x"82",
          6234 => x"06",
          6235 => x"54",
          6236 => x"cc",
          6237 => x"0d",
          6238 => x"0d",
          6239 => x"53",
          6240 => x"53",
          6241 => x"56",
          6242 => x"82",
          6243 => x"55",
          6244 => x"08",
          6245 => x"52",
          6246 => x"82",
          6247 => x"cc",
          6248 => x"87",
          6249 => x"38",
          6250 => x"05",
          6251 => x"2b",
          6252 => x"80",
          6253 => x"86",
          6254 => x"76",
          6255 => x"38",
          6256 => x"51",
          6257 => x"74",
          6258 => x"0c",
          6259 => x"04",
          6260 => x"63",
          6261 => x"80",
          6262 => x"ec",
          6263 => x"3d",
          6264 => x"3f",
          6265 => x"08",
          6266 => x"cc",
          6267 => x"38",
          6268 => x"73",
          6269 => x"08",
          6270 => x"13",
          6271 => x"58",
          6272 => x"26",
          6273 => x"7c",
          6274 => x"39",
          6275 => x"cc",
          6276 => x"81",
          6277 => x"87",
          6278 => x"33",
          6279 => x"81",
          6280 => x"06",
          6281 => x"75",
          6282 => x"52",
          6283 => x"05",
          6284 => x"3f",
          6285 => x"08",
          6286 => x"38",
          6287 => x"08",
          6288 => x"38",
          6289 => x"08",
          6290 => x"87",
          6291 => x"80",
          6292 => x"81",
          6293 => x"59",
          6294 => x"14",
          6295 => x"ca",
          6296 => x"39",
          6297 => x"82",
          6298 => x"57",
          6299 => x"38",
          6300 => x"18",
          6301 => x"ff",
          6302 => x"82",
          6303 => x"5b",
          6304 => x"08",
          6305 => x"7c",
          6306 => x"12",
          6307 => x"52",
          6308 => x"82",
          6309 => x"06",
          6310 => x"14",
          6311 => x"cc",
          6312 => x"cc",
          6313 => x"ff",
          6314 => x"70",
          6315 => x"82",
          6316 => x"51",
          6317 => x"b4",
          6318 => x"bb",
          6319 => x"87",
          6320 => x"0a",
          6321 => x"70",
          6322 => x"84",
          6323 => x"51",
          6324 => x"ff",
          6325 => x"56",
          6326 => x"38",
          6327 => x"7c",
          6328 => x"0c",
          6329 => x"81",
          6330 => x"74",
          6331 => x"7a",
          6332 => x"0c",
          6333 => x"04",
          6334 => x"79",
          6335 => x"05",
          6336 => x"57",
          6337 => x"82",
          6338 => x"56",
          6339 => x"08",
          6340 => x"91",
          6341 => x"75",
          6342 => x"90",
          6343 => x"81",
          6344 => x"06",
          6345 => x"87",
          6346 => x"2e",
          6347 => x"94",
          6348 => x"73",
          6349 => x"27",
          6350 => x"73",
          6351 => x"87",
          6352 => x"88",
          6353 => x"76",
          6354 => x"3f",
          6355 => x"08",
          6356 => x"0c",
          6357 => x"39",
          6358 => x"52",
          6359 => x"bf",
          6360 => x"87",
          6361 => x"2e",
          6362 => x"83",
          6363 => x"82",
          6364 => x"81",
          6365 => x"06",
          6366 => x"56",
          6367 => x"a0",
          6368 => x"82",
          6369 => x"98",
          6370 => x"94",
          6371 => x"08",
          6372 => x"cc",
          6373 => x"51",
          6374 => x"82",
          6375 => x"56",
          6376 => x"8c",
          6377 => x"17",
          6378 => x"07",
          6379 => x"18",
          6380 => x"2e",
          6381 => x"91",
          6382 => x"55",
          6383 => x"cc",
          6384 => x"0d",
          6385 => x"0d",
          6386 => x"3d",
          6387 => x"52",
          6388 => x"da",
          6389 => x"87",
          6390 => x"82",
          6391 => x"81",
          6392 => x"45",
          6393 => x"52",
          6394 => x"52",
          6395 => x"3f",
          6396 => x"08",
          6397 => x"cc",
          6398 => x"38",
          6399 => x"05",
          6400 => x"2a",
          6401 => x"51",
          6402 => x"55",
          6403 => x"38",
          6404 => x"54",
          6405 => x"81",
          6406 => x"80",
          6407 => x"70",
          6408 => x"54",
          6409 => x"81",
          6410 => x"52",
          6411 => x"c6",
          6412 => x"cc",
          6413 => x"2a",
          6414 => x"51",
          6415 => x"80",
          6416 => x"38",
          6417 => x"87",
          6418 => x"15",
          6419 => x"86",
          6420 => x"82",
          6421 => x"5c",
          6422 => x"3d",
          6423 => x"c7",
          6424 => x"87",
          6425 => x"82",
          6426 => x"80",
          6427 => x"87",
          6428 => x"73",
          6429 => x"3f",
          6430 => x"08",
          6431 => x"cc",
          6432 => x"87",
          6433 => x"39",
          6434 => x"08",
          6435 => x"38",
          6436 => x"08",
          6437 => x"77",
          6438 => x"3f",
          6439 => x"08",
          6440 => x"08",
          6441 => x"87",
          6442 => x"80",
          6443 => x"55",
          6444 => x"94",
          6445 => x"2e",
          6446 => x"53",
          6447 => x"51",
          6448 => x"82",
          6449 => x"55",
          6450 => x"78",
          6451 => x"ff",
          6452 => x"cc",
          6453 => x"82",
          6454 => x"a0",
          6455 => x"e9",
          6456 => x"53",
          6457 => x"05",
          6458 => x"51",
          6459 => x"82",
          6460 => x"54",
          6461 => x"08",
          6462 => x"78",
          6463 => x"8e",
          6464 => x"58",
          6465 => x"82",
          6466 => x"54",
          6467 => x"08",
          6468 => x"54",
          6469 => x"82",
          6470 => x"84",
          6471 => x"06",
          6472 => x"02",
          6473 => x"33",
          6474 => x"81",
          6475 => x"86",
          6476 => x"f6",
          6477 => x"74",
          6478 => x"70",
          6479 => x"c4",
          6480 => x"cc",
          6481 => x"56",
          6482 => x"08",
          6483 => x"54",
          6484 => x"08",
          6485 => x"81",
          6486 => x"82",
          6487 => x"cc",
          6488 => x"09",
          6489 => x"38",
          6490 => x"b4",
          6491 => x"b0",
          6492 => x"cc",
          6493 => x"51",
          6494 => x"82",
          6495 => x"54",
          6496 => x"08",
          6497 => x"8b",
          6498 => x"b4",
          6499 => x"b7",
          6500 => x"54",
          6501 => x"15",
          6502 => x"90",
          6503 => x"34",
          6504 => x"0a",
          6505 => x"19",
          6506 => x"a0",
          6507 => x"78",
          6508 => x"51",
          6509 => x"a0",
          6510 => x"11",
          6511 => x"05",
          6512 => x"b7",
          6513 => x"ae",
          6514 => x"15",
          6515 => x"78",
          6516 => x"53",
          6517 => x"3f",
          6518 => x"0b",
          6519 => x"77",
          6520 => x"3f",
          6521 => x"08",
          6522 => x"cc",
          6523 => x"82",
          6524 => x"52",
          6525 => x"51",
          6526 => x"3f",
          6527 => x"52",
          6528 => x"ab",
          6529 => x"90",
          6530 => x"34",
          6531 => x"0b",
          6532 => x"78",
          6533 => x"b7",
          6534 => x"cc",
          6535 => x"39",
          6536 => x"52",
          6537 => x"be",
          6538 => x"82",
          6539 => x"99",
          6540 => x"da",
          6541 => x"3d",
          6542 => x"d2",
          6543 => x"53",
          6544 => x"84",
          6545 => x"3d",
          6546 => x"3f",
          6547 => x"08",
          6548 => x"cc",
          6549 => x"38",
          6550 => x"3d",
          6551 => x"3d",
          6552 => x"cc",
          6553 => x"87",
          6554 => x"82",
          6555 => x"82",
          6556 => x"81",
          6557 => x"81",
          6558 => x"86",
          6559 => x"aa",
          6560 => x"a4",
          6561 => x"a8",
          6562 => x"05",
          6563 => x"eb",
          6564 => x"77",
          6565 => x"70",
          6566 => x"b4",
          6567 => x"3d",
          6568 => x"51",
          6569 => x"82",
          6570 => x"55",
          6571 => x"08",
          6572 => x"6f",
          6573 => x"06",
          6574 => x"a2",
          6575 => x"92",
          6576 => x"81",
          6577 => x"87",
          6578 => x"2e",
          6579 => x"81",
          6580 => x"51",
          6581 => x"82",
          6582 => x"55",
          6583 => x"08",
          6584 => x"68",
          6585 => x"a8",
          6586 => x"05",
          6587 => x"51",
          6588 => x"3f",
          6589 => x"33",
          6590 => x"8b",
          6591 => x"84",
          6592 => x"06",
          6593 => x"73",
          6594 => x"a0",
          6595 => x"8b",
          6596 => x"54",
          6597 => x"15",
          6598 => x"33",
          6599 => x"70",
          6600 => x"55",
          6601 => x"2e",
          6602 => x"6e",
          6603 => x"df",
          6604 => x"78",
          6605 => x"3f",
          6606 => x"08",
          6607 => x"ff",
          6608 => x"82",
          6609 => x"cc",
          6610 => x"80",
          6611 => x"87",
          6612 => x"78",
          6613 => x"b0",
          6614 => x"cc",
          6615 => x"d4",
          6616 => x"55",
          6617 => x"08",
          6618 => x"81",
          6619 => x"73",
          6620 => x"81",
          6621 => x"63",
          6622 => x"76",
          6623 => x"3f",
          6624 => x"0b",
          6625 => x"87",
          6626 => x"cc",
          6627 => x"77",
          6628 => x"3f",
          6629 => x"08",
          6630 => x"cc",
          6631 => x"78",
          6632 => x"ab",
          6633 => x"cc",
          6634 => x"82",
          6635 => x"a8",
          6636 => x"ed",
          6637 => x"80",
          6638 => x"02",
          6639 => x"df",
          6640 => x"57",
          6641 => x"3d",
          6642 => x"96",
          6643 => x"ea",
          6644 => x"cc",
          6645 => x"87",
          6646 => x"cf",
          6647 => x"65",
          6648 => x"d4",
          6649 => x"b6",
          6650 => x"cc",
          6651 => x"87",
          6652 => x"38",
          6653 => x"05",
          6654 => x"06",
          6655 => x"73",
          6656 => x"a7",
          6657 => x"09",
          6658 => x"71",
          6659 => x"06",
          6660 => x"55",
          6661 => x"15",
          6662 => x"81",
          6663 => x"34",
          6664 => x"b4",
          6665 => x"87",
          6666 => x"74",
          6667 => x"0c",
          6668 => x"04",
          6669 => x"64",
          6670 => x"93",
          6671 => x"52",
          6672 => x"d1",
          6673 => x"87",
          6674 => x"82",
          6675 => x"80",
          6676 => x"58",
          6677 => x"3d",
          6678 => x"c8",
          6679 => x"87",
          6680 => x"82",
          6681 => x"b4",
          6682 => x"c7",
          6683 => x"a0",
          6684 => x"55",
          6685 => x"84",
          6686 => x"17",
          6687 => x"2b",
          6688 => x"96",
          6689 => x"b0",
          6690 => x"54",
          6691 => x"15",
          6692 => x"ff",
          6693 => x"82",
          6694 => x"55",
          6695 => x"cc",
          6696 => x"0d",
          6697 => x"0d",
          6698 => x"5a",
          6699 => x"3d",
          6700 => x"99",
          6701 => x"82",
          6702 => x"cc",
          6703 => x"cc",
          6704 => x"82",
          6705 => x"07",
          6706 => x"55",
          6707 => x"2e",
          6708 => x"81",
          6709 => x"55",
          6710 => x"2e",
          6711 => x"7b",
          6712 => x"80",
          6713 => x"70",
          6714 => x"be",
          6715 => x"87",
          6716 => x"82",
          6717 => x"80",
          6718 => x"52",
          6719 => x"dd",
          6720 => x"cc",
          6721 => x"87",
          6722 => x"38",
          6723 => x"08",
          6724 => x"08",
          6725 => x"56",
          6726 => x"19",
          6727 => x"59",
          6728 => x"74",
          6729 => x"56",
          6730 => x"ec",
          6731 => x"75",
          6732 => x"74",
          6733 => x"2e",
          6734 => x"16",
          6735 => x"33",
          6736 => x"73",
          6737 => x"38",
          6738 => x"84",
          6739 => x"06",
          6740 => x"7a",
          6741 => x"76",
          6742 => x"07",
          6743 => x"54",
          6744 => x"80",
          6745 => x"80",
          6746 => x"7b",
          6747 => x"53",
          6748 => x"94",
          6749 => x"cc",
          6750 => x"87",
          6751 => x"38",
          6752 => x"55",
          6753 => x"56",
          6754 => x"8b",
          6755 => x"56",
          6756 => x"83",
          6757 => x"75",
          6758 => x"51",
          6759 => x"3f",
          6760 => x"08",
          6761 => x"82",
          6762 => x"98",
          6763 => x"e6",
          6764 => x"53",
          6765 => x"b8",
          6766 => x"3d",
          6767 => x"3f",
          6768 => x"08",
          6769 => x"08",
          6770 => x"87",
          6771 => x"98",
          6772 => x"a0",
          6773 => x"70",
          6774 => x"ae",
          6775 => x"6d",
          6776 => x"81",
          6777 => x"57",
          6778 => x"74",
          6779 => x"38",
          6780 => x"81",
          6781 => x"81",
          6782 => x"52",
          6783 => x"8a",
          6784 => x"cc",
          6785 => x"a5",
          6786 => x"33",
          6787 => x"54",
          6788 => x"3f",
          6789 => x"08",
          6790 => x"38",
          6791 => x"76",
          6792 => x"05",
          6793 => x"39",
          6794 => x"08",
          6795 => x"15",
          6796 => x"ff",
          6797 => x"73",
          6798 => x"38",
          6799 => x"83",
          6800 => x"56",
          6801 => x"75",
          6802 => x"82",
          6803 => x"33",
          6804 => x"2e",
          6805 => x"52",
          6806 => x"51",
          6807 => x"3f",
          6808 => x"08",
          6809 => x"ff",
          6810 => x"38",
          6811 => x"88",
          6812 => x"8a",
          6813 => x"38",
          6814 => x"ec",
          6815 => x"75",
          6816 => x"74",
          6817 => x"73",
          6818 => x"05",
          6819 => x"17",
          6820 => x"70",
          6821 => x"34",
          6822 => x"70",
          6823 => x"ff",
          6824 => x"55",
          6825 => x"26",
          6826 => x"8b",
          6827 => x"86",
          6828 => x"e5",
          6829 => x"38",
          6830 => x"99",
          6831 => x"05",
          6832 => x"70",
          6833 => x"73",
          6834 => x"81",
          6835 => x"ff",
          6836 => x"ed",
          6837 => x"80",
          6838 => x"91",
          6839 => x"55",
          6840 => x"3f",
          6841 => x"08",
          6842 => x"cc",
          6843 => x"38",
          6844 => x"51",
          6845 => x"3f",
          6846 => x"08",
          6847 => x"cc",
          6848 => x"76",
          6849 => x"67",
          6850 => x"34",
          6851 => x"82",
          6852 => x"84",
          6853 => x"06",
          6854 => x"80",
          6855 => x"2e",
          6856 => x"81",
          6857 => x"ff",
          6858 => x"82",
          6859 => x"54",
          6860 => x"08",
          6861 => x"53",
          6862 => x"08",
          6863 => x"ff",
          6864 => x"67",
          6865 => x"8b",
          6866 => x"53",
          6867 => x"51",
          6868 => x"3f",
          6869 => x"0b",
          6870 => x"79",
          6871 => x"ef",
          6872 => x"cc",
          6873 => x"55",
          6874 => x"cc",
          6875 => x"0d",
          6876 => x"0d",
          6877 => x"88",
          6878 => x"05",
          6879 => x"fc",
          6880 => x"54",
          6881 => x"d2",
          6882 => x"87",
          6883 => x"82",
          6884 => x"82",
          6885 => x"1a",
          6886 => x"82",
          6887 => x"80",
          6888 => x"8c",
          6889 => x"78",
          6890 => x"1a",
          6891 => x"2a",
          6892 => x"51",
          6893 => x"90",
          6894 => x"82",
          6895 => x"58",
          6896 => x"81",
          6897 => x"39",
          6898 => x"22",
          6899 => x"70",
          6900 => x"56",
          6901 => x"94",
          6902 => x"14",
          6903 => x"30",
          6904 => x"9f",
          6905 => x"cc",
          6906 => x"19",
          6907 => x"5a",
          6908 => x"81",
          6909 => x"38",
          6910 => x"77",
          6911 => x"82",
          6912 => x"56",
          6913 => x"74",
          6914 => x"ff",
          6915 => x"81",
          6916 => x"55",
          6917 => x"75",
          6918 => x"82",
          6919 => x"cc",
          6920 => x"ff",
          6921 => x"87",
          6922 => x"2e",
          6923 => x"82",
          6924 => x"8e",
          6925 => x"56",
          6926 => x"09",
          6927 => x"38",
          6928 => x"59",
          6929 => x"77",
          6930 => x"06",
          6931 => x"87",
          6932 => x"39",
          6933 => x"ba",
          6934 => x"55",
          6935 => x"2e",
          6936 => x"15",
          6937 => x"2e",
          6938 => x"83",
          6939 => x"75",
          6940 => x"7e",
          6941 => x"a9",
          6942 => x"cc",
          6943 => x"87",
          6944 => x"ce",
          6945 => x"16",
          6946 => x"56",
          6947 => x"38",
          6948 => x"19",
          6949 => x"8c",
          6950 => x"7d",
          6951 => x"38",
          6952 => x"0c",
          6953 => x"0c",
          6954 => x"80",
          6955 => x"73",
          6956 => x"98",
          6957 => x"05",
          6958 => x"57",
          6959 => x"26",
          6960 => x"7b",
          6961 => x"0c",
          6962 => x"81",
          6963 => x"84",
          6964 => x"54",
          6965 => x"cc",
          6966 => x"0d",
          6967 => x"0d",
          6968 => x"88",
          6969 => x"05",
          6970 => x"54",
          6971 => x"c5",
          6972 => x"56",
          6973 => x"87",
          6974 => x"8b",
          6975 => x"87",
          6976 => x"29",
          6977 => x"05",
          6978 => x"55",
          6979 => x"84",
          6980 => x"34",
          6981 => x"08",
          6982 => x"5f",
          6983 => x"51",
          6984 => x"3f",
          6985 => x"08",
          6986 => x"70",
          6987 => x"57",
          6988 => x"8b",
          6989 => x"82",
          6990 => x"06",
          6991 => x"56",
          6992 => x"38",
          6993 => x"05",
          6994 => x"7e",
          6995 => x"f1",
          6996 => x"cc",
          6997 => x"67",
          6998 => x"2e",
          6999 => x"82",
          7000 => x"8b",
          7001 => x"75",
          7002 => x"80",
          7003 => x"81",
          7004 => x"2e",
          7005 => x"80",
          7006 => x"38",
          7007 => x"0a",
          7008 => x"ff",
          7009 => x"55",
          7010 => x"86",
          7011 => x"8a",
          7012 => x"89",
          7013 => x"2a",
          7014 => x"77",
          7015 => x"59",
          7016 => x"81",
          7017 => x"70",
          7018 => x"07",
          7019 => x"56",
          7020 => x"38",
          7021 => x"05",
          7022 => x"7e",
          7023 => x"81",
          7024 => x"82",
          7025 => x"8a",
          7026 => x"83",
          7027 => x"06",
          7028 => x"08",
          7029 => x"74",
          7030 => x"41",
          7031 => x"56",
          7032 => x"8a",
          7033 => x"61",
          7034 => x"55",
          7035 => x"27",
          7036 => x"93",
          7037 => x"80",
          7038 => x"38",
          7039 => x"70",
          7040 => x"43",
          7041 => x"95",
          7042 => x"06",
          7043 => x"2e",
          7044 => x"77",
          7045 => x"74",
          7046 => x"83",
          7047 => x"06",
          7048 => x"82",
          7049 => x"2e",
          7050 => x"78",
          7051 => x"2e",
          7052 => x"80",
          7053 => x"ae",
          7054 => x"2a",
          7055 => x"82",
          7056 => x"56",
          7057 => x"2e",
          7058 => x"77",
          7059 => x"82",
          7060 => x"79",
          7061 => x"70",
          7062 => x"5a",
          7063 => x"86",
          7064 => x"27",
          7065 => x"52",
          7066 => x"8e",
          7067 => x"87",
          7068 => x"29",
          7069 => x"70",
          7070 => x"55",
          7071 => x"0b",
          7072 => x"08",
          7073 => x"05",
          7074 => x"ff",
          7075 => x"27",
          7076 => x"88",
          7077 => x"ae",
          7078 => x"2a",
          7079 => x"82",
          7080 => x"56",
          7081 => x"2e",
          7082 => x"77",
          7083 => x"82",
          7084 => x"79",
          7085 => x"70",
          7086 => x"5a",
          7087 => x"86",
          7088 => x"27",
          7089 => x"52",
          7090 => x"8e",
          7091 => x"87",
          7092 => x"84",
          7093 => x"87",
          7094 => x"f5",
          7095 => x"81",
          7096 => x"cc",
          7097 => x"87",
          7098 => x"71",
          7099 => x"83",
          7100 => x"5e",
          7101 => x"89",
          7102 => x"5c",
          7103 => x"1c",
          7104 => x"05",
          7105 => x"ff",
          7106 => x"70",
          7107 => x"31",
          7108 => x"57",
          7109 => x"83",
          7110 => x"06",
          7111 => x"1c",
          7112 => x"5c",
          7113 => x"1d",
          7114 => x"29",
          7115 => x"31",
          7116 => x"55",
          7117 => x"87",
          7118 => x"7c",
          7119 => x"7a",
          7120 => x"31",
          7121 => x"8d",
          7122 => x"87",
          7123 => x"7d",
          7124 => x"81",
          7125 => x"82",
          7126 => x"83",
          7127 => x"80",
          7128 => x"87",
          7129 => x"81",
          7130 => x"fd",
          7131 => x"f8",
          7132 => x"2e",
          7133 => x"80",
          7134 => x"ff",
          7135 => x"87",
          7136 => x"a0",
          7137 => x"38",
          7138 => x"74",
          7139 => x"86",
          7140 => x"fd",
          7141 => x"81",
          7142 => x"80",
          7143 => x"83",
          7144 => x"39",
          7145 => x"08",
          7146 => x"92",
          7147 => x"b8",
          7148 => x"59",
          7149 => x"27",
          7150 => x"86",
          7151 => x"55",
          7152 => x"09",
          7153 => x"38",
          7154 => x"f5",
          7155 => x"38",
          7156 => x"55",
          7157 => x"86",
          7158 => x"80",
          7159 => x"7a",
          7160 => x"ba",
          7161 => x"82",
          7162 => x"7a",
          7163 => x"8b",
          7164 => x"52",
          7165 => x"ff",
          7166 => x"79",
          7167 => x"7b",
          7168 => x"06",
          7169 => x"51",
          7170 => x"3f",
          7171 => x"1c",
          7172 => x"32",
          7173 => x"96",
          7174 => x"06",
          7175 => x"91",
          7176 => x"a1",
          7177 => x"55",
          7178 => x"ff",
          7179 => x"74",
          7180 => x"06",
          7181 => x"51",
          7182 => x"3f",
          7183 => x"52",
          7184 => x"ff",
          7185 => x"f8",
          7186 => x"34",
          7187 => x"1b",
          7188 => x"da",
          7189 => x"52",
          7190 => x"ff",
          7191 => x"60",
          7192 => x"51",
          7193 => x"3f",
          7194 => x"09",
          7195 => x"cb",
          7196 => x"b2",
          7197 => x"c3",
          7198 => x"a0",
          7199 => x"52",
          7200 => x"ff",
          7201 => x"82",
          7202 => x"51",
          7203 => x"3f",
          7204 => x"1b",
          7205 => x"96",
          7206 => x"b2",
          7207 => x"a0",
          7208 => x"80",
          7209 => x"1c",
          7210 => x"80",
          7211 => x"93",
          7212 => x"dc",
          7213 => x"1b",
          7214 => x"82",
          7215 => x"52",
          7216 => x"ff",
          7217 => x"7c",
          7218 => x"06",
          7219 => x"51",
          7220 => x"3f",
          7221 => x"a4",
          7222 => x"0b",
          7223 => x"93",
          7224 => x"f0",
          7225 => x"51",
          7226 => x"3f",
          7227 => x"52",
          7228 => x"70",
          7229 => x"9f",
          7230 => x"54",
          7231 => x"52",
          7232 => x"9b",
          7233 => x"56",
          7234 => x"08",
          7235 => x"7d",
          7236 => x"81",
          7237 => x"38",
          7238 => x"86",
          7239 => x"52",
          7240 => x"9b",
          7241 => x"80",
          7242 => x"7a",
          7243 => x"ee",
          7244 => x"85",
          7245 => x"7a",
          7246 => x"90",
          7247 => x"85",
          7248 => x"83",
          7249 => x"ff",
          7250 => x"ff",
          7251 => x"e8",
          7252 => x"9e",
          7253 => x"52",
          7254 => x"51",
          7255 => x"3f",
          7256 => x"52",
          7257 => x"9e",
          7258 => x"54",
          7259 => x"53",
          7260 => x"51",
          7261 => x"3f",
          7262 => x"16",
          7263 => x"7e",
          7264 => x"d9",
          7265 => x"80",
          7266 => x"ff",
          7267 => x"7f",
          7268 => x"7d",
          7269 => x"81",
          7270 => x"f8",
          7271 => x"ff",
          7272 => x"ff",
          7273 => x"51",
          7274 => x"3f",
          7275 => x"88",
          7276 => x"39",
          7277 => x"f8",
          7278 => x"2e",
          7279 => x"55",
          7280 => x"51",
          7281 => x"3f",
          7282 => x"57",
          7283 => x"83",
          7284 => x"76",
          7285 => x"7a",
          7286 => x"ff",
          7287 => x"82",
          7288 => x"82",
          7289 => x"80",
          7290 => x"cc",
          7291 => x"51",
          7292 => x"3f",
          7293 => x"78",
          7294 => x"74",
          7295 => x"18",
          7296 => x"2e",
          7297 => x"79",
          7298 => x"2e",
          7299 => x"55",
          7300 => x"62",
          7301 => x"74",
          7302 => x"75",
          7303 => x"7e",
          7304 => x"b9",
          7305 => x"cc",
          7306 => x"38",
          7307 => x"78",
          7308 => x"74",
          7309 => x"56",
          7310 => x"93",
          7311 => x"66",
          7312 => x"26",
          7313 => x"56",
          7314 => x"83",
          7315 => x"64",
          7316 => x"77",
          7317 => x"84",
          7318 => x"52",
          7319 => x"9d",
          7320 => x"d4",
          7321 => x"51",
          7322 => x"3f",
          7323 => x"55",
          7324 => x"81",
          7325 => x"34",
          7326 => x"16",
          7327 => x"16",
          7328 => x"16",
          7329 => x"05",
          7330 => x"c1",
          7331 => x"ff",
          7332 => x"fe",
          7333 => x"34",
          7334 => x"08",
          7335 => x"07",
          7336 => x"16",
          7337 => x"cc",
          7338 => x"34",
          7339 => x"c6",
          7340 => x"9c",
          7341 => x"52",
          7342 => x"51",
          7343 => x"3f",
          7344 => x"53",
          7345 => x"51",
          7346 => x"3f",
          7347 => x"87",
          7348 => x"38",
          7349 => x"52",
          7350 => x"99",
          7351 => x"56",
          7352 => x"08",
          7353 => x"39",
          7354 => x"39",
          7355 => x"39",
          7356 => x"08",
          7357 => x"87",
          7358 => x"3d",
          7359 => x"3d",
          7360 => x"5b",
          7361 => x"60",
          7362 => x"57",
          7363 => x"25",
          7364 => x"3d",
          7365 => x"55",
          7366 => x"15",
          7367 => x"c9",
          7368 => x"81",
          7369 => x"06",
          7370 => x"3d",
          7371 => x"8d",
          7372 => x"74",
          7373 => x"05",
          7374 => x"17",
          7375 => x"2e",
          7376 => x"c9",
          7377 => x"34",
          7378 => x"83",
          7379 => x"74",
          7380 => x"0c",
          7381 => x"04",
          7382 => x"7b",
          7383 => x"b3",
          7384 => x"57",
          7385 => x"09",
          7386 => x"38",
          7387 => x"51",
          7388 => x"17",
          7389 => x"76",
          7390 => x"88",
          7391 => x"17",
          7392 => x"59",
          7393 => x"81",
          7394 => x"76",
          7395 => x"8b",
          7396 => x"54",
          7397 => x"17",
          7398 => x"51",
          7399 => x"79",
          7400 => x"30",
          7401 => x"9f",
          7402 => x"53",
          7403 => x"75",
          7404 => x"81",
          7405 => x"0c",
          7406 => x"04",
          7407 => x"79",
          7408 => x"56",
          7409 => x"24",
          7410 => x"3d",
          7411 => x"74",
          7412 => x"52",
          7413 => x"cb",
          7414 => x"87",
          7415 => x"38",
          7416 => x"78",
          7417 => x"06",
          7418 => x"16",
          7419 => x"39",
          7420 => x"82",
          7421 => x"89",
          7422 => x"fd",
          7423 => x"54",
          7424 => x"80",
          7425 => x"ff",
          7426 => x"76",
          7427 => x"3d",
          7428 => x"3d",
          7429 => x"e3",
          7430 => x"53",
          7431 => x"53",
          7432 => x"3f",
          7433 => x"51",
          7434 => x"72",
          7435 => x"3f",
          7436 => x"04",
          7437 => x"ff",
          7438 => x"ff",
          7439 => x"00",
          7440 => x"ff",
          7441 => x"0e",
          7442 => x"0d",
          7443 => x"0d",
          7444 => x"0d",
          7445 => x"0d",
          7446 => x"0d",
          7447 => x"0d",
          7448 => x"0d",
          7449 => x"0d",
          7450 => x"0d",
          7451 => x"0d",
          7452 => x"0d",
          7453 => x"0d",
          7454 => x"0d",
          7455 => x"0d",
          7456 => x"0d",
          7457 => x"0d",
          7458 => x"0d",
          7459 => x"0d",
          7460 => x"0e",
          7461 => x"25",
          7462 => x"25",
          7463 => x"25",
          7464 => x"25",
          7465 => x"25",
          7466 => x"31",
          7467 => x"32",
          7468 => x"33",
          7469 => x"35",
          7470 => x"32",
          7471 => x"30",
          7472 => x"34",
          7473 => x"35",
          7474 => x"34",
          7475 => x"34",
          7476 => x"34",
          7477 => x"33",
          7478 => x"30",
          7479 => x"33",
          7480 => x"33",
          7481 => x"34",
          7482 => x"30",
          7483 => x"30",
          7484 => x"34",
          7485 => x"34",
          7486 => x"35",
          7487 => x"35",
          7488 => x"6e",
          7489 => x"00",
          7490 => x"6f",
          7491 => x"00",
          7492 => x"6e",
          7493 => x"00",
          7494 => x"6f",
          7495 => x"00",
          7496 => x"78",
          7497 => x"00",
          7498 => x"6c",
          7499 => x"00",
          7500 => x"6f",
          7501 => x"00",
          7502 => x"69",
          7503 => x"00",
          7504 => x"75",
          7505 => x"00",
          7506 => x"62",
          7507 => x"68",
          7508 => x"77",
          7509 => x"64",
          7510 => x"65",
          7511 => x"64",
          7512 => x"65",
          7513 => x"6c",
          7514 => x"00",
          7515 => x"70",
          7516 => x"73",
          7517 => x"74",
          7518 => x"73",
          7519 => x"00",
          7520 => x"66",
          7521 => x"00",
          7522 => x"73",
          7523 => x"00",
          7524 => x"61",
          7525 => x"00",
          7526 => x"61",
          7527 => x"00",
          7528 => x"6c",
          7529 => x"00",
          7530 => x"00",
          7531 => x"73",
          7532 => x"72",
          7533 => x"0a",
          7534 => x"74",
          7535 => x"61",
          7536 => x"72",
          7537 => x"2e",
          7538 => x"00",
          7539 => x"73",
          7540 => x"6f",
          7541 => x"65",
          7542 => x"2e",
          7543 => x"00",
          7544 => x"20",
          7545 => x"65",
          7546 => x"75",
          7547 => x"0a",
          7548 => x"20",
          7549 => x"68",
          7550 => x"75",
          7551 => x"0a",
          7552 => x"76",
          7553 => x"64",
          7554 => x"6c",
          7555 => x"6d",
          7556 => x"00",
          7557 => x"63",
          7558 => x"20",
          7559 => x"69",
          7560 => x"0a",
          7561 => x"6c",
          7562 => x"6c",
          7563 => x"64",
          7564 => x"78",
          7565 => x"73",
          7566 => x"00",
          7567 => x"6c",
          7568 => x"61",
          7569 => x"65",
          7570 => x"76",
          7571 => x"64",
          7572 => x"00",
          7573 => x"20",
          7574 => x"77",
          7575 => x"65",
          7576 => x"6f",
          7577 => x"74",
          7578 => x"0a",
          7579 => x"69",
          7580 => x"6e",
          7581 => x"65",
          7582 => x"73",
          7583 => x"76",
          7584 => x"64",
          7585 => x"00",
          7586 => x"73",
          7587 => x"6f",
          7588 => x"6e",
          7589 => x"65",
          7590 => x"00",
          7591 => x"20",
          7592 => x"70",
          7593 => x"62",
          7594 => x"66",
          7595 => x"73",
          7596 => x"65",
          7597 => x"6f",
          7598 => x"20",
          7599 => x"64",
          7600 => x"2e",
          7601 => x"00",
          7602 => x"72",
          7603 => x"20",
          7604 => x"72",
          7605 => x"2e",
          7606 => x"00",
          7607 => x"6d",
          7608 => x"74",
          7609 => x"70",
          7610 => x"74",
          7611 => x"20",
          7612 => x"63",
          7613 => x"65",
          7614 => x"00",
          7615 => x"6c",
          7616 => x"73",
          7617 => x"63",
          7618 => x"2e",
          7619 => x"00",
          7620 => x"73",
          7621 => x"69",
          7622 => x"6e",
          7623 => x"65",
          7624 => x"79",
          7625 => x"00",
          7626 => x"6f",
          7627 => x"6e",
          7628 => x"70",
          7629 => x"66",
          7630 => x"73",
          7631 => x"00",
          7632 => x"72",
          7633 => x"74",
          7634 => x"20",
          7635 => x"6f",
          7636 => x"63",
          7637 => x"00",
          7638 => x"63",
          7639 => x"73",
          7640 => x"00",
          7641 => x"6b",
          7642 => x"6e",
          7643 => x"72",
          7644 => x"0a",
          7645 => x"6c",
          7646 => x"79",
          7647 => x"20",
          7648 => x"61",
          7649 => x"6c",
          7650 => x"79",
          7651 => x"2f",
          7652 => x"2e",
          7653 => x"00",
          7654 => x"61",
          7655 => x"00",
          7656 => x"38",
          7657 => x"00",
          7658 => x"20",
          7659 => x"34",
          7660 => x"00",
          7661 => x"20",
          7662 => x"20",
          7663 => x"00",
          7664 => x"32",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"0a",
          7669 => x"55",
          7670 => x"00",
          7671 => x"2a",
          7672 => x"20",
          7673 => x"00",
          7674 => x"2f",
          7675 => x"32",
          7676 => x"00",
          7677 => x"2e",
          7678 => x"00",
          7679 => x"50",
          7680 => x"72",
          7681 => x"25",
          7682 => x"29",
          7683 => x"20",
          7684 => x"2a",
          7685 => x"00",
          7686 => x"55",
          7687 => x"49",
          7688 => x"72",
          7689 => x"74",
          7690 => x"6e",
          7691 => x"72",
          7692 => x"00",
          7693 => x"6d",
          7694 => x"69",
          7695 => x"72",
          7696 => x"74",
          7697 => x"00",
          7698 => x"32",
          7699 => x"74",
          7700 => x"75",
          7701 => x"00",
          7702 => x"43",
          7703 => x"52",
          7704 => x"6e",
          7705 => x"72",
          7706 => x"0a",
          7707 => x"43",
          7708 => x"57",
          7709 => x"6e",
          7710 => x"72",
          7711 => x"0a",
          7712 => x"52",
          7713 => x"52",
          7714 => x"6e",
          7715 => x"72",
          7716 => x"0a",
          7717 => x"52",
          7718 => x"54",
          7719 => x"6e",
          7720 => x"72",
          7721 => x"0a",
          7722 => x"52",
          7723 => x"52",
          7724 => x"6e",
          7725 => x"72",
          7726 => x"0a",
          7727 => x"52",
          7728 => x"54",
          7729 => x"6e",
          7730 => x"72",
          7731 => x"0a",
          7732 => x"74",
          7733 => x"67",
          7734 => x"20",
          7735 => x"65",
          7736 => x"2e",
          7737 => x"00",
          7738 => x"61",
          7739 => x"6e",
          7740 => x"69",
          7741 => x"2e",
          7742 => x"00",
          7743 => x"74",
          7744 => x"65",
          7745 => x"61",
          7746 => x"00",
          7747 => x"75",
          7748 => x"68",
          7749 => x"00",
          7750 => x"00",
          7751 => x"69",
          7752 => x"20",
          7753 => x"69",
          7754 => x"69",
          7755 => x"73",
          7756 => x"64",
          7757 => x"72",
          7758 => x"2c",
          7759 => x"65",
          7760 => x"20",
          7761 => x"74",
          7762 => x"6e",
          7763 => x"6c",
          7764 => x"00",
          7765 => x"00",
          7766 => x"64",
          7767 => x"73",
          7768 => x"64",
          7769 => x"00",
          7770 => x"69",
          7771 => x"6c",
          7772 => x"64",
          7773 => x"00",
          7774 => x"69",
          7775 => x"20",
          7776 => x"69",
          7777 => x"69",
          7778 => x"73",
          7779 => x"00",
          7780 => x"3d",
          7781 => x"00",
          7782 => x"3a",
          7783 => x"65",
          7784 => x"6e",
          7785 => x"2e",
          7786 => x"00",
          7787 => x"70",
          7788 => x"67",
          7789 => x"00",
          7790 => x"6d",
          7791 => x"69",
          7792 => x"2e",
          7793 => x"00",
          7794 => x"38",
          7795 => x"25",
          7796 => x"29",
          7797 => x"30",
          7798 => x"28",
          7799 => x"78",
          7800 => x"00",
          7801 => x"6d",
          7802 => x"65",
          7803 => x"79",
          7804 => x"00",
          7805 => x"6f",
          7806 => x"65",
          7807 => x"0a",
          7808 => x"38",
          7809 => x"30",
          7810 => x"00",
          7811 => x"3f",
          7812 => x"00",
          7813 => x"38",
          7814 => x"30",
          7815 => x"00",
          7816 => x"38",
          7817 => x"30",
          7818 => x"00",
          7819 => x"73",
          7820 => x"69",
          7821 => x"69",
          7822 => x"72",
          7823 => x"74",
          7824 => x"00",
          7825 => x"61",
          7826 => x"6e",
          7827 => x"6e",
          7828 => x"72",
          7829 => x"73",
          7830 => x"00",
          7831 => x"73",
          7832 => x"65",
          7833 => x"61",
          7834 => x"66",
          7835 => x"0a",
          7836 => x"61",
          7837 => x"6e",
          7838 => x"61",
          7839 => x"66",
          7840 => x"0a",
          7841 => x"65",
          7842 => x"69",
          7843 => x"63",
          7844 => x"20",
          7845 => x"30",
          7846 => x"2e",
          7847 => x"00",
          7848 => x"6c",
          7849 => x"67",
          7850 => x"64",
          7851 => x"20",
          7852 => x"78",
          7853 => x"2e",
          7854 => x"00",
          7855 => x"6c",
          7856 => x"65",
          7857 => x"6e",
          7858 => x"63",
          7859 => x"20",
          7860 => x"29",
          7861 => x"00",
          7862 => x"73",
          7863 => x"74",
          7864 => x"20",
          7865 => x"6c",
          7866 => x"74",
          7867 => x"2e",
          7868 => x"00",
          7869 => x"6c",
          7870 => x"65",
          7871 => x"74",
          7872 => x"2e",
          7873 => x"00",
          7874 => x"55",
          7875 => x"6e",
          7876 => x"3a",
          7877 => x"5c",
          7878 => x"25",
          7879 => x"00",
          7880 => x"3a",
          7881 => x"5c",
          7882 => x"00",
          7883 => x"3a",
          7884 => x"00",
          7885 => x"64",
          7886 => x"6d",
          7887 => x"64",
          7888 => x"00",
          7889 => x"6e",
          7890 => x"67",
          7891 => x"0a",
          7892 => x"61",
          7893 => x"6e",
          7894 => x"6e",
          7895 => x"72",
          7896 => x"73",
          7897 => x"0a",
          7898 => x"2f",
          7899 => x"25",
          7900 => x"64",
          7901 => x"3a",
          7902 => x"25",
          7903 => x"0a",
          7904 => x"43",
          7905 => x"6e",
          7906 => x"75",
          7907 => x"69",
          7908 => x"00",
          7909 => x"66",
          7910 => x"20",
          7911 => x"20",
          7912 => x"66",
          7913 => x"00",
          7914 => x"44",
          7915 => x"63",
          7916 => x"69",
          7917 => x"65",
          7918 => x"74",
          7919 => x"0a",
          7920 => x"20",
          7921 => x"20",
          7922 => x"41",
          7923 => x"28",
          7924 => x"58",
          7925 => x"38",
          7926 => x"0a",
          7927 => x"20",
          7928 => x"52",
          7929 => x"20",
          7930 => x"28",
          7931 => x"58",
          7932 => x"38",
          7933 => x"0a",
          7934 => x"20",
          7935 => x"53",
          7936 => x"52",
          7937 => x"28",
          7938 => x"58",
          7939 => x"38",
          7940 => x"0a",
          7941 => x"20",
          7942 => x"41",
          7943 => x"20",
          7944 => x"28",
          7945 => x"58",
          7946 => x"38",
          7947 => x"0a",
          7948 => x"20",
          7949 => x"4d",
          7950 => x"20",
          7951 => x"28",
          7952 => x"58",
          7953 => x"38",
          7954 => x"0a",
          7955 => x"20",
          7956 => x"20",
          7957 => x"44",
          7958 => x"28",
          7959 => x"69",
          7960 => x"20",
          7961 => x"32",
          7962 => x"0a",
          7963 => x"20",
          7964 => x"4d",
          7965 => x"20",
          7966 => x"28",
          7967 => x"65",
          7968 => x"20",
          7969 => x"32",
          7970 => x"0a",
          7971 => x"20",
          7972 => x"54",
          7973 => x"54",
          7974 => x"28",
          7975 => x"6e",
          7976 => x"73",
          7977 => x"32",
          7978 => x"0a",
          7979 => x"20",
          7980 => x"53",
          7981 => x"4e",
          7982 => x"55",
          7983 => x"00",
          7984 => x"20",
          7985 => x"20",
          7986 => x"0a",
          7987 => x"20",
          7988 => x"43",
          7989 => x"00",
          7990 => x"20",
          7991 => x"32",
          7992 => x"00",
          7993 => x"20",
          7994 => x"49",
          7995 => x"00",
          7996 => x"64",
          7997 => x"73",
          7998 => x"0a",
          7999 => x"20",
          8000 => x"55",
          8001 => x"73",
          8002 => x"56",
          8003 => x"6f",
          8004 => x"64",
          8005 => x"73",
          8006 => x"20",
          8007 => x"58",
          8008 => x"00",
          8009 => x"20",
          8010 => x"55",
          8011 => x"6d",
          8012 => x"20",
          8013 => x"72",
          8014 => x"64",
          8015 => x"73",
          8016 => x"20",
          8017 => x"58",
          8018 => x"00",
          8019 => x"20",
          8020 => x"61",
          8021 => x"53",
          8022 => x"74",
          8023 => x"64",
          8024 => x"73",
          8025 => x"20",
          8026 => x"20",
          8027 => x"58",
          8028 => x"00",
          8029 => x"73",
          8030 => x"00",
          8031 => x"20",
          8032 => x"55",
          8033 => x"20",
          8034 => x"20",
          8035 => x"20",
          8036 => x"20",
          8037 => x"20",
          8038 => x"20",
          8039 => x"58",
          8040 => x"00",
          8041 => x"20",
          8042 => x"73",
          8043 => x"20",
          8044 => x"63",
          8045 => x"72",
          8046 => x"20",
          8047 => x"20",
          8048 => x"20",
          8049 => x"25",
          8050 => x"4d",
          8051 => x"00",
          8052 => x"20",
          8053 => x"52",
          8054 => x"43",
          8055 => x"6b",
          8056 => x"65",
          8057 => x"20",
          8058 => x"20",
          8059 => x"20",
          8060 => x"25",
          8061 => x"4d",
          8062 => x"00",
          8063 => x"20",
          8064 => x"73",
          8065 => x"6e",
          8066 => x"44",
          8067 => x"20",
          8068 => x"63",
          8069 => x"72",
          8070 => x"20",
          8071 => x"25",
          8072 => x"4d",
          8073 => x"00",
          8074 => x"61",
          8075 => x"00",
          8076 => x"64",
          8077 => x"00",
          8078 => x"65",
          8079 => x"00",
          8080 => x"4f",
          8081 => x"4f",
          8082 => x"00",
          8083 => x"6b",
          8084 => x"6e",
          8085 => x"7f",
          8086 => x"00",
          8087 => x"00",
          8088 => x"7f",
          8089 => x"00",
          8090 => x"00",
          8091 => x"7f",
          8092 => x"00",
          8093 => x"00",
          8094 => x"7f",
          8095 => x"00",
          8096 => x"00",
          8097 => x"7f",
          8098 => x"00",
          8099 => x"00",
          8100 => x"7f",
          8101 => x"00",
          8102 => x"00",
          8103 => x"7f",
          8104 => x"00",
          8105 => x"00",
          8106 => x"7f",
          8107 => x"00",
          8108 => x"00",
          8109 => x"7f",
          8110 => x"00",
          8111 => x"00",
          8112 => x"7f",
          8113 => x"00",
          8114 => x"00",
          8115 => x"7f",
          8116 => x"00",
          8117 => x"00",
          8118 => x"7f",
          8119 => x"00",
          8120 => x"00",
          8121 => x"7f",
          8122 => x"00",
          8123 => x"00",
          8124 => x"7f",
          8125 => x"00",
          8126 => x"00",
          8127 => x"7f",
          8128 => x"00",
          8129 => x"00",
          8130 => x"7f",
          8131 => x"00",
          8132 => x"00",
          8133 => x"7f",
          8134 => x"00",
          8135 => x"00",
          8136 => x"7f",
          8137 => x"00",
          8138 => x"00",
          8139 => x"7f",
          8140 => x"00",
          8141 => x"00",
          8142 => x"7f",
          8143 => x"00",
          8144 => x"00",
          8145 => x"7f",
          8146 => x"00",
          8147 => x"00",
          8148 => x"7f",
          8149 => x"00",
          8150 => x"00",
          8151 => x"44",
          8152 => x"43",
          8153 => x"42",
          8154 => x"41",
          8155 => x"36",
          8156 => x"35",
          8157 => x"34",
          8158 => x"46",
          8159 => x"33",
          8160 => x"32",
          8161 => x"31",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"73",
          8174 => x"79",
          8175 => x"73",
          8176 => x"00",
          8177 => x"00",
          8178 => x"34",
          8179 => x"25",
          8180 => x"00",
          8181 => x"69",
          8182 => x"20",
          8183 => x"72",
          8184 => x"74",
          8185 => x"65",
          8186 => x"73",
          8187 => x"79",
          8188 => x"6c",
          8189 => x"6f",
          8190 => x"46",
          8191 => x"00",
          8192 => x"6e",
          8193 => x"20",
          8194 => x"6e",
          8195 => x"65",
          8196 => x"20",
          8197 => x"74",
          8198 => x"20",
          8199 => x"65",
          8200 => x"69",
          8201 => x"6c",
          8202 => x"2e",
          8203 => x"00",
          8204 => x"00",
          8205 => x"2b",
          8206 => x"3c",
          8207 => x"5b",
          8208 => x"00",
          8209 => x"54",
          8210 => x"54",
          8211 => x"00",
          8212 => x"90",
          8213 => x"4f",
          8214 => x"30",
          8215 => x"20",
          8216 => x"45",
          8217 => x"20",
          8218 => x"33",
          8219 => x"20",
          8220 => x"20",
          8221 => x"45",
          8222 => x"20",
          8223 => x"20",
          8224 => x"20",
          8225 => x"80",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"45",
          8230 => x"8f",
          8231 => x"45",
          8232 => x"8e",
          8233 => x"92",
          8234 => x"55",
          8235 => x"9a",
          8236 => x"9e",
          8237 => x"4f",
          8238 => x"a6",
          8239 => x"aa",
          8240 => x"ae",
          8241 => x"b2",
          8242 => x"b6",
          8243 => x"ba",
          8244 => x"be",
          8245 => x"c2",
          8246 => x"c6",
          8247 => x"ca",
          8248 => x"ce",
          8249 => x"d2",
          8250 => x"d6",
          8251 => x"da",
          8252 => x"de",
          8253 => x"e2",
          8254 => x"e6",
          8255 => x"ea",
          8256 => x"ee",
          8257 => x"f2",
          8258 => x"f6",
          8259 => x"fa",
          8260 => x"fe",
          8261 => x"2c",
          8262 => x"5d",
          8263 => x"2a",
          8264 => x"3f",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"02",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"75",
          8276 => x"01",
          8277 => x"00",
          8278 => x"00",
          8279 => x"75",
          8280 => x"01",
          8281 => x"00",
          8282 => x"00",
          8283 => x"75",
          8284 => x"03",
          8285 => x"00",
          8286 => x"00",
          8287 => x"75",
          8288 => x"03",
          8289 => x"00",
          8290 => x"00",
          8291 => x"75",
          8292 => x"03",
          8293 => x"00",
          8294 => x"00",
          8295 => x"75",
          8296 => x"04",
          8297 => x"00",
          8298 => x"00",
          8299 => x"75",
          8300 => x"04",
          8301 => x"00",
          8302 => x"00",
          8303 => x"75",
          8304 => x"04",
          8305 => x"00",
          8306 => x"00",
          8307 => x"75",
          8308 => x"04",
          8309 => x"00",
          8310 => x"00",
          8311 => x"75",
          8312 => x"04",
          8313 => x"00",
          8314 => x"00",
          8315 => x"75",
          8316 => x"04",
          8317 => x"00",
          8318 => x"00",
          8319 => x"75",
          8320 => x"04",
          8321 => x"00",
          8322 => x"00",
          8323 => x"75",
          8324 => x"05",
          8325 => x"00",
          8326 => x"00",
          8327 => x"75",
          8328 => x"05",
          8329 => x"00",
          8330 => x"00",
          8331 => x"75",
          8332 => x"05",
          8333 => x"00",
          8334 => x"00",
          8335 => x"75",
          8336 => x"05",
          8337 => x"00",
          8338 => x"00",
          8339 => x"75",
          8340 => x"07",
          8341 => x"00",
          8342 => x"00",
          8343 => x"75",
          8344 => x"07",
          8345 => x"00",
          8346 => x"00",
          8347 => x"75",
          8348 => x"08",
          8349 => x"00",
          8350 => x"00",
          8351 => x"75",
          8352 => x"08",
          8353 => x"00",
          8354 => x"00",
          8355 => x"75",
          8356 => x"08",
          8357 => x"00",
          8358 => x"00",
          8359 => x"75",
          8360 => x"08",
          8361 => x"00",
          8362 => x"00",
          8363 => x"75",
          8364 => x"09",
          8365 => x"00",
          8366 => x"00",
          8367 => x"75",
          8368 => x"09",
          8369 => x"00",
          8370 => x"00",
          8371 => x"75",
          8372 => x"09",
          8373 => x"00",
          8374 => x"00",
          8375 => x"75",
          8376 => x"09",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"7f",
          8382 => x"00",
          8383 => x"7f",
          8384 => x"00",
          8385 => x"7f",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"ff",
          8390 => x"00",
          8391 => x"00",
          8392 => x"78",
          8393 => x"00",
          8394 => x"e1",
          8395 => x"e1",
          8396 => x"e1",
          8397 => x"00",
          8398 => x"01",
          8399 => x"01",
          8400 => x"10",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"7f",
          8427 => x"00",
          8428 => x"7f",
          8429 => x"00",
          8430 => x"7f",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"e5",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"be",
           387 => x"87",
           388 => x"a0",
           389 => x"87",
           390 => x"cb",
           391 => x"87",
           392 => x"a0",
           393 => x"87",
           394 => x"cc",
           395 => x"87",
           396 => x"a0",
           397 => x"87",
           398 => x"cc",
           399 => x"87",
           400 => x"a0",
           401 => x"87",
           402 => x"d2",
           403 => x"87",
           404 => x"a0",
           405 => x"87",
           406 => x"d3",
           407 => x"87",
           408 => x"a0",
           409 => x"87",
           410 => x"cc",
           411 => x"87",
           412 => x"a0",
           413 => x"87",
           414 => x"d3",
           415 => x"87",
           416 => x"a0",
           417 => x"87",
           418 => x"d5",
           419 => x"87",
           420 => x"a0",
           421 => x"87",
           422 => x"d2",
           423 => x"87",
           424 => x"a0",
           425 => x"87",
           426 => x"cc",
           427 => x"87",
           428 => x"a0",
           429 => x"87",
           430 => x"d2",
           431 => x"87",
           432 => x"a0",
           433 => x"87",
           434 => x"d2",
           435 => x"87",
           436 => x"a0",
           437 => x"87",
           438 => x"c0",
           439 => x"87",
           440 => x"a0",
           441 => x"87",
           442 => x"c0",
           443 => x"87",
           444 => x"a0",
           445 => x"87",
           446 => x"d3",
           447 => x"d8",
           448 => x"90",
           449 => x"d8",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"82",
           455 => x"82",
           456 => x"82",
           457 => x"81",
           458 => x"82",
           459 => x"82",
           460 => x"82",
           461 => x"81",
           462 => x"82",
           463 => x"82",
           464 => x"82",
           465 => x"81",
           466 => x"82",
           467 => x"82",
           468 => x"82",
           469 => x"81",
           470 => x"82",
           471 => x"82",
           472 => x"82",
           473 => x"81",
           474 => x"82",
           475 => x"82",
           476 => x"82",
           477 => x"81",
           478 => x"82",
           479 => x"82",
           480 => x"82",
           481 => x"81",
           482 => x"82",
           483 => x"82",
           484 => x"82",
           485 => x"81",
           486 => x"82",
           487 => x"82",
           488 => x"82",
           489 => x"81",
           490 => x"82",
           491 => x"82",
           492 => x"82",
           493 => x"81",
           494 => x"82",
           495 => x"82",
           496 => x"82",
           497 => x"81",
           498 => x"82",
           499 => x"82",
           500 => x"82",
           501 => x"81",
           502 => x"82",
           503 => x"82",
           504 => x"82",
           505 => x"81",
           506 => x"82",
           507 => x"82",
           508 => x"82",
           509 => x"81",
           510 => x"82",
           511 => x"82",
           512 => x"82",
           513 => x"81",
           514 => x"82",
           515 => x"82",
           516 => x"82",
           517 => x"81",
           518 => x"82",
           519 => x"82",
           520 => x"82",
           521 => x"81",
           522 => x"82",
           523 => x"82",
           524 => x"82",
           525 => x"81",
           526 => x"82",
           527 => x"82",
           528 => x"82",
           529 => x"81",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"81",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"81",
           538 => x"82",
           539 => x"82",
           540 => x"82",
           541 => x"81",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"81",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"81",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"81",
           554 => x"82",
           555 => x"82",
           556 => x"82",
           557 => x"81",
           558 => x"82",
           559 => x"82",
           560 => x"82",
           561 => x"81",
           562 => x"82",
           563 => x"82",
           564 => x"82",
           565 => x"80",
           566 => x"82",
           567 => x"82",
           568 => x"82",
           569 => x"80",
           570 => x"82",
           571 => x"82",
           572 => x"82",
           573 => x"80",
           574 => x"82",
           575 => x"82",
           576 => x"82",
           577 => x"b8",
           578 => x"87",
           579 => x"a0",
           580 => x"87",
           581 => x"a0",
           582 => x"d8",
           583 => x"90",
           584 => x"d8",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"82",
           590 => x"82",
           591 => x"3c",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"51",
           601 => x"73",
           602 => x"73",
           603 => x"81",
           604 => x"10",
           605 => x"07",
           606 => x"0c",
           607 => x"72",
           608 => x"81",
           609 => x"09",
           610 => x"71",
           611 => x"0a",
           612 => x"72",
           613 => x"51",
           614 => x"82",
           615 => x"82",
           616 => x"8e",
           617 => x"70",
           618 => x"0c",
           619 => x"93",
           620 => x"81",
           621 => x"04",
           622 => x"d8",
           623 => x"87",
           624 => x"3d",
           625 => x"d8",
           626 => x"08",
           627 => x"08",
           628 => x"82",
           629 => x"fc",
           630 => x"71",
           631 => x"d8",
           632 => x"08",
           633 => x"87",
           634 => x"05",
           635 => x"ff",
           636 => x"70",
           637 => x"38",
           638 => x"87",
           639 => x"05",
           640 => x"82",
           641 => x"fc",
           642 => x"87",
           643 => x"05",
           644 => x"d8",
           645 => x"08",
           646 => x"87",
           647 => x"84",
           648 => x"87",
           649 => x"82",
           650 => x"02",
           651 => x"0c",
           652 => x"82",
           653 => x"88",
           654 => x"87",
           655 => x"05",
           656 => x"d8",
           657 => x"08",
           658 => x"82",
           659 => x"8c",
           660 => x"05",
           661 => x"08",
           662 => x"82",
           663 => x"fc",
           664 => x"51",
           665 => x"82",
           666 => x"fc",
           667 => x"05",
           668 => x"08",
           669 => x"70",
           670 => x"51",
           671 => x"84",
           672 => x"39",
           673 => x"08",
           674 => x"70",
           675 => x"0c",
           676 => x"0d",
           677 => x"0c",
           678 => x"d8",
           679 => x"87",
           680 => x"3d",
           681 => x"d8",
           682 => x"08",
           683 => x"08",
           684 => x"82",
           685 => x"8c",
           686 => x"87",
           687 => x"05",
           688 => x"d8",
           689 => x"08",
           690 => x"e5",
           691 => x"d8",
           692 => x"08",
           693 => x"87",
           694 => x"05",
           695 => x"d8",
           696 => x"08",
           697 => x"87",
           698 => x"05",
           699 => x"d8",
           700 => x"08",
           701 => x"38",
           702 => x"08",
           703 => x"51",
           704 => x"87",
           705 => x"05",
           706 => x"82",
           707 => x"f8",
           708 => x"87",
           709 => x"05",
           710 => x"71",
           711 => x"87",
           712 => x"05",
           713 => x"82",
           714 => x"fc",
           715 => x"ad",
           716 => x"d8",
           717 => x"08",
           718 => x"cc",
           719 => x"3d",
           720 => x"d8",
           721 => x"87",
           722 => x"82",
           723 => x"fd",
           724 => x"87",
           725 => x"05",
           726 => x"81",
           727 => x"87",
           728 => x"05",
           729 => x"33",
           730 => x"08",
           731 => x"81",
           732 => x"d8",
           733 => x"0c",
           734 => x"08",
           735 => x"70",
           736 => x"ff",
           737 => x"54",
           738 => x"2e",
           739 => x"ce",
           740 => x"d8",
           741 => x"08",
           742 => x"82",
           743 => x"88",
           744 => x"05",
           745 => x"08",
           746 => x"70",
           747 => x"51",
           748 => x"38",
           749 => x"87",
           750 => x"05",
           751 => x"39",
           752 => x"08",
           753 => x"ff",
           754 => x"d8",
           755 => x"0c",
           756 => x"08",
           757 => x"80",
           758 => x"ff",
           759 => x"87",
           760 => x"05",
           761 => x"80",
           762 => x"87",
           763 => x"05",
           764 => x"52",
           765 => x"38",
           766 => x"87",
           767 => x"05",
           768 => x"39",
           769 => x"08",
           770 => x"ff",
           771 => x"d8",
           772 => x"0c",
           773 => x"08",
           774 => x"70",
           775 => x"70",
           776 => x"0b",
           777 => x"08",
           778 => x"ae",
           779 => x"d8",
           780 => x"08",
           781 => x"87",
           782 => x"05",
           783 => x"72",
           784 => x"82",
           785 => x"fc",
           786 => x"55",
           787 => x"8a",
           788 => x"82",
           789 => x"fc",
           790 => x"87",
           791 => x"05",
           792 => x"cc",
           793 => x"0d",
           794 => x"0c",
           795 => x"d8",
           796 => x"87",
           797 => x"3d",
           798 => x"d8",
           799 => x"08",
           800 => x"08",
           801 => x"82",
           802 => x"90",
           803 => x"2e",
           804 => x"82",
           805 => x"90",
           806 => x"05",
           807 => x"08",
           808 => x"82",
           809 => x"90",
           810 => x"05",
           811 => x"08",
           812 => x"82",
           813 => x"90",
           814 => x"2e",
           815 => x"87",
           816 => x"05",
           817 => x"82",
           818 => x"fc",
           819 => x"52",
           820 => x"82",
           821 => x"fc",
           822 => x"05",
           823 => x"08",
           824 => x"ff",
           825 => x"87",
           826 => x"05",
           827 => x"87",
           828 => x"84",
           829 => x"87",
           830 => x"f9",
           831 => x"70",
           832 => x"56",
           833 => x"2e",
           834 => x"95",
           835 => x"51",
           836 => x"82",
           837 => x"15",
           838 => x"16",
           839 => x"cd",
           840 => x"54",
           841 => x"09",
           842 => x"38",
           843 => x"f1",
           844 => x"76",
           845 => x"82",
           846 => x"08",
           847 => x"f9",
           848 => x"cc",
           849 => x"52",
           850 => x"fb",
           851 => x"87",
           852 => x"38",
           853 => x"54",
           854 => x"ff",
           855 => x"17",
           856 => x"06",
           857 => x"77",
           858 => x"ff",
           859 => x"87",
           860 => x"3d",
           861 => x"3d",
           862 => x"71",
           863 => x"8e",
           864 => x"29",
           865 => x"05",
           866 => x"04",
           867 => x"51",
           868 => x"81",
           869 => x"80",
           870 => x"eb",
           871 => x"f2",
           872 => x"e0",
           873 => x"39",
           874 => x"51",
           875 => x"81",
           876 => x"80",
           877 => x"ec",
           878 => x"d6",
           879 => x"a4",
           880 => x"39",
           881 => x"51",
           882 => x"81",
           883 => x"80",
           884 => x"ec",
           885 => x"39",
           886 => x"51",
           887 => x"ed",
           888 => x"39",
           889 => x"51",
           890 => x"ed",
           891 => x"39",
           892 => x"51",
           893 => x"ee",
           894 => x"39",
           895 => x"51",
           896 => x"ee",
           897 => x"39",
           898 => x"51",
           899 => x"ee",
           900 => x"8e",
           901 => x"0d",
           902 => x"0d",
           903 => x"56",
           904 => x"26",
           905 => x"52",
           906 => x"29",
           907 => x"87",
           908 => x"51",
           909 => x"3f",
           910 => x"08",
           911 => x"80",
           912 => x"82",
           913 => x"54",
           914 => x"52",
           915 => x"51",
           916 => x"87",
           917 => x"ec",
           918 => x"02",
           919 => x"e3",
           920 => x"57",
           921 => x"30",
           922 => x"73",
           923 => x"59",
           924 => x"77",
           925 => x"83",
           926 => x"74",
           927 => x"81",
           928 => x"55",
           929 => x"81",
           930 => x"53",
           931 => x"3d",
           932 => x"81",
           933 => x"82",
           934 => x"57",
           935 => x"08",
           936 => x"87",
           937 => x"c0",
           938 => x"82",
           939 => x"59",
           940 => x"05",
           941 => x"53",
           942 => x"51",
           943 => x"3f",
           944 => x"08",
           945 => x"cc",
           946 => x"7a",
           947 => x"2e",
           948 => x"19",
           949 => x"59",
           950 => x"3d",
           951 => x"81",
           952 => x"76",
           953 => x"07",
           954 => x"30",
           955 => x"72",
           956 => x"51",
           957 => x"2e",
           958 => x"ef",
           959 => x"c0",
           960 => x"52",
           961 => x"91",
           962 => x"75",
           963 => x"0c",
           964 => x"04",
           965 => x"7b",
           966 => x"b3",
           967 => x"58",
           968 => x"53",
           969 => x"51",
           970 => x"82",
           971 => x"a4",
           972 => x"2e",
           973 => x"81",
           974 => x"98",
           975 => x"7f",
           976 => x"cc",
           977 => x"7d",
           978 => x"82",
           979 => x"57",
           980 => x"04",
           981 => x"cc",
           982 => x"0d",
           983 => x"0d",
           984 => x"02",
           985 => x"cf",
           986 => x"73",
           987 => x"5f",
           988 => x"5e",
           989 => x"81",
           990 => x"b3",
           991 => x"ef",
           992 => x"9e",
           993 => x"74",
           994 => x"f4",
           995 => x"2e",
           996 => x"a0",
           997 => x"80",
           998 => x"18",
           999 => x"27",
          1000 => x"22",
          1001 => x"ac",
          1002 => x"3f",
          1003 => x"ef",
          1004 => x"ee",
          1005 => x"55",
          1006 => x"18",
          1007 => x"27",
          1008 => x"08",
          1009 => x"a0",
          1010 => x"3f",
          1011 => x"ef",
          1012 => x"ce",
          1013 => x"55",
          1014 => x"18",
          1015 => x"27",
          1016 => x"33",
          1017 => x"c0",
          1018 => x"3f",
          1019 => x"ef",
          1020 => x"ae",
          1021 => x"55",
          1022 => x"c9",
          1023 => x"39",
          1024 => x"51",
          1025 => x"80",
          1026 => x"27",
          1027 => x"18",
          1028 => x"53",
          1029 => x"7a",
          1030 => x"81",
          1031 => x"9f",
          1032 => x"38",
          1033 => x"73",
          1034 => x"ff",
          1035 => x"72",
          1036 => x"38",
          1037 => x"26",
          1038 => x"51",
          1039 => x"51",
          1040 => x"81",
          1041 => x"39",
          1042 => x"51",
          1043 => x"78",
          1044 => x"5c",
          1045 => x"3f",
          1046 => x"08",
          1047 => x"98",
          1048 => x"76",
          1049 => x"81",
          1050 => x"a0",
          1051 => x"87",
          1052 => x"2b",
          1053 => x"70",
          1054 => x"30",
          1055 => x"70",
          1056 => x"07",
          1057 => x"06",
          1058 => x"59",
          1059 => x"80",
          1060 => x"38",
          1061 => x"09",
          1062 => x"38",
          1063 => x"39",
          1064 => x"72",
          1065 => x"cd",
          1066 => x"72",
          1067 => x"0c",
          1068 => x"04",
          1069 => x"02",
          1070 => x"81",
          1071 => x"81",
          1072 => x"55",
          1073 => x"82",
          1074 => x"51",
          1075 => x"81",
          1076 => x"81",
          1077 => x"82",
          1078 => x"52",
          1079 => x"51",
          1080 => x"74",
          1081 => x"38",
          1082 => x"86",
          1083 => x"fe",
          1084 => x"c0",
          1085 => x"53",
          1086 => x"81",
          1087 => x"3f",
          1088 => x"51",
          1089 => x"80",
          1090 => x"3f",
          1091 => x"70",
          1092 => x"52",
          1093 => x"92",
          1094 => x"9a",
          1095 => x"f0",
          1096 => x"e5",
          1097 => x"9a",
          1098 => x"82",
          1099 => x"06",
          1100 => x"80",
          1101 => x"81",
          1102 => x"3f",
          1103 => x"51",
          1104 => x"80",
          1105 => x"3f",
          1106 => x"70",
          1107 => x"52",
          1108 => x"92",
          1109 => x"9a",
          1110 => x"f0",
          1111 => x"a9",
          1112 => x"9a",
          1113 => x"84",
          1114 => x"06",
          1115 => x"80",
          1116 => x"81",
          1117 => x"3f",
          1118 => x"51",
          1119 => x"80",
          1120 => x"3f",
          1121 => x"70",
          1122 => x"52",
          1123 => x"92",
          1124 => x"99",
          1125 => x"f1",
          1126 => x"ed",
          1127 => x"99",
          1128 => x"86",
          1129 => x"06",
          1130 => x"80",
          1131 => x"81",
          1132 => x"3f",
          1133 => x"51",
          1134 => x"80",
          1135 => x"3f",
          1136 => x"70",
          1137 => x"52",
          1138 => x"92",
          1139 => x"99",
          1140 => x"f1",
          1141 => x"b1",
          1142 => x"99",
          1143 => x"88",
          1144 => x"06",
          1145 => x"80",
          1146 => x"81",
          1147 => x"3f",
          1148 => x"51",
          1149 => x"80",
          1150 => x"3f",
          1151 => x"84",
          1152 => x"fb",
          1153 => x"02",
          1154 => x"05",
          1155 => x"56",
          1156 => x"75",
          1157 => x"3f",
          1158 => x"82",
          1159 => x"73",
          1160 => x"53",
          1161 => x"52",
          1162 => x"51",
          1163 => x"3f",
          1164 => x"08",
          1165 => x"87",
          1166 => x"80",
          1167 => x"31",
          1168 => x"73",
          1169 => x"82",
          1170 => x"0b",
          1171 => x"33",
          1172 => x"2e",
          1173 => x"af",
          1174 => x"ac",
          1175 => x"75",
          1176 => x"9b",
          1177 => x"cc",
          1178 => x"8b",
          1179 => x"cc",
          1180 => x"ae",
          1181 => x"82",
          1182 => x"81",
          1183 => x"82",
          1184 => x"82",
          1185 => x"0b",
          1186 => x"c8",
          1187 => x"82",
          1188 => x"06",
          1189 => x"f2",
          1190 => x"52",
          1191 => x"ba",
          1192 => x"82",
          1193 => x"87",
          1194 => x"ce",
          1195 => x"70",
          1196 => x"a8",
          1197 => x"81",
          1198 => x"80",
          1199 => x"82",
          1200 => x"81",
          1201 => x"78",
          1202 => x"81",
          1203 => x"81",
          1204 => x"96",
          1205 => x"59",
          1206 => x"7c",
          1207 => x"82",
          1208 => x"81",
          1209 => x"82",
          1210 => x"7d",
          1211 => x"81",
          1212 => x"91",
          1213 => x"70",
          1214 => x"f2",
          1215 => x"a2",
          1216 => x"70",
          1217 => x"f8",
          1218 => x"fd",
          1219 => x"3d",
          1220 => x"51",
          1221 => x"82",
          1222 => x"90",
          1223 => x"2c",
          1224 => x"80",
          1225 => x"d1",
          1226 => x"c1",
          1227 => x"38",
          1228 => x"83",
          1229 => x"ab",
          1230 => x"78",
          1231 => x"b3",
          1232 => x"24",
          1233 => x"80",
          1234 => x"38",
          1235 => x"78",
          1236 => x"83",
          1237 => x"2e",
          1238 => x"8e",
          1239 => x"bd",
          1240 => x"38",
          1241 => x"90",
          1242 => x"2e",
          1243 => x"78",
          1244 => x"83",
          1245 => x"39",
          1246 => x"85",
          1247 => x"80",
          1248 => x"b7",
          1249 => x"39",
          1250 => x"2e",
          1251 => x"78",
          1252 => x"b0",
          1253 => x"d0",
          1254 => x"38",
          1255 => x"24",
          1256 => x"80",
          1257 => x"f2",
          1258 => x"c3",
          1259 => x"38",
          1260 => x"78",
          1261 => x"8c",
          1262 => x"80",
          1263 => x"ba",
          1264 => x"39",
          1265 => x"2e",
          1266 => x"78",
          1267 => x"92",
          1268 => x"f8",
          1269 => x"38",
          1270 => x"2e",
          1271 => x"8d",
          1272 => x"81",
          1273 => x"b5",
          1274 => x"85",
          1275 => x"38",
          1276 => x"b4",
          1277 => x"11",
          1278 => x"05",
          1279 => x"3f",
          1280 => x"08",
          1281 => x"f2",
          1282 => x"9d",
          1283 => x"fe",
          1284 => x"ff",
          1285 => x"ab",
          1286 => x"87",
          1287 => x"2e",
          1288 => x"63",
          1289 => x"80",
          1290 => x"cb",
          1291 => x"02",
          1292 => x"33",
          1293 => x"bd",
          1294 => x"cc",
          1295 => x"06",
          1296 => x"38",
          1297 => x"51",
          1298 => x"81",
          1299 => x"39",
          1300 => x"51",
          1301 => x"b4",
          1302 => x"11",
          1303 => x"05",
          1304 => x"3f",
          1305 => x"08",
          1306 => x"8e",
          1307 => x"80",
          1308 => x"cf",
          1309 => x"80",
          1310 => x"82",
          1311 => x"52",
          1312 => x"51",
          1313 => x"b4",
          1314 => x"11",
          1315 => x"05",
          1316 => x"3f",
          1317 => x"08",
          1318 => x"38",
          1319 => x"fc",
          1320 => x"3d",
          1321 => x"53",
          1322 => x"51",
          1323 => x"82",
          1324 => x"86",
          1325 => x"cc",
          1326 => x"53",
          1327 => x"52",
          1328 => x"d8",
          1329 => x"cb",
          1330 => x"79",
          1331 => x"b4",
          1332 => x"d8",
          1333 => x"80",
          1334 => x"87",
          1335 => x"8c",
          1336 => x"e8",
          1337 => x"3f",
          1338 => x"8e",
          1339 => x"ff",
          1340 => x"8f",
          1341 => x"87",
          1342 => x"3d",
          1343 => x"52",
          1344 => x"3f",
          1345 => x"87",
          1346 => x"7a",
          1347 => x"3f",
          1348 => x"b4",
          1349 => x"05",
          1350 => x"3f",
          1351 => x"08",
          1352 => x"84",
          1353 => x"8f",
          1354 => x"87",
          1355 => x"3d",
          1356 => x"52",
          1357 => x"3f",
          1358 => x"08",
          1359 => x"84",
          1360 => x"8f",
          1361 => x"85",
          1362 => x"87",
          1363 => x"56",
          1364 => x"87",
          1365 => x"ff",
          1366 => x"53",
          1367 => x"51",
          1368 => x"82",
          1369 => x"80",
          1370 => x"38",
          1371 => x"08",
          1372 => x"3f",
          1373 => x"b4",
          1374 => x"11",
          1375 => x"05",
          1376 => x"3f",
          1377 => x"08",
          1378 => x"ee",
          1379 => x"fe",
          1380 => x"ff",
          1381 => x"a8",
          1382 => x"87",
          1383 => x"2e",
          1384 => x"b4",
          1385 => x"11",
          1386 => x"05",
          1387 => x"3f",
          1388 => x"08",
          1389 => x"87",
          1390 => x"81",
          1391 => x"a0",
          1392 => x"63",
          1393 => x"7b",
          1394 => x"38",
          1395 => x"7a",
          1396 => x"5c",
          1397 => x"26",
          1398 => x"d8",
          1399 => x"ff",
          1400 => x"ff",
          1401 => x"a8",
          1402 => x"87",
          1403 => x"2e",
          1404 => x"b4",
          1405 => x"11",
          1406 => x"05",
          1407 => x"3f",
          1408 => x"08",
          1409 => x"f2",
          1410 => x"fe",
          1411 => x"ff",
          1412 => x"a7",
          1413 => x"87",
          1414 => x"2e",
          1415 => x"81",
          1416 => x"9f",
          1417 => x"5a",
          1418 => x"81",
          1419 => x"59",
          1420 => x"05",
          1421 => x"34",
          1422 => x"42",
          1423 => x"3d",
          1424 => x"53",
          1425 => x"51",
          1426 => x"82",
          1427 => x"80",
          1428 => x"38",
          1429 => x"fc",
          1430 => x"84",
          1431 => x"9b",
          1432 => x"cc",
          1433 => x"f9",
          1434 => x"3d",
          1435 => x"53",
          1436 => x"51",
          1437 => x"82",
          1438 => x"80",
          1439 => x"38",
          1440 => x"51",
          1441 => x"63",
          1442 => x"27",
          1443 => x"70",
          1444 => x"5e",
          1445 => x"7c",
          1446 => x"78",
          1447 => x"79",
          1448 => x"52",
          1449 => x"51",
          1450 => x"81",
          1451 => x"05",
          1452 => x"39",
          1453 => x"51",
          1454 => x"b4",
          1455 => x"11",
          1456 => x"05",
          1457 => x"3f",
          1458 => x"08",
          1459 => x"82",
          1460 => x"59",
          1461 => x"89",
          1462 => x"f0",
          1463 => x"cd",
          1464 => x"b9",
          1465 => x"80",
          1466 => x"82",
          1467 => x"44",
          1468 => x"86",
          1469 => x"78",
          1470 => x"38",
          1471 => x"08",
          1472 => x"82",
          1473 => x"59",
          1474 => x"88",
          1475 => x"88",
          1476 => x"39",
          1477 => x"33",
          1478 => x"2e",
          1479 => x"86",
          1480 => x"89",
          1481 => x"a0",
          1482 => x"05",
          1483 => x"fe",
          1484 => x"ff",
          1485 => x"a5",
          1486 => x"87",
          1487 => x"de",
          1488 => x"b8",
          1489 => x"80",
          1490 => x"82",
          1491 => x"43",
          1492 => x"82",
          1493 => x"59",
          1494 => x"88",
          1495 => x"fc",
          1496 => x"39",
          1497 => x"33",
          1498 => x"2e",
          1499 => x"86",
          1500 => x"aa",
          1501 => x"bb",
          1502 => x"80",
          1503 => x"82",
          1504 => x"43",
          1505 => x"86",
          1506 => x"78",
          1507 => x"38",
          1508 => x"08",
          1509 => x"82",
          1510 => x"88",
          1511 => x"3d",
          1512 => x"53",
          1513 => x"51",
          1514 => x"82",
          1515 => x"80",
          1516 => x"80",
          1517 => x"7a",
          1518 => x"38",
          1519 => x"90",
          1520 => x"70",
          1521 => x"2a",
          1522 => x"51",
          1523 => x"78",
          1524 => x"38",
          1525 => x"83",
          1526 => x"81",
          1527 => x"9c",
          1528 => x"55",
          1529 => x"53",
          1530 => x"51",
          1531 => x"81",
          1532 => x"9c",
          1533 => x"82",
          1534 => x"ff",
          1535 => x"ff",
          1536 => x"a3",
          1537 => x"87",
          1538 => x"2e",
          1539 => x"b4",
          1540 => x"11",
          1541 => x"05",
          1542 => x"3f",
          1543 => x"08",
          1544 => x"38",
          1545 => x"80",
          1546 => x"79",
          1547 => x"05",
          1548 => x"fe",
          1549 => x"ff",
          1550 => x"a3",
          1551 => x"87",
          1552 => x"38",
          1553 => x"63",
          1554 => x"52",
          1555 => x"51",
          1556 => x"80",
          1557 => x"51",
          1558 => x"79",
          1559 => x"59",
          1560 => x"f5",
          1561 => x"79",
          1562 => x"b4",
          1563 => x"11",
          1564 => x"05",
          1565 => x"3f",
          1566 => x"08",
          1567 => x"38",
          1568 => x"80",
          1569 => x"79",
          1570 => x"05",
          1571 => x"39",
          1572 => x"51",
          1573 => x"ff",
          1574 => x"3d",
          1575 => x"53",
          1576 => x"51",
          1577 => x"82",
          1578 => x"80",
          1579 => x"38",
          1580 => x"f0",
          1581 => x"84",
          1582 => x"b1",
          1583 => x"cc",
          1584 => x"a5",
          1585 => x"02",
          1586 => x"79",
          1587 => x"5b",
          1588 => x"b4",
          1589 => x"11",
          1590 => x"05",
          1591 => x"3f",
          1592 => x"08",
          1593 => x"92",
          1594 => x"22",
          1595 => x"f4",
          1596 => x"92",
          1597 => x"52",
          1598 => x"e4",
          1599 => x"79",
          1600 => x"ae",
          1601 => x"38",
          1602 => x"87",
          1603 => x"05",
          1604 => x"b4",
          1605 => x"11",
          1606 => x"05",
          1607 => x"3f",
          1608 => x"08",
          1609 => x"38",
          1610 => x"be",
          1611 => x"70",
          1612 => x"23",
          1613 => x"b1",
          1614 => x"8c",
          1615 => x"3f",
          1616 => x"b4",
          1617 => x"11",
          1618 => x"05",
          1619 => x"3f",
          1620 => x"08",
          1621 => x"a2",
          1622 => x"fe",
          1623 => x"ff",
          1624 => x"a3",
          1625 => x"87",
          1626 => x"2e",
          1627 => x"60",
          1628 => x"60",
          1629 => x"b4",
          1630 => x"11",
          1631 => x"05",
          1632 => x"3f",
          1633 => x"08",
          1634 => x"ee",
          1635 => x"08",
          1636 => x"f4",
          1637 => x"ee",
          1638 => x"52",
          1639 => x"c0",
          1640 => x"79",
          1641 => x"ae",
          1642 => x"38",
          1643 => x"9b",
          1644 => x"fe",
          1645 => x"ff",
          1646 => x"a2",
          1647 => x"87",
          1648 => x"2e",
          1649 => x"60",
          1650 => x"60",
          1651 => x"ff",
          1652 => x"f4",
          1653 => x"ca",
          1654 => x"39",
          1655 => x"51",
          1656 => x"82",
          1657 => x"3f",
          1658 => x"81",
          1659 => x"98",
          1660 => x"51",
          1661 => x"f2",
          1662 => x"f4",
          1663 => x"a2",
          1664 => x"81",
          1665 => x"94",
          1666 => x"80",
          1667 => x"c0",
          1668 => x"f1",
          1669 => x"f4",
          1670 => x"86",
          1671 => x"83",
          1672 => x"94",
          1673 => x"80",
          1674 => x"c0",
          1675 => x"f1",
          1676 => x"3d",
          1677 => x"53",
          1678 => x"51",
          1679 => x"82",
          1680 => x"80",
          1681 => x"38",
          1682 => x"f5",
          1683 => x"b6",
          1684 => x"78",
          1685 => x"ff",
          1686 => x"ff",
          1687 => x"9f",
          1688 => x"87",
          1689 => x"2e",
          1690 => x"63",
          1691 => x"a0",
          1692 => x"3f",
          1693 => x"2d",
          1694 => x"08",
          1695 => x"fa",
          1696 => x"cc",
          1697 => x"f5",
          1698 => x"fa",
          1699 => x"39",
          1700 => x"51",
          1701 => x"de",
          1702 => x"de",
          1703 => x"f4",
          1704 => x"3f",
          1705 => x"ab",
          1706 => x"3f",
          1707 => x"79",
          1708 => x"59",
          1709 => x"f0",
          1710 => x"7d",
          1711 => x"80",
          1712 => x"38",
          1713 => x"84",
          1714 => x"b2",
          1715 => x"cc",
          1716 => x"5c",
          1717 => x"b1",
          1718 => x"24",
          1719 => x"81",
          1720 => x"80",
          1721 => x"83",
          1722 => x"80",
          1723 => x"f6",
          1724 => x"55",
          1725 => x"54",
          1726 => x"f6",
          1727 => x"3d",
          1728 => x"51",
          1729 => x"b8",
          1730 => x"b0",
          1731 => x"ff",
          1732 => x"9c",
          1733 => x"39",
          1734 => x"f6",
          1735 => x"53",
          1736 => x"52",
          1737 => x"b0",
          1738 => x"f0",
          1739 => x"7a",
          1740 => x"81",
          1741 => x"b4",
          1742 => x"05",
          1743 => x"3f",
          1744 => x"58",
          1745 => x"57",
          1746 => x"55",
          1747 => x"a0",
          1748 => x"a0",
          1749 => x"3d",
          1750 => x"51",
          1751 => x"82",
          1752 => x"82",
          1753 => x"09",
          1754 => x"72",
          1755 => x"51",
          1756 => x"80",
          1757 => x"26",
          1758 => x"5a",
          1759 => x"59",
          1760 => x"8d",
          1761 => x"70",
          1762 => x"5d",
          1763 => x"c4",
          1764 => x"32",
          1765 => x"07",
          1766 => x"38",
          1767 => x"09",
          1768 => x"d6",
          1769 => x"b4",
          1770 => x"3f",
          1771 => x"fc",
          1772 => x"0b",
          1773 => x"34",
          1774 => x"8c",
          1775 => x"55",
          1776 => x"52",
          1777 => x"a5",
          1778 => x"cc",
          1779 => x"75",
          1780 => x"87",
          1781 => x"73",
          1782 => x"3f",
          1783 => x"cc",
          1784 => x"0c",
          1785 => x"9c",
          1786 => x"55",
          1787 => x"52",
          1788 => x"f9",
          1789 => x"cc",
          1790 => x"75",
          1791 => x"87",
          1792 => x"73",
          1793 => x"3f",
          1794 => x"cc",
          1795 => x"0c",
          1796 => x"0b",
          1797 => x"84",
          1798 => x"83",
          1799 => x"94",
          1800 => x"a5",
          1801 => x"d4",
          1802 => x"a0",
          1803 => x"d8",
          1804 => x"3f",
          1805 => x"81",
          1806 => x"93",
          1807 => x"f6",
          1808 => x"de",
          1809 => x"51",
          1810 => x"81",
          1811 => x"3f",
          1812 => x"80",
          1813 => x"0d",
          1814 => x"53",
          1815 => x"52",
          1816 => x"82",
          1817 => x"81",
          1818 => x"07",
          1819 => x"52",
          1820 => x"e8",
          1821 => x"87",
          1822 => x"3d",
          1823 => x"3d",
          1824 => x"08",
          1825 => x"73",
          1826 => x"74",
          1827 => x"38",
          1828 => x"70",
          1829 => x"81",
          1830 => x"81",
          1831 => x"39",
          1832 => x"70",
          1833 => x"81",
          1834 => x"81",
          1835 => x"54",
          1836 => x"81",
          1837 => x"06",
          1838 => x"39",
          1839 => x"80",
          1840 => x"54",
          1841 => x"83",
          1842 => x"70",
          1843 => x"38",
          1844 => x"98",
          1845 => x"52",
          1846 => x"52",
          1847 => x"2e",
          1848 => x"54",
          1849 => x"84",
          1850 => x"38",
          1851 => x"52",
          1852 => x"2e",
          1853 => x"83",
          1854 => x"70",
          1855 => x"30",
          1856 => x"76",
          1857 => x"51",
          1858 => x"88",
          1859 => x"70",
          1860 => x"34",
          1861 => x"72",
          1862 => x"87",
          1863 => x"3d",
          1864 => x"3d",
          1865 => x"72",
          1866 => x"91",
          1867 => x"fc",
          1868 => x"51",
          1869 => x"82",
          1870 => x"85",
          1871 => x"83",
          1872 => x"72",
          1873 => x"0c",
          1874 => x"04",
          1875 => x"76",
          1876 => x"ff",
          1877 => x"81",
          1878 => x"26",
          1879 => x"83",
          1880 => x"05",
          1881 => x"70",
          1882 => x"8a",
          1883 => x"33",
          1884 => x"70",
          1885 => x"fe",
          1886 => x"33",
          1887 => x"70",
          1888 => x"f2",
          1889 => x"33",
          1890 => x"70",
          1891 => x"e6",
          1892 => x"22",
          1893 => x"74",
          1894 => x"80",
          1895 => x"13",
          1896 => x"52",
          1897 => x"26",
          1898 => x"81",
          1899 => x"98",
          1900 => x"22",
          1901 => x"bc",
          1902 => x"33",
          1903 => x"b8",
          1904 => x"33",
          1905 => x"b4",
          1906 => x"33",
          1907 => x"b0",
          1908 => x"33",
          1909 => x"ac",
          1910 => x"33",
          1911 => x"a8",
          1912 => x"c0",
          1913 => x"73",
          1914 => x"a0",
          1915 => x"87",
          1916 => x"0c",
          1917 => x"82",
          1918 => x"86",
          1919 => x"f3",
          1920 => x"5b",
          1921 => x"9c",
          1922 => x"0c",
          1923 => x"bc",
          1924 => x"7b",
          1925 => x"98",
          1926 => x"79",
          1927 => x"87",
          1928 => x"08",
          1929 => x"1c",
          1930 => x"98",
          1931 => x"79",
          1932 => x"87",
          1933 => x"08",
          1934 => x"1c",
          1935 => x"98",
          1936 => x"79",
          1937 => x"87",
          1938 => x"08",
          1939 => x"1c",
          1940 => x"98",
          1941 => x"79",
          1942 => x"80",
          1943 => x"83",
          1944 => x"59",
          1945 => x"ff",
          1946 => x"1b",
          1947 => x"1b",
          1948 => x"1b",
          1949 => x"1b",
          1950 => x"1b",
          1951 => x"83",
          1952 => x"52",
          1953 => x"51",
          1954 => x"8f",
          1955 => x"ff",
          1956 => x"8f",
          1957 => x"30",
          1958 => x"51",
          1959 => x"82",
          1960 => x"83",
          1961 => x"fb",
          1962 => x"82",
          1963 => x"70",
          1964 => x"57",
          1965 => x"c0",
          1966 => x"74",
          1967 => x"38",
          1968 => x"94",
          1969 => x"70",
          1970 => x"81",
          1971 => x"52",
          1972 => x"8c",
          1973 => x"2a",
          1974 => x"51",
          1975 => x"38",
          1976 => x"70",
          1977 => x"51",
          1978 => x"8d",
          1979 => x"2a",
          1980 => x"51",
          1981 => x"be",
          1982 => x"ff",
          1983 => x"c0",
          1984 => x"70",
          1985 => x"38",
          1986 => x"90",
          1987 => x"0c",
          1988 => x"cc",
          1989 => x"0d",
          1990 => x"0d",
          1991 => x"33",
          1992 => x"33",
          1993 => x"06",
          1994 => x"87",
          1995 => x"51",
          1996 => x"86",
          1997 => x"94",
          1998 => x"08",
          1999 => x"70",
          2000 => x"54",
          2001 => x"2e",
          2002 => x"91",
          2003 => x"06",
          2004 => x"d7",
          2005 => x"32",
          2006 => x"51",
          2007 => x"2e",
          2008 => x"93",
          2009 => x"06",
          2010 => x"ff",
          2011 => x"81",
          2012 => x"87",
          2013 => x"52",
          2014 => x"86",
          2015 => x"94",
          2016 => x"72",
          2017 => x"0d",
          2018 => x"0d",
          2019 => x"74",
          2020 => x"ff",
          2021 => x"57",
          2022 => x"80",
          2023 => x"81",
          2024 => x"15",
          2025 => x"33",
          2026 => x"06",
          2027 => x"58",
          2028 => x"84",
          2029 => x"2e",
          2030 => x"c0",
          2031 => x"70",
          2032 => x"2a",
          2033 => x"53",
          2034 => x"80",
          2035 => x"71",
          2036 => x"81",
          2037 => x"70",
          2038 => x"81",
          2039 => x"06",
          2040 => x"80",
          2041 => x"71",
          2042 => x"81",
          2043 => x"70",
          2044 => x"74",
          2045 => x"51",
          2046 => x"80",
          2047 => x"2e",
          2048 => x"c0",
          2049 => x"77",
          2050 => x"17",
          2051 => x"81",
          2052 => x"53",
          2053 => x"86",
          2054 => x"87",
          2055 => x"3d",
          2056 => x"3d",
          2057 => x"ec",
          2058 => x"ff",
          2059 => x"87",
          2060 => x"51",
          2061 => x"86",
          2062 => x"94",
          2063 => x"08",
          2064 => x"70",
          2065 => x"51",
          2066 => x"2e",
          2067 => x"81",
          2068 => x"87",
          2069 => x"52",
          2070 => x"86",
          2071 => x"94",
          2072 => x"08",
          2073 => x"06",
          2074 => x"0c",
          2075 => x"0d",
          2076 => x"0d",
          2077 => x"33",
          2078 => x"06",
          2079 => x"c0",
          2080 => x"70",
          2081 => x"38",
          2082 => x"94",
          2083 => x"70",
          2084 => x"81",
          2085 => x"51",
          2086 => x"80",
          2087 => x"72",
          2088 => x"51",
          2089 => x"80",
          2090 => x"2e",
          2091 => x"c0",
          2092 => x"71",
          2093 => x"2b",
          2094 => x"51",
          2095 => x"82",
          2096 => x"84",
          2097 => x"ff",
          2098 => x"c0",
          2099 => x"70",
          2100 => x"06",
          2101 => x"80",
          2102 => x"38",
          2103 => x"a4",
          2104 => x"f0",
          2105 => x"9e",
          2106 => x"85",
          2107 => x"c0",
          2108 => x"82",
          2109 => x"87",
          2110 => x"08",
          2111 => x"0c",
          2112 => x"9c",
          2113 => x"80",
          2114 => x"9e",
          2115 => x"86",
          2116 => x"c0",
          2117 => x"82",
          2118 => x"87",
          2119 => x"08",
          2120 => x"0c",
          2121 => x"b4",
          2122 => x"90",
          2123 => x"9e",
          2124 => x"86",
          2125 => x"c0",
          2126 => x"82",
          2127 => x"87",
          2128 => x"08",
          2129 => x"0c",
          2130 => x"c4",
          2131 => x"a0",
          2132 => x"9e",
          2133 => x"70",
          2134 => x"23",
          2135 => x"84",
          2136 => x"a8",
          2137 => x"9e",
          2138 => x"86",
          2139 => x"c0",
          2140 => x"82",
          2141 => x"81",
          2142 => x"b4",
          2143 => x"87",
          2144 => x"08",
          2145 => x"0a",
          2146 => x"52",
          2147 => x"83",
          2148 => x"71",
          2149 => x"34",
          2150 => x"c0",
          2151 => x"70",
          2152 => x"06",
          2153 => x"70",
          2154 => x"38",
          2155 => x"82",
          2156 => x"80",
          2157 => x"9e",
          2158 => x"90",
          2159 => x"51",
          2160 => x"80",
          2161 => x"81",
          2162 => x"86",
          2163 => x"0b",
          2164 => x"90",
          2165 => x"80",
          2166 => x"52",
          2167 => x"2e",
          2168 => x"52",
          2169 => x"b8",
          2170 => x"87",
          2171 => x"08",
          2172 => x"80",
          2173 => x"52",
          2174 => x"83",
          2175 => x"71",
          2176 => x"34",
          2177 => x"c0",
          2178 => x"70",
          2179 => x"06",
          2180 => x"70",
          2181 => x"38",
          2182 => x"82",
          2183 => x"80",
          2184 => x"9e",
          2185 => x"84",
          2186 => x"51",
          2187 => x"80",
          2188 => x"81",
          2189 => x"86",
          2190 => x"0b",
          2191 => x"90",
          2192 => x"80",
          2193 => x"52",
          2194 => x"2e",
          2195 => x"52",
          2196 => x"bc",
          2197 => x"87",
          2198 => x"08",
          2199 => x"80",
          2200 => x"52",
          2201 => x"83",
          2202 => x"71",
          2203 => x"34",
          2204 => x"c0",
          2205 => x"70",
          2206 => x"06",
          2207 => x"70",
          2208 => x"38",
          2209 => x"82",
          2210 => x"80",
          2211 => x"9e",
          2212 => x"a0",
          2213 => x"52",
          2214 => x"2e",
          2215 => x"52",
          2216 => x"bf",
          2217 => x"9e",
          2218 => x"98",
          2219 => x"8a",
          2220 => x"51",
          2221 => x"c0",
          2222 => x"87",
          2223 => x"08",
          2224 => x"06",
          2225 => x"70",
          2226 => x"38",
          2227 => x"82",
          2228 => x"87",
          2229 => x"08",
          2230 => x"06",
          2231 => x"51",
          2232 => x"82",
          2233 => x"80",
          2234 => x"9e",
          2235 => x"88",
          2236 => x"52",
          2237 => x"83",
          2238 => x"71",
          2239 => x"34",
          2240 => x"90",
          2241 => x"06",
          2242 => x"82",
          2243 => x"83",
          2244 => x"fb",
          2245 => x"f7",
          2246 => x"86",
          2247 => x"b4",
          2248 => x"80",
          2249 => x"81",
          2250 => x"85",
          2251 => x"f7",
          2252 => x"ee",
          2253 => x"b6",
          2254 => x"80",
          2255 => x"82",
          2256 => x"82",
          2257 => x"11",
          2258 => x"f7",
          2259 => x"b6",
          2260 => x"bb",
          2261 => x"80",
          2262 => x"82",
          2263 => x"82",
          2264 => x"11",
          2265 => x"f7",
          2266 => x"9a",
          2267 => x"b8",
          2268 => x"80",
          2269 => x"82",
          2270 => x"82",
          2271 => x"11",
          2272 => x"f7",
          2273 => x"fe",
          2274 => x"b9",
          2275 => x"80",
          2276 => x"82",
          2277 => x"82",
          2278 => x"11",
          2279 => x"f8",
          2280 => x"e2",
          2281 => x"ba",
          2282 => x"80",
          2283 => x"82",
          2284 => x"82",
          2285 => x"11",
          2286 => x"f8",
          2287 => x"c6",
          2288 => x"bf",
          2289 => x"80",
          2290 => x"82",
          2291 => x"52",
          2292 => x"51",
          2293 => x"82",
          2294 => x"54",
          2295 => x"8d",
          2296 => x"c4",
          2297 => x"f8",
          2298 => x"9a",
          2299 => x"c1",
          2300 => x"80",
          2301 => x"82",
          2302 => x"52",
          2303 => x"51",
          2304 => x"82",
          2305 => x"54",
          2306 => x"88",
          2307 => x"ac",
          2308 => x"3f",
          2309 => x"33",
          2310 => x"2e",
          2311 => x"f9",
          2312 => x"fe",
          2313 => x"bc",
          2314 => x"80",
          2315 => x"81",
          2316 => x"83",
          2317 => x"86",
          2318 => x"73",
          2319 => x"38",
          2320 => x"51",
          2321 => x"82",
          2322 => x"54",
          2323 => x"88",
          2324 => x"e4",
          2325 => x"3f",
          2326 => x"51",
          2327 => x"82",
          2328 => x"52",
          2329 => x"51",
          2330 => x"82",
          2331 => x"52",
          2332 => x"51",
          2333 => x"82",
          2334 => x"52",
          2335 => x"51",
          2336 => x"81",
          2337 => x"83",
          2338 => x"86",
          2339 => x"81",
          2340 => x"88",
          2341 => x"86",
          2342 => x"bd",
          2343 => x"75",
          2344 => x"3f",
          2345 => x"08",
          2346 => x"29",
          2347 => x"54",
          2348 => x"cc",
          2349 => x"fb",
          2350 => x"ca",
          2351 => x"bb",
          2352 => x"80",
          2353 => x"82",
          2354 => x"56",
          2355 => x"52",
          2356 => x"99",
          2357 => x"cc",
          2358 => x"c0",
          2359 => x"31",
          2360 => x"87",
          2361 => x"81",
          2362 => x"88",
          2363 => x"86",
          2364 => x"73",
          2365 => x"38",
          2366 => x"08",
          2367 => x"c0",
          2368 => x"a1",
          2369 => x"87",
          2370 => x"84",
          2371 => x"71",
          2372 => x"82",
          2373 => x"52",
          2374 => x"51",
          2375 => x"81",
          2376 => x"81",
          2377 => x"3d",
          2378 => x"3d",
          2379 => x"05",
          2380 => x"52",
          2381 => x"aa",
          2382 => x"29",
          2383 => x"05",
          2384 => x"04",
          2385 => x"51",
          2386 => x"fc",
          2387 => x"39",
          2388 => x"51",
          2389 => x"fc",
          2390 => x"39",
          2391 => x"51",
          2392 => x"fc",
          2393 => x"ba",
          2394 => x"0d",
          2395 => x"80",
          2396 => x"3d",
          2397 => x"96",
          2398 => x"52",
          2399 => x"0c",
          2400 => x"70",
          2401 => x"0c",
          2402 => x"3d",
          2403 => x"3d",
          2404 => x"96",
          2405 => x"82",
          2406 => x"52",
          2407 => x"73",
          2408 => x"86",
          2409 => x"70",
          2410 => x"0c",
          2411 => x"83",
          2412 => x"80",
          2413 => x"96",
          2414 => x"82",
          2415 => x"87",
          2416 => x"0c",
          2417 => x"0d",
          2418 => x"33",
          2419 => x"2e",
          2420 => x"85",
          2421 => x"ed",
          2422 => x"dc",
          2423 => x"80",
          2424 => x"72",
          2425 => x"9e",
          2426 => x"05",
          2427 => x"0c",
          2428 => x"9e",
          2429 => x"71",
          2430 => x"38",
          2431 => x"2d",
          2432 => x"04",
          2433 => x"02",
          2434 => x"82",
          2435 => x"76",
          2436 => x"0c",
          2437 => x"ad",
          2438 => x"9e",
          2439 => x"3d",
          2440 => x"3d",
          2441 => x"73",
          2442 => x"ff",
          2443 => x"71",
          2444 => x"38",
          2445 => x"06",
          2446 => x"54",
          2447 => x"e7",
          2448 => x"0d",
          2449 => x"0d",
          2450 => x"d4",
          2451 => x"9e",
          2452 => x"54",
          2453 => x"81",
          2454 => x"53",
          2455 => x"8e",
          2456 => x"ff",
          2457 => x"14",
          2458 => x"3f",
          2459 => x"82",
          2460 => x"86",
          2461 => x"ec",
          2462 => x"68",
          2463 => x"70",
          2464 => x"33",
          2465 => x"2e",
          2466 => x"75",
          2467 => x"81",
          2468 => x"38",
          2469 => x"70",
          2470 => x"33",
          2471 => x"75",
          2472 => x"81",
          2473 => x"81",
          2474 => x"75",
          2475 => x"81",
          2476 => x"82",
          2477 => x"81",
          2478 => x"56",
          2479 => x"09",
          2480 => x"38",
          2481 => x"71",
          2482 => x"81",
          2483 => x"59",
          2484 => x"9d",
          2485 => x"53",
          2486 => x"95",
          2487 => x"29",
          2488 => x"76",
          2489 => x"79",
          2490 => x"5b",
          2491 => x"e5",
          2492 => x"ec",
          2493 => x"70",
          2494 => x"25",
          2495 => x"32",
          2496 => x"72",
          2497 => x"73",
          2498 => x"58",
          2499 => x"73",
          2500 => x"38",
          2501 => x"79",
          2502 => x"5b",
          2503 => x"75",
          2504 => x"de",
          2505 => x"80",
          2506 => x"89",
          2507 => x"70",
          2508 => x"55",
          2509 => x"cf",
          2510 => x"38",
          2511 => x"24",
          2512 => x"80",
          2513 => x"8e",
          2514 => x"c3",
          2515 => x"73",
          2516 => x"81",
          2517 => x"99",
          2518 => x"c4",
          2519 => x"38",
          2520 => x"73",
          2521 => x"81",
          2522 => x"80",
          2523 => x"38",
          2524 => x"2e",
          2525 => x"f9",
          2526 => x"d8",
          2527 => x"38",
          2528 => x"77",
          2529 => x"08",
          2530 => x"80",
          2531 => x"55",
          2532 => x"8d",
          2533 => x"70",
          2534 => x"51",
          2535 => x"f5",
          2536 => x"2a",
          2537 => x"74",
          2538 => x"53",
          2539 => x"8f",
          2540 => x"fc",
          2541 => x"81",
          2542 => x"80",
          2543 => x"73",
          2544 => x"3f",
          2545 => x"56",
          2546 => x"27",
          2547 => x"a0",
          2548 => x"3f",
          2549 => x"84",
          2550 => x"33",
          2551 => x"93",
          2552 => x"95",
          2553 => x"91",
          2554 => x"8d",
          2555 => x"89",
          2556 => x"fb",
          2557 => x"86",
          2558 => x"2a",
          2559 => x"51",
          2560 => x"2e",
          2561 => x"84",
          2562 => x"86",
          2563 => x"78",
          2564 => x"08",
          2565 => x"32",
          2566 => x"72",
          2567 => x"51",
          2568 => x"74",
          2569 => x"38",
          2570 => x"88",
          2571 => x"7a",
          2572 => x"55",
          2573 => x"3d",
          2574 => x"52",
          2575 => x"d4",
          2576 => x"cc",
          2577 => x"06",
          2578 => x"52",
          2579 => x"3f",
          2580 => x"08",
          2581 => x"27",
          2582 => x"14",
          2583 => x"f8",
          2584 => x"87",
          2585 => x"81",
          2586 => x"b0",
          2587 => x"7d",
          2588 => x"5f",
          2589 => x"75",
          2590 => x"07",
          2591 => x"54",
          2592 => x"26",
          2593 => x"ff",
          2594 => x"84",
          2595 => x"06",
          2596 => x"80",
          2597 => x"96",
          2598 => x"e0",
          2599 => x"73",
          2600 => x"57",
          2601 => x"06",
          2602 => x"54",
          2603 => x"a0",
          2604 => x"2a",
          2605 => x"54",
          2606 => x"38",
          2607 => x"76",
          2608 => x"38",
          2609 => x"fd",
          2610 => x"06",
          2611 => x"38",
          2612 => x"56",
          2613 => x"26",
          2614 => x"3d",
          2615 => x"05",
          2616 => x"ff",
          2617 => x"53",
          2618 => x"d9",
          2619 => x"38",
          2620 => x"56",
          2621 => x"27",
          2622 => x"a0",
          2623 => x"3f",
          2624 => x"3d",
          2625 => x"3d",
          2626 => x"70",
          2627 => x"52",
          2628 => x"73",
          2629 => x"3f",
          2630 => x"04",
          2631 => x"74",
          2632 => x"0c",
          2633 => x"05",
          2634 => x"fa",
          2635 => x"9e",
          2636 => x"80",
          2637 => x"0b",
          2638 => x"0c",
          2639 => x"04",
          2640 => x"82",
          2641 => x"76",
          2642 => x"0c",
          2643 => x"05",
          2644 => x"53",
          2645 => x"72",
          2646 => x"0c",
          2647 => x"04",
          2648 => x"77",
          2649 => x"d8",
          2650 => x"54",
          2651 => x"54",
          2652 => x"80",
          2653 => x"9e",
          2654 => x"71",
          2655 => x"cc",
          2656 => x"06",
          2657 => x"2e",
          2658 => x"72",
          2659 => x"38",
          2660 => x"70",
          2661 => x"25",
          2662 => x"73",
          2663 => x"38",
          2664 => x"86",
          2665 => x"54",
          2666 => x"73",
          2667 => x"ff",
          2668 => x"72",
          2669 => x"74",
          2670 => x"72",
          2671 => x"54",
          2672 => x"81",
          2673 => x"39",
          2674 => x"80",
          2675 => x"51",
          2676 => x"81",
          2677 => x"87",
          2678 => x"3d",
          2679 => x"3d",
          2680 => x"d8",
          2681 => x"9e",
          2682 => x"53",
          2683 => x"fe",
          2684 => x"82",
          2685 => x"84",
          2686 => x"f8",
          2687 => x"7c",
          2688 => x"70",
          2689 => x"75",
          2690 => x"55",
          2691 => x"2e",
          2692 => x"87",
          2693 => x"76",
          2694 => x"73",
          2695 => x"81",
          2696 => x"81",
          2697 => x"77",
          2698 => x"70",
          2699 => x"58",
          2700 => x"09",
          2701 => x"c2",
          2702 => x"81",
          2703 => x"75",
          2704 => x"55",
          2705 => x"e2",
          2706 => x"90",
          2707 => x"f8",
          2708 => x"8f",
          2709 => x"81",
          2710 => x"75",
          2711 => x"55",
          2712 => x"81",
          2713 => x"27",
          2714 => x"d0",
          2715 => x"55",
          2716 => x"73",
          2717 => x"80",
          2718 => x"14",
          2719 => x"72",
          2720 => x"e0",
          2721 => x"80",
          2722 => x"39",
          2723 => x"55",
          2724 => x"80",
          2725 => x"e0",
          2726 => x"38",
          2727 => x"81",
          2728 => x"53",
          2729 => x"81",
          2730 => x"53",
          2731 => x"8e",
          2732 => x"70",
          2733 => x"55",
          2734 => x"27",
          2735 => x"77",
          2736 => x"74",
          2737 => x"76",
          2738 => x"77",
          2739 => x"70",
          2740 => x"55",
          2741 => x"77",
          2742 => x"38",
          2743 => x"74",
          2744 => x"55",
          2745 => x"cc",
          2746 => x"0d",
          2747 => x"0d",
          2748 => x"56",
          2749 => x"0c",
          2750 => x"70",
          2751 => x"73",
          2752 => x"81",
          2753 => x"81",
          2754 => x"ed",
          2755 => x"2e",
          2756 => x"8e",
          2757 => x"08",
          2758 => x"76",
          2759 => x"56",
          2760 => x"b0",
          2761 => x"06",
          2762 => x"75",
          2763 => x"76",
          2764 => x"70",
          2765 => x"73",
          2766 => x"8b",
          2767 => x"73",
          2768 => x"85",
          2769 => x"82",
          2770 => x"76",
          2771 => x"70",
          2772 => x"ac",
          2773 => x"a0",
          2774 => x"fa",
          2775 => x"53",
          2776 => x"57",
          2777 => x"98",
          2778 => x"39",
          2779 => x"80",
          2780 => x"26",
          2781 => x"86",
          2782 => x"80",
          2783 => x"57",
          2784 => x"74",
          2785 => x"38",
          2786 => x"27",
          2787 => x"14",
          2788 => x"06",
          2789 => x"14",
          2790 => x"06",
          2791 => x"74",
          2792 => x"f9",
          2793 => x"ff",
          2794 => x"89",
          2795 => x"38",
          2796 => x"c5",
          2797 => x"29",
          2798 => x"81",
          2799 => x"76",
          2800 => x"56",
          2801 => x"ba",
          2802 => x"2e",
          2803 => x"30",
          2804 => x"0c",
          2805 => x"82",
          2806 => x"8a",
          2807 => x"fd",
          2808 => x"98",
          2809 => x"2c",
          2810 => x"70",
          2811 => x"10",
          2812 => x"2b",
          2813 => x"54",
          2814 => x"0b",
          2815 => x"12",
          2816 => x"71",
          2817 => x"38",
          2818 => x"11",
          2819 => x"84",
          2820 => x"33",
          2821 => x"52",
          2822 => x"2e",
          2823 => x"83",
          2824 => x"72",
          2825 => x"0c",
          2826 => x"04",
          2827 => x"78",
          2828 => x"9f",
          2829 => x"33",
          2830 => x"71",
          2831 => x"38",
          2832 => x"81",
          2833 => x"f2",
          2834 => x"51",
          2835 => x"72",
          2836 => x"52",
          2837 => x"71",
          2838 => x"52",
          2839 => x"51",
          2840 => x"73",
          2841 => x"3d",
          2842 => x"3d",
          2843 => x"84",
          2844 => x"33",
          2845 => x"bb",
          2846 => x"87",
          2847 => x"84",
          2848 => x"cc",
          2849 => x"51",
          2850 => x"58",
          2851 => x"2e",
          2852 => x"51",
          2853 => x"82",
          2854 => x"70",
          2855 => x"86",
          2856 => x"19",
          2857 => x"56",
          2858 => x"3f",
          2859 => x"08",
          2860 => x"87",
          2861 => x"84",
          2862 => x"cc",
          2863 => x"51",
          2864 => x"80",
          2865 => x"75",
          2866 => x"74",
          2867 => x"c9",
          2868 => x"a4",
          2869 => x"55",
          2870 => x"a4",
          2871 => x"ff",
          2872 => x"75",
          2873 => x"80",
          2874 => x"a4",
          2875 => x"2e",
          2876 => x"87",
          2877 => x"75",
          2878 => x"38",
          2879 => x"33",
          2880 => x"38",
          2881 => x"05",
          2882 => x"78",
          2883 => x"80",
          2884 => x"82",
          2885 => x"52",
          2886 => x"8d",
          2887 => x"87",
          2888 => x"80",
          2889 => x"8c",
          2890 => x"fd",
          2891 => x"86",
          2892 => x"54",
          2893 => x"71",
          2894 => x"38",
          2895 => x"d9",
          2896 => x"0c",
          2897 => x"14",
          2898 => x"80",
          2899 => x"80",
          2900 => x"a4",
          2901 => x"a0",
          2902 => x"80",
          2903 => x"71",
          2904 => x"a6",
          2905 => x"a0",
          2906 => x"ad",
          2907 => x"82",
          2908 => x"85",
          2909 => x"dc",
          2910 => x"57",
          2911 => x"87",
          2912 => x"80",
          2913 => x"82",
          2914 => x"80",
          2915 => x"87",
          2916 => x"80",
          2917 => x"3d",
          2918 => x"81",
          2919 => x"82",
          2920 => x"80",
          2921 => x"75",
          2922 => x"8d",
          2923 => x"cc",
          2924 => x"0b",
          2925 => x"08",
          2926 => x"82",
          2927 => x"ff",
          2928 => x"55",
          2929 => x"34",
          2930 => x"52",
          2931 => x"ff",
          2932 => x"f6",
          2933 => x"ff",
          2934 => x"06",
          2935 => x"a6",
          2936 => x"d9",
          2937 => x"3d",
          2938 => x"08",
          2939 => x"70",
          2940 => x"52",
          2941 => x"08",
          2942 => x"9d",
          2943 => x"cc",
          2944 => x"38",
          2945 => x"87",
          2946 => x"55",
          2947 => x"8b",
          2948 => x"56",
          2949 => x"3f",
          2950 => x"08",
          2951 => x"38",
          2952 => x"b7",
          2953 => x"87",
          2954 => x"18",
          2955 => x"0b",
          2956 => x"08",
          2957 => x"82",
          2958 => x"ff",
          2959 => x"55",
          2960 => x"34",
          2961 => x"30",
          2962 => x"9f",
          2963 => x"55",
          2964 => x"85",
          2965 => x"ac",
          2966 => x"a0",
          2967 => x"08",
          2968 => x"e0",
          2969 => x"87",
          2970 => x"2e",
          2971 => x"ff",
          2972 => x"ae",
          2973 => x"2e",
          2974 => x"9b",
          2975 => x"79",
          2976 => x"a3",
          2977 => x"ff",
          2978 => x"ab",
          2979 => x"82",
          2980 => x"74",
          2981 => x"77",
          2982 => x"0c",
          2983 => x"04",
          2984 => x"7c",
          2985 => x"71",
          2986 => x"59",
          2987 => x"a0",
          2988 => x"06",
          2989 => x"33",
          2990 => x"77",
          2991 => x"38",
          2992 => x"5b",
          2993 => x"56",
          2994 => x"a0",
          2995 => x"06",
          2996 => x"75",
          2997 => x"80",
          2998 => x"29",
          2999 => x"05",
          3000 => x"55",
          3001 => x"3f",
          3002 => x"08",
          3003 => x"74",
          3004 => x"b8",
          3005 => x"87",
          3006 => x"c5",
          3007 => x"33",
          3008 => x"2e",
          3009 => x"82",
          3010 => x"b5",
          3011 => x"3f",
          3012 => x"1a",
          3013 => x"fc",
          3014 => x"05",
          3015 => x"3f",
          3016 => x"08",
          3017 => x"38",
          3018 => x"78",
          3019 => x"fd",
          3020 => x"87",
          3021 => x"ff",
          3022 => x"85",
          3023 => x"91",
          3024 => x"70",
          3025 => x"51",
          3026 => x"27",
          3027 => x"80",
          3028 => x"87",
          3029 => x"3d",
          3030 => x"3d",
          3031 => x"08",
          3032 => x"b4",
          3033 => x"5f",
          3034 => x"af",
          3035 => x"87",
          3036 => x"87",
          3037 => x"5b",
          3038 => x"38",
          3039 => x"9c",
          3040 => x"73",
          3041 => x"55",
          3042 => x"81",
          3043 => x"70",
          3044 => x"56",
          3045 => x"81",
          3046 => x"51",
          3047 => x"82",
          3048 => x"82",
          3049 => x"82",
          3050 => x"80",
          3051 => x"38",
          3052 => x"52",
          3053 => x"08",
          3054 => x"dd",
          3055 => x"cc",
          3056 => x"8b",
          3057 => x"80",
          3058 => x"3f",
          3059 => x"82",
          3060 => x"5b",
          3061 => x"08",
          3062 => x"52",
          3063 => x"52",
          3064 => x"9b",
          3065 => x"cc",
          3066 => x"87",
          3067 => x"2e",
          3068 => x"80",
          3069 => x"87",
          3070 => x"ff",
          3071 => x"82",
          3072 => x"55",
          3073 => x"87",
          3074 => x"a9",
          3075 => x"cc",
          3076 => x"70",
          3077 => x"80",
          3078 => x"53",
          3079 => x"06",
          3080 => x"f8",
          3081 => x"1b",
          3082 => x"06",
          3083 => x"7b",
          3084 => x"80",
          3085 => x"2e",
          3086 => x"ff",
          3087 => x"39",
          3088 => x"9c",
          3089 => x"38",
          3090 => x"08",
          3091 => x"38",
          3092 => x"8f",
          3093 => x"99",
          3094 => x"cc",
          3095 => x"70",
          3096 => x"59",
          3097 => x"ee",
          3098 => x"ff",
          3099 => x"e4",
          3100 => x"2b",
          3101 => x"82",
          3102 => x"70",
          3103 => x"97",
          3104 => x"2c",
          3105 => x"29",
          3106 => x"05",
          3107 => x"70",
          3108 => x"51",
          3109 => x"51",
          3110 => x"81",
          3111 => x"2e",
          3112 => x"77",
          3113 => x"38",
          3114 => x"0a",
          3115 => x"0a",
          3116 => x"2c",
          3117 => x"75",
          3118 => x"38",
          3119 => x"52",
          3120 => x"9b",
          3121 => x"cc",
          3122 => x"06",
          3123 => x"2e",
          3124 => x"82",
          3125 => x"81",
          3126 => x"74",
          3127 => x"29",
          3128 => x"05",
          3129 => x"70",
          3130 => x"56",
          3131 => x"95",
          3132 => x"76",
          3133 => x"77",
          3134 => x"3f",
          3135 => x"08",
          3136 => x"54",
          3137 => x"d3",
          3138 => x"75",
          3139 => x"ca",
          3140 => x"55",
          3141 => x"e4",
          3142 => x"2b",
          3143 => x"82",
          3144 => x"70",
          3145 => x"98",
          3146 => x"11",
          3147 => x"81",
          3148 => x"33",
          3149 => x"51",
          3150 => x"55",
          3151 => x"09",
          3152 => x"92",
          3153 => x"dc",
          3154 => x"0c",
          3155 => x"9e",
          3156 => x"0b",
          3157 => x"34",
          3158 => x"82",
          3159 => x"75",
          3160 => x"34",
          3161 => x"34",
          3162 => x"7e",
          3163 => x"26",
          3164 => x"73",
          3165 => x"e9",
          3166 => x"73",
          3167 => x"9e",
          3168 => x"73",
          3169 => x"cb",
          3170 => x"e8",
          3171 => x"75",
          3172 => x"74",
          3173 => x"98",
          3174 => x"73",
          3175 => x"38",
          3176 => x"73",
          3177 => x"34",
          3178 => x"0a",
          3179 => x"0a",
          3180 => x"2c",
          3181 => x"33",
          3182 => x"df",
          3183 => x"ec",
          3184 => x"56",
          3185 => x"9e",
          3186 => x"1a",
          3187 => x"33",
          3188 => x"9e",
          3189 => x"73",
          3190 => x"38",
          3191 => x"73",
          3192 => x"34",
          3193 => x"33",
          3194 => x"0a",
          3195 => x"0a",
          3196 => x"2c",
          3197 => x"33",
          3198 => x"56",
          3199 => x"a2",
          3200 => x"70",
          3201 => x"e7",
          3202 => x"81",
          3203 => x"81",
          3204 => x"70",
          3205 => x"9e",
          3206 => x"51",
          3207 => x"24",
          3208 => x"9e",
          3209 => x"98",
          3210 => x"2c",
          3211 => x"33",
          3212 => x"56",
          3213 => x"fc",
          3214 => x"51",
          3215 => x"74",
          3216 => x"29",
          3217 => x"05",
          3218 => x"82",
          3219 => x"56",
          3220 => x"75",
          3221 => x"fb",
          3222 => x"7a",
          3223 => x"81",
          3224 => x"9e",
          3225 => x"52",
          3226 => x"51",
          3227 => x"81",
          3228 => x"9e",
          3229 => x"81",
          3230 => x"55",
          3231 => x"fb",
          3232 => x"9e",
          3233 => x"05",
          3234 => x"9e",
          3235 => x"15",
          3236 => x"9e",
          3237 => x"51",
          3238 => x"82",
          3239 => x"70",
          3240 => x"98",
          3241 => x"e8",
          3242 => x"56",
          3243 => x"25",
          3244 => x"1a",
          3245 => x"33",
          3246 => x"33",
          3247 => x"3f",
          3248 => x"0a",
          3249 => x"0a",
          3250 => x"2c",
          3251 => x"33",
          3252 => x"75",
          3253 => x"38",
          3254 => x"e9",
          3255 => x"ec",
          3256 => x"2b",
          3257 => x"82",
          3258 => x"57",
          3259 => x"74",
          3260 => x"df",
          3261 => x"e5",
          3262 => x"81",
          3263 => x"81",
          3264 => x"70",
          3265 => x"9e",
          3266 => x"51",
          3267 => x"25",
          3268 => x"bf",
          3269 => x"e8",
          3270 => x"54",
          3271 => x"8a",
          3272 => x"3f",
          3273 => x"52",
          3274 => x"f4",
          3275 => x"cc",
          3276 => x"06",
          3277 => x"38",
          3278 => x"33",
          3279 => x"2e",
          3280 => x"53",
          3281 => x"51",
          3282 => x"84",
          3283 => x"34",
          3284 => x"9e",
          3285 => x"0b",
          3286 => x"34",
          3287 => x"cc",
          3288 => x"0d",
          3289 => x"ec",
          3290 => x"80",
          3291 => x"38",
          3292 => x"d1",
          3293 => x"ec",
          3294 => x"54",
          3295 => x"ec",
          3296 => x"ff",
          3297 => x"39",
          3298 => x"33",
          3299 => x"33",
          3300 => x"75",
          3301 => x"38",
          3302 => x"73",
          3303 => x"34",
          3304 => x"70",
          3305 => x"81",
          3306 => x"51",
          3307 => x"25",
          3308 => x"1a",
          3309 => x"33",
          3310 => x"33",
          3311 => x"3f",
          3312 => x"0a",
          3313 => x"0a",
          3314 => x"2c",
          3315 => x"33",
          3316 => x"75",
          3317 => x"38",
          3318 => x"e9",
          3319 => x"ec",
          3320 => x"2b",
          3321 => x"82",
          3322 => x"57",
          3323 => x"74",
          3324 => x"df",
          3325 => x"e3",
          3326 => x"81",
          3327 => x"81",
          3328 => x"70",
          3329 => x"9e",
          3330 => x"51",
          3331 => x"25",
          3332 => x"bf",
          3333 => x"ec",
          3334 => x"ff",
          3335 => x"e8",
          3336 => x"54",
          3337 => x"f8",
          3338 => x"14",
          3339 => x"9e",
          3340 => x"1a",
          3341 => x"54",
          3342 => x"82",
          3343 => x"70",
          3344 => x"82",
          3345 => x"58",
          3346 => x"75",
          3347 => x"f8",
          3348 => x"9e",
          3349 => x"52",
          3350 => x"51",
          3351 => x"80",
          3352 => x"ec",
          3353 => x"82",
          3354 => x"f7",
          3355 => x"b0",
          3356 => x"98",
          3357 => x"80",
          3358 => x"74",
          3359 => x"b9",
          3360 => x"cc",
          3361 => x"e8",
          3362 => x"cc",
          3363 => x"06",
          3364 => x"74",
          3365 => x"ff",
          3366 => x"93",
          3367 => x"39",
          3368 => x"82",
          3369 => x"fc",
          3370 => x"54",
          3371 => x"a7",
          3372 => x"ff",
          3373 => x"82",
          3374 => x"82",
          3375 => x"82",
          3376 => x"81",
          3377 => x"05",
          3378 => x"79",
          3379 => x"c9",
          3380 => x"54",
          3381 => x"73",
          3382 => x"80",
          3383 => x"38",
          3384 => x"a9",
          3385 => x"39",
          3386 => x"09",
          3387 => x"38",
          3388 => x"08",
          3389 => x"2e",
          3390 => x"51",
          3391 => x"3f",
          3392 => x"08",
          3393 => x"34",
          3394 => x"08",
          3395 => x"81",
          3396 => x"52",
          3397 => x"ab",
          3398 => x"c3",
          3399 => x"29",
          3400 => x"05",
          3401 => x"54",
          3402 => x"ab",
          3403 => x"ff",
          3404 => x"82",
          3405 => x"82",
          3406 => x"82",
          3407 => x"81",
          3408 => x"05",
          3409 => x"79",
          3410 => x"cd",
          3411 => x"54",
          3412 => x"06",
          3413 => x"74",
          3414 => x"34",
          3415 => x"82",
          3416 => x"82",
          3417 => x"52",
          3418 => x"c0",
          3419 => x"39",
          3420 => x"33",
          3421 => x"06",
          3422 => x"33",
          3423 => x"74",
          3424 => x"cf",
          3425 => x"54",
          3426 => x"ec",
          3427 => x"70",
          3428 => x"e0",
          3429 => x"bb",
          3430 => x"ec",
          3431 => x"80",
          3432 => x"38",
          3433 => x"9d",
          3434 => x"ec",
          3435 => x"54",
          3436 => x"ec",
          3437 => x"39",
          3438 => x"77",
          3439 => x"9f",
          3440 => x"2c",
          3441 => x"73",
          3442 => x"2c",
          3443 => x"74",
          3444 => x"31",
          3445 => x"54",
          3446 => x"91",
          3447 => x"cc",
          3448 => x"74",
          3449 => x"cc",
          3450 => x"0d",
          3451 => x"0d",
          3452 => x"55",
          3453 => x"80",
          3454 => x"76",
          3455 => x"3f",
          3456 => x"08",
          3457 => x"53",
          3458 => x"8d",
          3459 => x"80",
          3460 => x"82",
          3461 => x"31",
          3462 => x"72",
          3463 => x"cb",
          3464 => x"72",
          3465 => x"c3",
          3466 => x"75",
          3467 => x"72",
          3468 => x"2b",
          3469 => x"53",
          3470 => x"76",
          3471 => x"73",
          3472 => x"2a",
          3473 => x"77",
          3474 => x"31",
          3475 => x"2c",
          3476 => x"7b",
          3477 => x"71",
          3478 => x"5a",
          3479 => x"51",
          3480 => x"72",
          3481 => x"10",
          3482 => x"71",
          3483 => x"0c",
          3484 => x"04",
          3485 => x"75",
          3486 => x"80",
          3487 => x"70",
          3488 => x"25",
          3489 => x"90",
          3490 => x"71",
          3491 => x"74",
          3492 => x"06",
          3493 => x"80",
          3494 => x"88",
          3495 => x"71",
          3496 => x"73",
          3497 => x"f0",
          3498 => x"70",
          3499 => x"2b",
          3500 => x"7b",
          3501 => x"52",
          3502 => x"8c",
          3503 => x"70",
          3504 => x"82",
          3505 => x"71",
          3506 => x"2a",
          3507 => x"81",
          3508 => x"82",
          3509 => x"75",
          3510 => x"87",
          3511 => x"52",
          3512 => x"51",
          3513 => x"52",
          3514 => x"53",
          3515 => x"52",
          3516 => x"04",
          3517 => x"75",
          3518 => x"71",
          3519 => x"fd",
          3520 => x"87",
          3521 => x"29",
          3522 => x"82",
          3523 => x"53",
          3524 => x"04",
          3525 => x"78",
          3526 => x"a0",
          3527 => x"2e",
          3528 => x"51",
          3529 => x"82",
          3530 => x"52",
          3531 => x"74",
          3532 => x"38",
          3533 => x"bc",
          3534 => x"87",
          3535 => x"53",
          3536 => x"9f",
          3537 => x"38",
          3538 => x"9f",
          3539 => x"38",
          3540 => x"71",
          3541 => x"31",
          3542 => x"58",
          3543 => x"80",
          3544 => x"2e",
          3545 => x"10",
          3546 => x"07",
          3547 => x"07",
          3548 => x"ff",
          3549 => x"70",
          3550 => x"72",
          3551 => x"31",
          3552 => x"56",
          3553 => x"54",
          3554 => x"da",
          3555 => x"71",
          3556 => x"0c",
          3557 => x"04",
          3558 => x"83",
          3559 => x"82",
          3560 => x"84",
          3561 => x"87",
          3562 => x"80",
          3563 => x"83",
          3564 => x"ff",
          3565 => x"82",
          3566 => x"54",
          3567 => x"74",
          3568 => x"76",
          3569 => x"82",
          3570 => x"54",
          3571 => x"34",
          3572 => x"34",
          3573 => x"08",
          3574 => x"15",
          3575 => x"15",
          3576 => x"c4",
          3577 => x"c0",
          3578 => x"fe",
          3579 => x"70",
          3580 => x"06",
          3581 => x"58",
          3582 => x"74",
          3583 => x"73",
          3584 => x"82",
          3585 => x"70",
          3586 => x"87",
          3587 => x"f8",
          3588 => x"55",
          3589 => x"34",
          3590 => x"34",
          3591 => x"04",
          3592 => x"73",
          3593 => x"84",
          3594 => x"38",
          3595 => x"2a",
          3596 => x"83",
          3597 => x"51",
          3598 => x"82",
          3599 => x"83",
          3600 => x"f9",
          3601 => x"a6",
          3602 => x"84",
          3603 => x"22",
          3604 => x"87",
          3605 => x"83",
          3606 => x"74",
          3607 => x"11",
          3608 => x"12",
          3609 => x"2b",
          3610 => x"05",
          3611 => x"71",
          3612 => x"06",
          3613 => x"2a",
          3614 => x"59",
          3615 => x"57",
          3616 => x"71",
          3617 => x"81",
          3618 => x"87",
          3619 => x"75",
          3620 => x"54",
          3621 => x"34",
          3622 => x"34",
          3623 => x"08",
          3624 => x"33",
          3625 => x"71",
          3626 => x"70",
          3627 => x"ff",
          3628 => x"52",
          3629 => x"05",
          3630 => x"ff",
          3631 => x"2a",
          3632 => x"71",
          3633 => x"72",
          3634 => x"53",
          3635 => x"34",
          3636 => x"08",
          3637 => x"76",
          3638 => x"17",
          3639 => x"0d",
          3640 => x"0d",
          3641 => x"08",
          3642 => x"9e",
          3643 => x"83",
          3644 => x"86",
          3645 => x"12",
          3646 => x"2b",
          3647 => x"07",
          3648 => x"52",
          3649 => x"05",
          3650 => x"85",
          3651 => x"88",
          3652 => x"88",
          3653 => x"56",
          3654 => x"13",
          3655 => x"13",
          3656 => x"c4",
          3657 => x"84",
          3658 => x"12",
          3659 => x"2b",
          3660 => x"07",
          3661 => x"52",
          3662 => x"12",
          3663 => x"33",
          3664 => x"07",
          3665 => x"54",
          3666 => x"70",
          3667 => x"73",
          3668 => x"82",
          3669 => x"13",
          3670 => x"12",
          3671 => x"2b",
          3672 => x"ff",
          3673 => x"88",
          3674 => x"53",
          3675 => x"73",
          3676 => x"14",
          3677 => x"0d",
          3678 => x"0d",
          3679 => x"22",
          3680 => x"08",
          3681 => x"71",
          3682 => x"81",
          3683 => x"88",
          3684 => x"88",
          3685 => x"33",
          3686 => x"71",
          3687 => x"90",
          3688 => x"5f",
          3689 => x"5a",
          3690 => x"54",
          3691 => x"80",
          3692 => x"51",
          3693 => x"82",
          3694 => x"70",
          3695 => x"81",
          3696 => x"8b",
          3697 => x"2b",
          3698 => x"70",
          3699 => x"33",
          3700 => x"07",
          3701 => x"8f",
          3702 => x"51",
          3703 => x"53",
          3704 => x"72",
          3705 => x"2a",
          3706 => x"82",
          3707 => x"83",
          3708 => x"87",
          3709 => x"16",
          3710 => x"12",
          3711 => x"2b",
          3712 => x"07",
          3713 => x"55",
          3714 => x"33",
          3715 => x"71",
          3716 => x"70",
          3717 => x"06",
          3718 => x"57",
          3719 => x"52",
          3720 => x"71",
          3721 => x"88",
          3722 => x"fb",
          3723 => x"87",
          3724 => x"84",
          3725 => x"22",
          3726 => x"72",
          3727 => x"33",
          3728 => x"71",
          3729 => x"83",
          3730 => x"5b",
          3731 => x"52",
          3732 => x"33",
          3733 => x"71",
          3734 => x"02",
          3735 => x"05",
          3736 => x"70",
          3737 => x"51",
          3738 => x"71",
          3739 => x"81",
          3740 => x"87",
          3741 => x"15",
          3742 => x"12",
          3743 => x"2b",
          3744 => x"07",
          3745 => x"52",
          3746 => x"12",
          3747 => x"33",
          3748 => x"07",
          3749 => x"54",
          3750 => x"70",
          3751 => x"72",
          3752 => x"82",
          3753 => x"14",
          3754 => x"83",
          3755 => x"88",
          3756 => x"87",
          3757 => x"54",
          3758 => x"04",
          3759 => x"7b",
          3760 => x"08",
          3761 => x"70",
          3762 => x"06",
          3763 => x"53",
          3764 => x"82",
          3765 => x"76",
          3766 => x"11",
          3767 => x"83",
          3768 => x"8b",
          3769 => x"2b",
          3770 => x"70",
          3771 => x"33",
          3772 => x"71",
          3773 => x"53",
          3774 => x"53",
          3775 => x"59",
          3776 => x"25",
          3777 => x"80",
          3778 => x"51",
          3779 => x"81",
          3780 => x"14",
          3781 => x"33",
          3782 => x"71",
          3783 => x"76",
          3784 => x"2a",
          3785 => x"58",
          3786 => x"14",
          3787 => x"ff",
          3788 => x"87",
          3789 => x"87",
          3790 => x"19",
          3791 => x"85",
          3792 => x"88",
          3793 => x"88",
          3794 => x"5b",
          3795 => x"84",
          3796 => x"85",
          3797 => x"87",
          3798 => x"53",
          3799 => x"14",
          3800 => x"87",
          3801 => x"87",
          3802 => x"76",
          3803 => x"75",
          3804 => x"82",
          3805 => x"18",
          3806 => x"12",
          3807 => x"2b",
          3808 => x"80",
          3809 => x"88",
          3810 => x"55",
          3811 => x"74",
          3812 => x"15",
          3813 => x"0d",
          3814 => x"0d",
          3815 => x"87",
          3816 => x"38",
          3817 => x"71",
          3818 => x"38",
          3819 => x"8c",
          3820 => x"0d",
          3821 => x"0d",
          3822 => x"58",
          3823 => x"82",
          3824 => x"83",
          3825 => x"82",
          3826 => x"84",
          3827 => x"12",
          3828 => x"2b",
          3829 => x"59",
          3830 => x"81",
          3831 => x"75",
          3832 => x"cb",
          3833 => x"29",
          3834 => x"81",
          3835 => x"88",
          3836 => x"81",
          3837 => x"79",
          3838 => x"ff",
          3839 => x"7f",
          3840 => x"51",
          3841 => x"77",
          3842 => x"38",
          3843 => x"85",
          3844 => x"5a",
          3845 => x"33",
          3846 => x"71",
          3847 => x"57",
          3848 => x"38",
          3849 => x"ff",
          3850 => x"7a",
          3851 => x"80",
          3852 => x"82",
          3853 => x"11",
          3854 => x"12",
          3855 => x"2b",
          3856 => x"ff",
          3857 => x"52",
          3858 => x"55",
          3859 => x"83",
          3860 => x"80",
          3861 => x"26",
          3862 => x"74",
          3863 => x"2e",
          3864 => x"77",
          3865 => x"81",
          3866 => x"75",
          3867 => x"3f",
          3868 => x"82",
          3869 => x"79",
          3870 => x"f7",
          3871 => x"87",
          3872 => x"1c",
          3873 => x"87",
          3874 => x"8b",
          3875 => x"2b",
          3876 => x"5e",
          3877 => x"7a",
          3878 => x"ff",
          3879 => x"88",
          3880 => x"56",
          3881 => x"15",
          3882 => x"ff",
          3883 => x"85",
          3884 => x"87",
          3885 => x"83",
          3886 => x"72",
          3887 => x"33",
          3888 => x"71",
          3889 => x"70",
          3890 => x"5b",
          3891 => x"56",
          3892 => x"19",
          3893 => x"19",
          3894 => x"c4",
          3895 => x"84",
          3896 => x"12",
          3897 => x"2b",
          3898 => x"07",
          3899 => x"55",
          3900 => x"78",
          3901 => x"76",
          3902 => x"82",
          3903 => x"70",
          3904 => x"84",
          3905 => x"12",
          3906 => x"2b",
          3907 => x"2a",
          3908 => x"52",
          3909 => x"84",
          3910 => x"85",
          3911 => x"87",
          3912 => x"84",
          3913 => x"82",
          3914 => x"8d",
          3915 => x"fe",
          3916 => x"52",
          3917 => x"08",
          3918 => x"dc",
          3919 => x"71",
          3920 => x"38",
          3921 => x"ed",
          3922 => x"cc",
          3923 => x"82",
          3924 => x"84",
          3925 => x"ff",
          3926 => x"8f",
          3927 => x"81",
          3928 => x"26",
          3929 => x"87",
          3930 => x"52",
          3931 => x"cc",
          3932 => x"0d",
          3933 => x"0d",
          3934 => x"33",
          3935 => x"9f",
          3936 => x"53",
          3937 => x"81",
          3938 => x"38",
          3939 => x"87",
          3940 => x"11",
          3941 => x"54",
          3942 => x"84",
          3943 => x"54",
          3944 => x"87",
          3945 => x"11",
          3946 => x"0c",
          3947 => x"c0",
          3948 => x"70",
          3949 => x"70",
          3950 => x"51",
          3951 => x"8a",
          3952 => x"98",
          3953 => x"70",
          3954 => x"08",
          3955 => x"06",
          3956 => x"38",
          3957 => x"8c",
          3958 => x"80",
          3959 => x"71",
          3960 => x"14",
          3961 => x"c8",
          3962 => x"70",
          3963 => x"0c",
          3964 => x"04",
          3965 => x"60",
          3966 => x"8c",
          3967 => x"33",
          3968 => x"5b",
          3969 => x"5a",
          3970 => x"82",
          3971 => x"81",
          3972 => x"52",
          3973 => x"38",
          3974 => x"84",
          3975 => x"92",
          3976 => x"c0",
          3977 => x"87",
          3978 => x"13",
          3979 => x"57",
          3980 => x"0b",
          3981 => x"8c",
          3982 => x"0c",
          3983 => x"75",
          3984 => x"2a",
          3985 => x"51",
          3986 => x"80",
          3987 => x"7b",
          3988 => x"7b",
          3989 => x"5d",
          3990 => x"59",
          3991 => x"06",
          3992 => x"73",
          3993 => x"81",
          3994 => x"ff",
          3995 => x"72",
          3996 => x"38",
          3997 => x"8c",
          3998 => x"c3",
          3999 => x"98",
          4000 => x"71",
          4001 => x"38",
          4002 => x"2e",
          4003 => x"76",
          4004 => x"92",
          4005 => x"72",
          4006 => x"06",
          4007 => x"f7",
          4008 => x"5a",
          4009 => x"80",
          4010 => x"70",
          4011 => x"5a",
          4012 => x"80",
          4013 => x"73",
          4014 => x"06",
          4015 => x"38",
          4016 => x"fe",
          4017 => x"fc",
          4018 => x"52",
          4019 => x"83",
          4020 => x"71",
          4021 => x"87",
          4022 => x"3d",
          4023 => x"3d",
          4024 => x"64",
          4025 => x"bf",
          4026 => x"40",
          4027 => x"59",
          4028 => x"58",
          4029 => x"82",
          4030 => x"81",
          4031 => x"52",
          4032 => x"09",
          4033 => x"b1",
          4034 => x"84",
          4035 => x"92",
          4036 => x"c0",
          4037 => x"87",
          4038 => x"13",
          4039 => x"56",
          4040 => x"87",
          4041 => x"0c",
          4042 => x"82",
          4043 => x"58",
          4044 => x"84",
          4045 => x"06",
          4046 => x"71",
          4047 => x"38",
          4048 => x"05",
          4049 => x"0c",
          4050 => x"73",
          4051 => x"81",
          4052 => x"71",
          4053 => x"38",
          4054 => x"8c",
          4055 => x"d0",
          4056 => x"98",
          4057 => x"71",
          4058 => x"38",
          4059 => x"2e",
          4060 => x"76",
          4061 => x"92",
          4062 => x"72",
          4063 => x"06",
          4064 => x"f7",
          4065 => x"59",
          4066 => x"1a",
          4067 => x"06",
          4068 => x"59",
          4069 => x"80",
          4070 => x"73",
          4071 => x"06",
          4072 => x"38",
          4073 => x"fe",
          4074 => x"fc",
          4075 => x"52",
          4076 => x"83",
          4077 => x"71",
          4078 => x"87",
          4079 => x"3d",
          4080 => x"3d",
          4081 => x"84",
          4082 => x"33",
          4083 => x"a7",
          4084 => x"54",
          4085 => x"fa",
          4086 => x"87",
          4087 => x"06",
          4088 => x"72",
          4089 => x"85",
          4090 => x"98",
          4091 => x"56",
          4092 => x"80",
          4093 => x"76",
          4094 => x"74",
          4095 => x"c0",
          4096 => x"54",
          4097 => x"2e",
          4098 => x"d4",
          4099 => x"2e",
          4100 => x"80",
          4101 => x"08",
          4102 => x"70",
          4103 => x"51",
          4104 => x"2e",
          4105 => x"c0",
          4106 => x"52",
          4107 => x"87",
          4108 => x"08",
          4109 => x"38",
          4110 => x"87",
          4111 => x"14",
          4112 => x"70",
          4113 => x"52",
          4114 => x"96",
          4115 => x"92",
          4116 => x"0a",
          4117 => x"39",
          4118 => x"0c",
          4119 => x"39",
          4120 => x"54",
          4121 => x"cc",
          4122 => x"0d",
          4123 => x"0d",
          4124 => x"33",
          4125 => x"88",
          4126 => x"87",
          4127 => x"51",
          4128 => x"04",
          4129 => x"75",
          4130 => x"82",
          4131 => x"90",
          4132 => x"2b",
          4133 => x"33",
          4134 => x"88",
          4135 => x"71",
          4136 => x"cc",
          4137 => x"54",
          4138 => x"85",
          4139 => x"ff",
          4140 => x"02",
          4141 => x"05",
          4142 => x"70",
          4143 => x"05",
          4144 => x"88",
          4145 => x"72",
          4146 => x"0d",
          4147 => x"0d",
          4148 => x"52",
          4149 => x"81",
          4150 => x"70",
          4151 => x"70",
          4152 => x"05",
          4153 => x"88",
          4154 => x"72",
          4155 => x"54",
          4156 => x"2a",
          4157 => x"34",
          4158 => x"04",
          4159 => x"76",
          4160 => x"54",
          4161 => x"2e",
          4162 => x"70",
          4163 => x"33",
          4164 => x"05",
          4165 => x"11",
          4166 => x"84",
          4167 => x"fe",
          4168 => x"77",
          4169 => x"53",
          4170 => x"81",
          4171 => x"ff",
          4172 => x"f4",
          4173 => x"0d",
          4174 => x"0d",
          4175 => x"56",
          4176 => x"70",
          4177 => x"33",
          4178 => x"05",
          4179 => x"71",
          4180 => x"56",
          4181 => x"72",
          4182 => x"38",
          4183 => x"e2",
          4184 => x"87",
          4185 => x"3d",
          4186 => x"3d",
          4187 => x"54",
          4188 => x"71",
          4189 => x"38",
          4190 => x"70",
          4191 => x"f3",
          4192 => x"82",
          4193 => x"84",
          4194 => x"80",
          4195 => x"cc",
          4196 => x"0b",
          4197 => x"0c",
          4198 => x"0d",
          4199 => x"0b",
          4200 => x"56",
          4201 => x"2e",
          4202 => x"81",
          4203 => x"08",
          4204 => x"70",
          4205 => x"33",
          4206 => x"a2",
          4207 => x"cc",
          4208 => x"09",
          4209 => x"38",
          4210 => x"08",
          4211 => x"b0",
          4212 => x"a4",
          4213 => x"9c",
          4214 => x"56",
          4215 => x"27",
          4216 => x"16",
          4217 => x"82",
          4218 => x"06",
          4219 => x"54",
          4220 => x"78",
          4221 => x"33",
          4222 => x"3f",
          4223 => x"5a",
          4224 => x"cc",
          4225 => x"0d",
          4226 => x"0d",
          4227 => x"56",
          4228 => x"b0",
          4229 => x"af",
          4230 => x"fe",
          4231 => x"87",
          4232 => x"82",
          4233 => x"9f",
          4234 => x"74",
          4235 => x"52",
          4236 => x"51",
          4237 => x"82",
          4238 => x"80",
          4239 => x"ff",
          4240 => x"74",
          4241 => x"76",
          4242 => x"0c",
          4243 => x"04",
          4244 => x"7a",
          4245 => x"fe",
          4246 => x"87",
          4247 => x"82",
          4248 => x"81",
          4249 => x"33",
          4250 => x"2e",
          4251 => x"80",
          4252 => x"17",
          4253 => x"81",
          4254 => x"06",
          4255 => x"84",
          4256 => x"87",
          4257 => x"b4",
          4258 => x"56",
          4259 => x"82",
          4260 => x"84",
          4261 => x"fc",
          4262 => x"8b",
          4263 => x"52",
          4264 => x"a9",
          4265 => x"85",
          4266 => x"84",
          4267 => x"fc",
          4268 => x"17",
          4269 => x"9c",
          4270 => x"91",
          4271 => x"08",
          4272 => x"17",
          4273 => x"3f",
          4274 => x"81",
          4275 => x"19",
          4276 => x"53",
          4277 => x"17",
          4278 => x"82",
          4279 => x"18",
          4280 => x"80",
          4281 => x"33",
          4282 => x"3f",
          4283 => x"08",
          4284 => x"38",
          4285 => x"82",
          4286 => x"8a",
          4287 => x"fb",
          4288 => x"fe",
          4289 => x"08",
          4290 => x"56",
          4291 => x"74",
          4292 => x"38",
          4293 => x"75",
          4294 => x"16",
          4295 => x"53",
          4296 => x"cc",
          4297 => x"0d",
          4298 => x"0d",
          4299 => x"08",
          4300 => x"81",
          4301 => x"df",
          4302 => x"15",
          4303 => x"d7",
          4304 => x"33",
          4305 => x"82",
          4306 => x"38",
          4307 => x"89",
          4308 => x"2e",
          4309 => x"bf",
          4310 => x"2e",
          4311 => x"81",
          4312 => x"81",
          4313 => x"89",
          4314 => x"08",
          4315 => x"52",
          4316 => x"3f",
          4317 => x"08",
          4318 => x"74",
          4319 => x"14",
          4320 => x"81",
          4321 => x"2a",
          4322 => x"05",
          4323 => x"57",
          4324 => x"f5",
          4325 => x"cc",
          4326 => x"38",
          4327 => x"06",
          4328 => x"33",
          4329 => x"78",
          4330 => x"06",
          4331 => x"5c",
          4332 => x"53",
          4333 => x"38",
          4334 => x"06",
          4335 => x"39",
          4336 => x"a4",
          4337 => x"52",
          4338 => x"bd",
          4339 => x"cc",
          4340 => x"38",
          4341 => x"fe",
          4342 => x"b4",
          4343 => x"8d",
          4344 => x"cc",
          4345 => x"ff",
          4346 => x"39",
          4347 => x"a4",
          4348 => x"52",
          4349 => x"91",
          4350 => x"cc",
          4351 => x"76",
          4352 => x"fc",
          4353 => x"b4",
          4354 => x"f8",
          4355 => x"cc",
          4356 => x"06",
          4357 => x"81",
          4358 => x"87",
          4359 => x"3d",
          4360 => x"3d",
          4361 => x"7e",
          4362 => x"82",
          4363 => x"27",
          4364 => x"76",
          4365 => x"27",
          4366 => x"75",
          4367 => x"79",
          4368 => x"38",
          4369 => x"89",
          4370 => x"2e",
          4371 => x"80",
          4372 => x"2e",
          4373 => x"81",
          4374 => x"81",
          4375 => x"89",
          4376 => x"08",
          4377 => x"52",
          4378 => x"3f",
          4379 => x"08",
          4380 => x"cc",
          4381 => x"38",
          4382 => x"06",
          4383 => x"81",
          4384 => x"06",
          4385 => x"77",
          4386 => x"2e",
          4387 => x"84",
          4388 => x"06",
          4389 => x"06",
          4390 => x"53",
          4391 => x"81",
          4392 => x"34",
          4393 => x"a4",
          4394 => x"52",
          4395 => x"d9",
          4396 => x"cc",
          4397 => x"87",
          4398 => x"94",
          4399 => x"ff",
          4400 => x"05",
          4401 => x"54",
          4402 => x"38",
          4403 => x"74",
          4404 => x"06",
          4405 => x"07",
          4406 => x"74",
          4407 => x"39",
          4408 => x"a4",
          4409 => x"52",
          4410 => x"9d",
          4411 => x"cc",
          4412 => x"87",
          4413 => x"d8",
          4414 => x"ff",
          4415 => x"76",
          4416 => x"06",
          4417 => x"05",
          4418 => x"3f",
          4419 => x"87",
          4420 => x"08",
          4421 => x"51",
          4422 => x"82",
          4423 => x"59",
          4424 => x"08",
          4425 => x"f0",
          4426 => x"82",
          4427 => x"06",
          4428 => x"05",
          4429 => x"54",
          4430 => x"3f",
          4431 => x"08",
          4432 => x"74",
          4433 => x"51",
          4434 => x"81",
          4435 => x"34",
          4436 => x"cc",
          4437 => x"0d",
          4438 => x"0d",
          4439 => x"72",
          4440 => x"56",
          4441 => x"27",
          4442 => x"98",
          4443 => x"9d",
          4444 => x"2e",
          4445 => x"53",
          4446 => x"51",
          4447 => x"82",
          4448 => x"54",
          4449 => x"08",
          4450 => x"93",
          4451 => x"80",
          4452 => x"54",
          4453 => x"82",
          4454 => x"54",
          4455 => x"74",
          4456 => x"fb",
          4457 => x"87",
          4458 => x"82",
          4459 => x"80",
          4460 => x"38",
          4461 => x"08",
          4462 => x"38",
          4463 => x"08",
          4464 => x"38",
          4465 => x"52",
          4466 => x"d6",
          4467 => x"cc",
          4468 => x"98",
          4469 => x"11",
          4470 => x"57",
          4471 => x"74",
          4472 => x"81",
          4473 => x"0c",
          4474 => x"81",
          4475 => x"84",
          4476 => x"55",
          4477 => x"ff",
          4478 => x"54",
          4479 => x"cc",
          4480 => x"0d",
          4481 => x"0d",
          4482 => x"08",
          4483 => x"79",
          4484 => x"17",
          4485 => x"80",
          4486 => x"98",
          4487 => x"26",
          4488 => x"58",
          4489 => x"52",
          4490 => x"fd",
          4491 => x"74",
          4492 => x"08",
          4493 => x"38",
          4494 => x"08",
          4495 => x"cc",
          4496 => x"82",
          4497 => x"17",
          4498 => x"cc",
          4499 => x"c7",
          4500 => x"90",
          4501 => x"56",
          4502 => x"2e",
          4503 => x"77",
          4504 => x"81",
          4505 => x"38",
          4506 => x"98",
          4507 => x"26",
          4508 => x"56",
          4509 => x"51",
          4510 => x"80",
          4511 => x"cc",
          4512 => x"09",
          4513 => x"38",
          4514 => x"08",
          4515 => x"cc",
          4516 => x"30",
          4517 => x"80",
          4518 => x"07",
          4519 => x"08",
          4520 => x"55",
          4521 => x"ef",
          4522 => x"cc",
          4523 => x"95",
          4524 => x"08",
          4525 => x"27",
          4526 => x"98",
          4527 => x"89",
          4528 => x"85",
          4529 => x"db",
          4530 => x"81",
          4531 => x"17",
          4532 => x"89",
          4533 => x"75",
          4534 => x"ac",
          4535 => x"7a",
          4536 => x"3f",
          4537 => x"08",
          4538 => x"38",
          4539 => x"87",
          4540 => x"2e",
          4541 => x"86",
          4542 => x"cc",
          4543 => x"87",
          4544 => x"70",
          4545 => x"07",
          4546 => x"7c",
          4547 => x"55",
          4548 => x"f8",
          4549 => x"2e",
          4550 => x"ff",
          4551 => x"55",
          4552 => x"ff",
          4553 => x"76",
          4554 => x"3f",
          4555 => x"08",
          4556 => x"08",
          4557 => x"87",
          4558 => x"80",
          4559 => x"55",
          4560 => x"94",
          4561 => x"2e",
          4562 => x"53",
          4563 => x"51",
          4564 => x"82",
          4565 => x"55",
          4566 => x"75",
          4567 => x"98",
          4568 => x"05",
          4569 => x"56",
          4570 => x"26",
          4571 => x"15",
          4572 => x"84",
          4573 => x"07",
          4574 => x"18",
          4575 => x"ff",
          4576 => x"2e",
          4577 => x"39",
          4578 => x"39",
          4579 => x"08",
          4580 => x"81",
          4581 => x"74",
          4582 => x"0c",
          4583 => x"04",
          4584 => x"7a",
          4585 => x"f3",
          4586 => x"87",
          4587 => x"81",
          4588 => x"cc",
          4589 => x"38",
          4590 => x"51",
          4591 => x"82",
          4592 => x"82",
          4593 => x"b0",
          4594 => x"84",
          4595 => x"52",
          4596 => x"52",
          4597 => x"3f",
          4598 => x"39",
          4599 => x"8a",
          4600 => x"75",
          4601 => x"38",
          4602 => x"19",
          4603 => x"81",
          4604 => x"ed",
          4605 => x"87",
          4606 => x"2e",
          4607 => x"15",
          4608 => x"70",
          4609 => x"07",
          4610 => x"53",
          4611 => x"75",
          4612 => x"0c",
          4613 => x"04",
          4614 => x"7a",
          4615 => x"58",
          4616 => x"f0",
          4617 => x"80",
          4618 => x"9f",
          4619 => x"80",
          4620 => x"90",
          4621 => x"17",
          4622 => x"aa",
          4623 => x"53",
          4624 => x"88",
          4625 => x"08",
          4626 => x"38",
          4627 => x"53",
          4628 => x"17",
          4629 => x"72",
          4630 => x"fe",
          4631 => x"08",
          4632 => x"80",
          4633 => x"16",
          4634 => x"2b",
          4635 => x"75",
          4636 => x"73",
          4637 => x"f5",
          4638 => x"87",
          4639 => x"82",
          4640 => x"ff",
          4641 => x"81",
          4642 => x"cc",
          4643 => x"38",
          4644 => x"82",
          4645 => x"26",
          4646 => x"58",
          4647 => x"73",
          4648 => x"39",
          4649 => x"51",
          4650 => x"82",
          4651 => x"98",
          4652 => x"94",
          4653 => x"17",
          4654 => x"58",
          4655 => x"9a",
          4656 => x"81",
          4657 => x"74",
          4658 => x"98",
          4659 => x"83",
          4660 => x"b4",
          4661 => x"0c",
          4662 => x"82",
          4663 => x"8a",
          4664 => x"f8",
          4665 => x"70",
          4666 => x"08",
          4667 => x"57",
          4668 => x"0a",
          4669 => x"38",
          4670 => x"15",
          4671 => x"08",
          4672 => x"72",
          4673 => x"cb",
          4674 => x"ff",
          4675 => x"81",
          4676 => x"13",
          4677 => x"94",
          4678 => x"74",
          4679 => x"85",
          4680 => x"22",
          4681 => x"73",
          4682 => x"38",
          4683 => x"8a",
          4684 => x"05",
          4685 => x"06",
          4686 => x"8a",
          4687 => x"73",
          4688 => x"3f",
          4689 => x"08",
          4690 => x"81",
          4691 => x"cc",
          4692 => x"ff",
          4693 => x"82",
          4694 => x"ff",
          4695 => x"38",
          4696 => x"82",
          4697 => x"26",
          4698 => x"7b",
          4699 => x"98",
          4700 => x"55",
          4701 => x"94",
          4702 => x"73",
          4703 => x"3f",
          4704 => x"08",
          4705 => x"82",
          4706 => x"80",
          4707 => x"38",
          4708 => x"87",
          4709 => x"2e",
          4710 => x"55",
          4711 => x"08",
          4712 => x"38",
          4713 => x"08",
          4714 => x"fb",
          4715 => x"87",
          4716 => x"38",
          4717 => x"0c",
          4718 => x"51",
          4719 => x"82",
          4720 => x"98",
          4721 => x"90",
          4722 => x"16",
          4723 => x"15",
          4724 => x"74",
          4725 => x"0c",
          4726 => x"04",
          4727 => x"7b",
          4728 => x"5b",
          4729 => x"52",
          4730 => x"ac",
          4731 => x"cc",
          4732 => x"87",
          4733 => x"ec",
          4734 => x"cc",
          4735 => x"17",
          4736 => x"51",
          4737 => x"82",
          4738 => x"54",
          4739 => x"08",
          4740 => x"82",
          4741 => x"9c",
          4742 => x"33",
          4743 => x"72",
          4744 => x"09",
          4745 => x"38",
          4746 => x"87",
          4747 => x"72",
          4748 => x"55",
          4749 => x"53",
          4750 => x"8e",
          4751 => x"56",
          4752 => x"09",
          4753 => x"38",
          4754 => x"87",
          4755 => x"81",
          4756 => x"fd",
          4757 => x"87",
          4758 => x"82",
          4759 => x"80",
          4760 => x"38",
          4761 => x"09",
          4762 => x"38",
          4763 => x"82",
          4764 => x"8b",
          4765 => x"fd",
          4766 => x"9a",
          4767 => x"eb",
          4768 => x"87",
          4769 => x"ff",
          4770 => x"70",
          4771 => x"53",
          4772 => x"09",
          4773 => x"38",
          4774 => x"eb",
          4775 => x"87",
          4776 => x"2b",
          4777 => x"72",
          4778 => x"0c",
          4779 => x"04",
          4780 => x"77",
          4781 => x"ff",
          4782 => x"9a",
          4783 => x"55",
          4784 => x"76",
          4785 => x"53",
          4786 => x"09",
          4787 => x"38",
          4788 => x"52",
          4789 => x"eb",
          4790 => x"3d",
          4791 => x"3d",
          4792 => x"5b",
          4793 => x"08",
          4794 => x"15",
          4795 => x"81",
          4796 => x"15",
          4797 => x"51",
          4798 => x"82",
          4799 => x"58",
          4800 => x"08",
          4801 => x"9c",
          4802 => x"33",
          4803 => x"86",
          4804 => x"80",
          4805 => x"13",
          4806 => x"06",
          4807 => x"06",
          4808 => x"72",
          4809 => x"82",
          4810 => x"53",
          4811 => x"2e",
          4812 => x"53",
          4813 => x"a9",
          4814 => x"74",
          4815 => x"72",
          4816 => x"38",
          4817 => x"99",
          4818 => x"cc",
          4819 => x"06",
          4820 => x"88",
          4821 => x"06",
          4822 => x"54",
          4823 => x"a0",
          4824 => x"74",
          4825 => x"3f",
          4826 => x"08",
          4827 => x"cc",
          4828 => x"98",
          4829 => x"fa",
          4830 => x"80",
          4831 => x"0c",
          4832 => x"cc",
          4833 => x"0d",
          4834 => x"0d",
          4835 => x"57",
          4836 => x"73",
          4837 => x"3f",
          4838 => x"08",
          4839 => x"cc",
          4840 => x"98",
          4841 => x"75",
          4842 => x"3f",
          4843 => x"08",
          4844 => x"cc",
          4845 => x"a0",
          4846 => x"cc",
          4847 => x"14",
          4848 => x"db",
          4849 => x"a0",
          4850 => x"14",
          4851 => x"ac",
          4852 => x"83",
          4853 => x"82",
          4854 => x"87",
          4855 => x"fd",
          4856 => x"70",
          4857 => x"08",
          4858 => x"55",
          4859 => x"3f",
          4860 => x"08",
          4861 => x"13",
          4862 => x"73",
          4863 => x"83",
          4864 => x"3d",
          4865 => x"3d",
          4866 => x"57",
          4867 => x"89",
          4868 => x"17",
          4869 => x"81",
          4870 => x"70",
          4871 => x"55",
          4872 => x"08",
          4873 => x"81",
          4874 => x"52",
          4875 => x"a8",
          4876 => x"2e",
          4877 => x"84",
          4878 => x"52",
          4879 => x"09",
          4880 => x"38",
          4881 => x"81",
          4882 => x"81",
          4883 => x"73",
          4884 => x"55",
          4885 => x"55",
          4886 => x"c5",
          4887 => x"88",
          4888 => x"0b",
          4889 => x"9c",
          4890 => x"8b",
          4891 => x"17",
          4892 => x"08",
          4893 => x"52",
          4894 => x"82",
          4895 => x"76",
          4896 => x"51",
          4897 => x"82",
          4898 => x"86",
          4899 => x"12",
          4900 => x"3f",
          4901 => x"08",
          4902 => x"88",
          4903 => x"f3",
          4904 => x"70",
          4905 => x"80",
          4906 => x"51",
          4907 => x"af",
          4908 => x"81",
          4909 => x"dc",
          4910 => x"74",
          4911 => x"38",
          4912 => x"88",
          4913 => x"39",
          4914 => x"80",
          4915 => x"56",
          4916 => x"af",
          4917 => x"06",
          4918 => x"56",
          4919 => x"32",
          4920 => x"80",
          4921 => x"51",
          4922 => x"dc",
          4923 => x"1c",
          4924 => x"33",
          4925 => x"9f",
          4926 => x"ff",
          4927 => x"1c",
          4928 => x"7a",
          4929 => x"3f",
          4930 => x"08",
          4931 => x"39",
          4932 => x"a0",
          4933 => x"5e",
          4934 => x"52",
          4935 => x"ff",
          4936 => x"59",
          4937 => x"33",
          4938 => x"ae",
          4939 => x"06",
          4940 => x"78",
          4941 => x"81",
          4942 => x"32",
          4943 => x"9f",
          4944 => x"26",
          4945 => x"53",
          4946 => x"73",
          4947 => x"17",
          4948 => x"34",
          4949 => x"db",
          4950 => x"32",
          4951 => x"9f",
          4952 => x"54",
          4953 => x"2e",
          4954 => x"80",
          4955 => x"75",
          4956 => x"bd",
          4957 => x"7e",
          4958 => x"a0",
          4959 => x"bd",
          4960 => x"82",
          4961 => x"18",
          4962 => x"1a",
          4963 => x"a0",
          4964 => x"fc",
          4965 => x"32",
          4966 => x"80",
          4967 => x"30",
          4968 => x"71",
          4969 => x"51",
          4970 => x"55",
          4971 => x"ac",
          4972 => x"81",
          4973 => x"78",
          4974 => x"51",
          4975 => x"af",
          4976 => x"06",
          4977 => x"55",
          4978 => x"32",
          4979 => x"80",
          4980 => x"51",
          4981 => x"db",
          4982 => x"39",
          4983 => x"09",
          4984 => x"38",
          4985 => x"7c",
          4986 => x"54",
          4987 => x"a2",
          4988 => x"32",
          4989 => x"ae",
          4990 => x"72",
          4991 => x"9f",
          4992 => x"51",
          4993 => x"74",
          4994 => x"88",
          4995 => x"fe",
          4996 => x"98",
          4997 => x"80",
          4998 => x"75",
          4999 => x"82",
          5000 => x"33",
          5001 => x"51",
          5002 => x"82",
          5003 => x"80",
          5004 => x"78",
          5005 => x"81",
          5006 => x"5a",
          5007 => x"d2",
          5008 => x"cc",
          5009 => x"80",
          5010 => x"1c",
          5011 => x"27",
          5012 => x"79",
          5013 => x"74",
          5014 => x"7a",
          5015 => x"74",
          5016 => x"39",
          5017 => x"80",
          5018 => x"fe",
          5019 => x"cc",
          5020 => x"ff",
          5021 => x"73",
          5022 => x"38",
          5023 => x"81",
          5024 => x"54",
          5025 => x"75",
          5026 => x"17",
          5027 => x"39",
          5028 => x"0c",
          5029 => x"99",
          5030 => x"54",
          5031 => x"2e",
          5032 => x"84",
          5033 => x"34",
          5034 => x"76",
          5035 => x"8b",
          5036 => x"81",
          5037 => x"56",
          5038 => x"80",
          5039 => x"1b",
          5040 => x"08",
          5041 => x"51",
          5042 => x"82",
          5043 => x"56",
          5044 => x"08",
          5045 => x"98",
          5046 => x"76",
          5047 => x"3f",
          5048 => x"08",
          5049 => x"cc",
          5050 => x"38",
          5051 => x"70",
          5052 => x"73",
          5053 => x"be",
          5054 => x"33",
          5055 => x"73",
          5056 => x"8b",
          5057 => x"83",
          5058 => x"06",
          5059 => x"73",
          5060 => x"53",
          5061 => x"51",
          5062 => x"82",
          5063 => x"80",
          5064 => x"75",
          5065 => x"f3",
          5066 => x"9f",
          5067 => x"1c",
          5068 => x"74",
          5069 => x"38",
          5070 => x"09",
          5071 => x"e7",
          5072 => x"2a",
          5073 => x"77",
          5074 => x"51",
          5075 => x"2e",
          5076 => x"81",
          5077 => x"80",
          5078 => x"38",
          5079 => x"ab",
          5080 => x"55",
          5081 => x"75",
          5082 => x"73",
          5083 => x"55",
          5084 => x"82",
          5085 => x"06",
          5086 => x"ab",
          5087 => x"33",
          5088 => x"70",
          5089 => x"55",
          5090 => x"2e",
          5091 => x"1b",
          5092 => x"06",
          5093 => x"52",
          5094 => x"db",
          5095 => x"cc",
          5096 => x"0c",
          5097 => x"74",
          5098 => x"0c",
          5099 => x"04",
          5100 => x"7c",
          5101 => x"08",
          5102 => x"55",
          5103 => x"59",
          5104 => x"81",
          5105 => x"70",
          5106 => x"33",
          5107 => x"52",
          5108 => x"2e",
          5109 => x"ee",
          5110 => x"2e",
          5111 => x"81",
          5112 => x"33",
          5113 => x"81",
          5114 => x"52",
          5115 => x"26",
          5116 => x"14",
          5117 => x"06",
          5118 => x"52",
          5119 => x"80",
          5120 => x"0b",
          5121 => x"59",
          5122 => x"7a",
          5123 => x"70",
          5124 => x"33",
          5125 => x"05",
          5126 => x"9f",
          5127 => x"53",
          5128 => x"89",
          5129 => x"70",
          5130 => x"54",
          5131 => x"12",
          5132 => x"26",
          5133 => x"12",
          5134 => x"06",
          5135 => x"30",
          5136 => x"51",
          5137 => x"2e",
          5138 => x"85",
          5139 => x"be",
          5140 => x"74",
          5141 => x"30",
          5142 => x"9f",
          5143 => x"2a",
          5144 => x"54",
          5145 => x"2e",
          5146 => x"15",
          5147 => x"55",
          5148 => x"ff",
          5149 => x"39",
          5150 => x"86",
          5151 => x"7c",
          5152 => x"51",
          5153 => x"9f",
          5154 => x"70",
          5155 => x"0c",
          5156 => x"04",
          5157 => x"78",
          5158 => x"83",
          5159 => x"0b",
          5160 => x"79",
          5161 => x"e2",
          5162 => x"55",
          5163 => x"08",
          5164 => x"84",
          5165 => x"df",
          5166 => x"87",
          5167 => x"ff",
          5168 => x"83",
          5169 => x"d4",
          5170 => x"81",
          5171 => x"38",
          5172 => x"17",
          5173 => x"74",
          5174 => x"09",
          5175 => x"38",
          5176 => x"81",
          5177 => x"30",
          5178 => x"79",
          5179 => x"54",
          5180 => x"74",
          5181 => x"09",
          5182 => x"38",
          5183 => x"80",
          5184 => x"ea",
          5185 => x"b1",
          5186 => x"cc",
          5187 => x"87",
          5188 => x"2e",
          5189 => x"53",
          5190 => x"52",
          5191 => x"51",
          5192 => x"82",
          5193 => x"55",
          5194 => x"08",
          5195 => x"38",
          5196 => x"82",
          5197 => x"88",
          5198 => x"f2",
          5199 => x"02",
          5200 => x"cb",
          5201 => x"55",
          5202 => x"60",
          5203 => x"3f",
          5204 => x"08",
          5205 => x"80",
          5206 => x"cc",
          5207 => x"fb",
          5208 => x"cc",
          5209 => x"82",
          5210 => x"70",
          5211 => x"8c",
          5212 => x"2e",
          5213 => x"73",
          5214 => x"81",
          5215 => x"33",
          5216 => x"80",
          5217 => x"81",
          5218 => x"d7",
          5219 => x"87",
          5220 => x"ff",
          5221 => x"06",
          5222 => x"98",
          5223 => x"2e",
          5224 => x"74",
          5225 => x"81",
          5226 => x"8a",
          5227 => x"ab",
          5228 => x"39",
          5229 => x"77",
          5230 => x"81",
          5231 => x"33",
          5232 => x"3f",
          5233 => x"08",
          5234 => x"70",
          5235 => x"55",
          5236 => x"86",
          5237 => x"80",
          5238 => x"74",
          5239 => x"81",
          5240 => x"8a",
          5241 => x"f3",
          5242 => x"53",
          5243 => x"fd",
          5244 => x"87",
          5245 => x"ff",
          5246 => x"82",
          5247 => x"06",
          5248 => x"8c",
          5249 => x"58",
          5250 => x"f6",
          5251 => x"58",
          5252 => x"2e",
          5253 => x"fa",
          5254 => x"e8",
          5255 => x"cc",
          5256 => x"78",
          5257 => x"5a",
          5258 => x"90",
          5259 => x"75",
          5260 => x"38",
          5261 => x"3d",
          5262 => x"70",
          5263 => x"08",
          5264 => x"7a",
          5265 => x"38",
          5266 => x"51",
          5267 => x"82",
          5268 => x"81",
          5269 => x"81",
          5270 => x"38",
          5271 => x"83",
          5272 => x"38",
          5273 => x"84",
          5274 => x"38",
          5275 => x"81",
          5276 => x"38",
          5277 => x"db",
          5278 => x"87",
          5279 => x"ff",
          5280 => x"72",
          5281 => x"09",
          5282 => x"cf",
          5283 => x"14",
          5284 => x"3f",
          5285 => x"08",
          5286 => x"06",
          5287 => x"38",
          5288 => x"51",
          5289 => x"82",
          5290 => x"58",
          5291 => x"0c",
          5292 => x"33",
          5293 => x"80",
          5294 => x"ff",
          5295 => x"ff",
          5296 => x"55",
          5297 => x"81",
          5298 => x"38",
          5299 => x"06",
          5300 => x"80",
          5301 => x"52",
          5302 => x"8a",
          5303 => x"80",
          5304 => x"ff",
          5305 => x"53",
          5306 => x"86",
          5307 => x"83",
          5308 => x"c5",
          5309 => x"f5",
          5310 => x"cc",
          5311 => x"87",
          5312 => x"15",
          5313 => x"06",
          5314 => x"76",
          5315 => x"80",
          5316 => x"da",
          5317 => x"87",
          5318 => x"ff",
          5319 => x"74",
          5320 => x"d4",
          5321 => x"dc",
          5322 => x"cc",
          5323 => x"c2",
          5324 => x"b9",
          5325 => x"cc",
          5326 => x"ff",
          5327 => x"56",
          5328 => x"83",
          5329 => x"14",
          5330 => x"71",
          5331 => x"5a",
          5332 => x"26",
          5333 => x"8a",
          5334 => x"74",
          5335 => x"c5",
          5336 => x"87",
          5337 => x"82",
          5338 => x"80",
          5339 => x"38",
          5340 => x"08",
          5341 => x"ff",
          5342 => x"38",
          5343 => x"83",
          5344 => x"83",
          5345 => x"74",
          5346 => x"85",
          5347 => x"89",
          5348 => x"76",
          5349 => x"c3",
          5350 => x"70",
          5351 => x"7b",
          5352 => x"73",
          5353 => x"17",
          5354 => x"ac",
          5355 => x"55",
          5356 => x"09",
          5357 => x"38",
          5358 => x"51",
          5359 => x"82",
          5360 => x"83",
          5361 => x"53",
          5362 => x"82",
          5363 => x"82",
          5364 => x"e0",
          5365 => x"ac",
          5366 => x"cc",
          5367 => x"0c",
          5368 => x"53",
          5369 => x"56",
          5370 => x"81",
          5371 => x"13",
          5372 => x"74",
          5373 => x"82",
          5374 => x"74",
          5375 => x"81",
          5376 => x"06",
          5377 => x"83",
          5378 => x"2a",
          5379 => x"72",
          5380 => x"26",
          5381 => x"ff",
          5382 => x"0c",
          5383 => x"15",
          5384 => x"0b",
          5385 => x"76",
          5386 => x"81",
          5387 => x"38",
          5388 => x"51",
          5389 => x"82",
          5390 => x"83",
          5391 => x"53",
          5392 => x"09",
          5393 => x"f9",
          5394 => x"52",
          5395 => x"b9",
          5396 => x"cc",
          5397 => x"38",
          5398 => x"08",
          5399 => x"84",
          5400 => x"d8",
          5401 => x"87",
          5402 => x"ff",
          5403 => x"72",
          5404 => x"2e",
          5405 => x"80",
          5406 => x"14",
          5407 => x"3f",
          5408 => x"08",
          5409 => x"a4",
          5410 => x"81",
          5411 => x"84",
          5412 => x"d7",
          5413 => x"87",
          5414 => x"8a",
          5415 => x"2e",
          5416 => x"9d",
          5417 => x"14",
          5418 => x"3f",
          5419 => x"08",
          5420 => x"84",
          5421 => x"d7",
          5422 => x"87",
          5423 => x"15",
          5424 => x"34",
          5425 => x"22",
          5426 => x"72",
          5427 => x"23",
          5428 => x"23",
          5429 => x"15",
          5430 => x"75",
          5431 => x"0c",
          5432 => x"04",
          5433 => x"77",
          5434 => x"73",
          5435 => x"38",
          5436 => x"72",
          5437 => x"38",
          5438 => x"71",
          5439 => x"38",
          5440 => x"84",
          5441 => x"52",
          5442 => x"09",
          5443 => x"38",
          5444 => x"51",
          5445 => x"82",
          5446 => x"81",
          5447 => x"88",
          5448 => x"08",
          5449 => x"39",
          5450 => x"73",
          5451 => x"74",
          5452 => x"0c",
          5453 => x"04",
          5454 => x"02",
          5455 => x"7a",
          5456 => x"fc",
          5457 => x"f4",
          5458 => x"54",
          5459 => x"87",
          5460 => x"bc",
          5461 => x"cc",
          5462 => x"82",
          5463 => x"70",
          5464 => x"73",
          5465 => x"38",
          5466 => x"78",
          5467 => x"2e",
          5468 => x"74",
          5469 => x"0c",
          5470 => x"80",
          5471 => x"80",
          5472 => x"70",
          5473 => x"51",
          5474 => x"82",
          5475 => x"54",
          5476 => x"cc",
          5477 => x"0d",
          5478 => x"0d",
          5479 => x"05",
          5480 => x"33",
          5481 => x"54",
          5482 => x"84",
          5483 => x"bf",
          5484 => x"98",
          5485 => x"53",
          5486 => x"05",
          5487 => x"fb",
          5488 => x"cc",
          5489 => x"87",
          5490 => x"a4",
          5491 => x"68",
          5492 => x"70",
          5493 => x"c7",
          5494 => x"cc",
          5495 => x"87",
          5496 => x"38",
          5497 => x"05",
          5498 => x"2b",
          5499 => x"80",
          5500 => x"86",
          5501 => x"06",
          5502 => x"2e",
          5503 => x"74",
          5504 => x"38",
          5505 => x"09",
          5506 => x"38",
          5507 => x"f9",
          5508 => x"cc",
          5509 => x"39",
          5510 => x"33",
          5511 => x"73",
          5512 => x"77",
          5513 => x"81",
          5514 => x"73",
          5515 => x"38",
          5516 => x"bc",
          5517 => x"07",
          5518 => x"b4",
          5519 => x"2a",
          5520 => x"51",
          5521 => x"2e",
          5522 => x"62",
          5523 => x"e8",
          5524 => x"87",
          5525 => x"82",
          5526 => x"52",
          5527 => x"51",
          5528 => x"62",
          5529 => x"8b",
          5530 => x"53",
          5531 => x"51",
          5532 => x"80",
          5533 => x"05",
          5534 => x"3f",
          5535 => x"0b",
          5536 => x"75",
          5537 => x"f1",
          5538 => x"11",
          5539 => x"80",
          5540 => x"97",
          5541 => x"51",
          5542 => x"82",
          5543 => x"55",
          5544 => x"08",
          5545 => x"b7",
          5546 => x"c4",
          5547 => x"05",
          5548 => x"2a",
          5549 => x"51",
          5550 => x"80",
          5551 => x"84",
          5552 => x"39",
          5553 => x"70",
          5554 => x"54",
          5555 => x"a9",
          5556 => x"06",
          5557 => x"2e",
          5558 => x"55",
          5559 => x"73",
          5560 => x"d6",
          5561 => x"87",
          5562 => x"ff",
          5563 => x"0c",
          5564 => x"87",
          5565 => x"f8",
          5566 => x"2a",
          5567 => x"51",
          5568 => x"2e",
          5569 => x"80",
          5570 => x"7a",
          5571 => x"a0",
          5572 => x"a4",
          5573 => x"53",
          5574 => x"e6",
          5575 => x"87",
          5576 => x"87",
          5577 => x"1b",
          5578 => x"05",
          5579 => x"d4",
          5580 => x"cc",
          5581 => x"cc",
          5582 => x"0c",
          5583 => x"56",
          5584 => x"84",
          5585 => x"90",
          5586 => x"0b",
          5587 => x"80",
          5588 => x"0c",
          5589 => x"1a",
          5590 => x"2a",
          5591 => x"51",
          5592 => x"2e",
          5593 => x"82",
          5594 => x"80",
          5595 => x"38",
          5596 => x"08",
          5597 => x"8a",
          5598 => x"89",
          5599 => x"59",
          5600 => x"76",
          5601 => x"d7",
          5602 => x"87",
          5603 => x"82",
          5604 => x"81",
          5605 => x"82",
          5606 => x"cc",
          5607 => x"09",
          5608 => x"38",
          5609 => x"78",
          5610 => x"30",
          5611 => x"80",
          5612 => x"77",
          5613 => x"38",
          5614 => x"06",
          5615 => x"c3",
          5616 => x"1a",
          5617 => x"38",
          5618 => x"06",
          5619 => x"2e",
          5620 => x"52",
          5621 => x"a7",
          5622 => x"cc",
          5623 => x"82",
          5624 => x"75",
          5625 => x"87",
          5626 => x"9c",
          5627 => x"39",
          5628 => x"74",
          5629 => x"87",
          5630 => x"3d",
          5631 => x"3d",
          5632 => x"65",
          5633 => x"5d",
          5634 => x"0c",
          5635 => x"05",
          5636 => x"f9",
          5637 => x"87",
          5638 => x"82",
          5639 => x"8a",
          5640 => x"33",
          5641 => x"2e",
          5642 => x"56",
          5643 => x"90",
          5644 => x"06",
          5645 => x"74",
          5646 => x"b6",
          5647 => x"82",
          5648 => x"34",
          5649 => x"aa",
          5650 => x"91",
          5651 => x"56",
          5652 => x"8c",
          5653 => x"1a",
          5654 => x"74",
          5655 => x"38",
          5656 => x"80",
          5657 => x"38",
          5658 => x"70",
          5659 => x"56",
          5660 => x"b2",
          5661 => x"11",
          5662 => x"77",
          5663 => x"5b",
          5664 => x"38",
          5665 => x"88",
          5666 => x"8f",
          5667 => x"08",
          5668 => x"d5",
          5669 => x"87",
          5670 => x"81",
          5671 => x"9f",
          5672 => x"2e",
          5673 => x"74",
          5674 => x"98",
          5675 => x"7e",
          5676 => x"3f",
          5677 => x"08",
          5678 => x"83",
          5679 => x"cc",
          5680 => x"89",
          5681 => x"77",
          5682 => x"d6",
          5683 => x"7f",
          5684 => x"58",
          5685 => x"75",
          5686 => x"75",
          5687 => x"77",
          5688 => x"7c",
          5689 => x"33",
          5690 => x"3f",
          5691 => x"08",
          5692 => x"7e",
          5693 => x"56",
          5694 => x"2e",
          5695 => x"16",
          5696 => x"55",
          5697 => x"94",
          5698 => x"53",
          5699 => x"b0",
          5700 => x"31",
          5701 => x"05",
          5702 => x"3f",
          5703 => x"56",
          5704 => x"9c",
          5705 => x"19",
          5706 => x"06",
          5707 => x"31",
          5708 => x"76",
          5709 => x"7b",
          5710 => x"08",
          5711 => x"d1",
          5712 => x"87",
          5713 => x"81",
          5714 => x"94",
          5715 => x"ff",
          5716 => x"05",
          5717 => x"cf",
          5718 => x"76",
          5719 => x"17",
          5720 => x"1e",
          5721 => x"18",
          5722 => x"5e",
          5723 => x"39",
          5724 => x"82",
          5725 => x"90",
          5726 => x"f2",
          5727 => x"63",
          5728 => x"40",
          5729 => x"7e",
          5730 => x"fc",
          5731 => x"51",
          5732 => x"82",
          5733 => x"55",
          5734 => x"08",
          5735 => x"18",
          5736 => x"80",
          5737 => x"74",
          5738 => x"39",
          5739 => x"70",
          5740 => x"81",
          5741 => x"56",
          5742 => x"80",
          5743 => x"38",
          5744 => x"0b",
          5745 => x"82",
          5746 => x"39",
          5747 => x"19",
          5748 => x"83",
          5749 => x"18",
          5750 => x"56",
          5751 => x"27",
          5752 => x"09",
          5753 => x"2e",
          5754 => x"94",
          5755 => x"83",
          5756 => x"56",
          5757 => x"38",
          5758 => x"22",
          5759 => x"89",
          5760 => x"55",
          5761 => x"75",
          5762 => x"18",
          5763 => x"9c",
          5764 => x"85",
          5765 => x"08",
          5766 => x"d7",
          5767 => x"87",
          5768 => x"82",
          5769 => x"80",
          5770 => x"38",
          5771 => x"ff",
          5772 => x"ff",
          5773 => x"38",
          5774 => x"0c",
          5775 => x"85",
          5776 => x"19",
          5777 => x"b0",
          5778 => x"19",
          5779 => x"81",
          5780 => x"74",
          5781 => x"3f",
          5782 => x"08",
          5783 => x"98",
          5784 => x"7e",
          5785 => x"3f",
          5786 => x"08",
          5787 => x"d2",
          5788 => x"cc",
          5789 => x"89",
          5790 => x"78",
          5791 => x"d5",
          5792 => x"7f",
          5793 => x"58",
          5794 => x"75",
          5795 => x"75",
          5796 => x"78",
          5797 => x"7c",
          5798 => x"33",
          5799 => x"3f",
          5800 => x"08",
          5801 => x"7e",
          5802 => x"78",
          5803 => x"74",
          5804 => x"38",
          5805 => x"b0",
          5806 => x"31",
          5807 => x"05",
          5808 => x"51",
          5809 => x"7e",
          5810 => x"83",
          5811 => x"89",
          5812 => x"db",
          5813 => x"08",
          5814 => x"26",
          5815 => x"51",
          5816 => x"82",
          5817 => x"fd",
          5818 => x"77",
          5819 => x"55",
          5820 => x"0c",
          5821 => x"83",
          5822 => x"80",
          5823 => x"55",
          5824 => x"83",
          5825 => x"9c",
          5826 => x"7e",
          5827 => x"3f",
          5828 => x"08",
          5829 => x"75",
          5830 => x"94",
          5831 => x"ff",
          5832 => x"05",
          5833 => x"3f",
          5834 => x"0b",
          5835 => x"7b",
          5836 => x"08",
          5837 => x"76",
          5838 => x"08",
          5839 => x"1c",
          5840 => x"08",
          5841 => x"5c",
          5842 => x"83",
          5843 => x"74",
          5844 => x"fd",
          5845 => x"18",
          5846 => x"07",
          5847 => x"19",
          5848 => x"75",
          5849 => x"0c",
          5850 => x"04",
          5851 => x"7a",
          5852 => x"05",
          5853 => x"56",
          5854 => x"82",
          5855 => x"57",
          5856 => x"08",
          5857 => x"90",
          5858 => x"86",
          5859 => x"06",
          5860 => x"73",
          5861 => x"e9",
          5862 => x"08",
          5863 => x"cc",
          5864 => x"87",
          5865 => x"82",
          5866 => x"80",
          5867 => x"16",
          5868 => x"33",
          5869 => x"55",
          5870 => x"34",
          5871 => x"53",
          5872 => x"08",
          5873 => x"3f",
          5874 => x"52",
          5875 => x"c9",
          5876 => x"88",
          5877 => x"96",
          5878 => x"f1",
          5879 => x"92",
          5880 => x"cb",
          5881 => x"81",
          5882 => x"34",
          5883 => x"e0",
          5884 => x"cc",
          5885 => x"33",
          5886 => x"55",
          5887 => x"17",
          5888 => x"87",
          5889 => x"3d",
          5890 => x"3d",
          5891 => x"52",
          5892 => x"3f",
          5893 => x"08",
          5894 => x"cc",
          5895 => x"86",
          5896 => x"52",
          5897 => x"bc",
          5898 => x"cc",
          5899 => x"87",
          5900 => x"38",
          5901 => x"08",
          5902 => x"82",
          5903 => x"86",
          5904 => x"ff",
          5905 => x"3d",
          5906 => x"3f",
          5907 => x"0b",
          5908 => x"08",
          5909 => x"82",
          5910 => x"82",
          5911 => x"80",
          5912 => x"87",
          5913 => x"3d",
          5914 => x"3d",
          5915 => x"93",
          5916 => x"52",
          5917 => x"e9",
          5918 => x"87",
          5919 => x"82",
          5920 => x"80",
          5921 => x"58",
          5922 => x"3d",
          5923 => x"e0",
          5924 => x"87",
          5925 => x"82",
          5926 => x"bc",
          5927 => x"c7",
          5928 => x"98",
          5929 => x"73",
          5930 => x"38",
          5931 => x"12",
          5932 => x"39",
          5933 => x"33",
          5934 => x"70",
          5935 => x"55",
          5936 => x"2e",
          5937 => x"7f",
          5938 => x"54",
          5939 => x"82",
          5940 => x"94",
          5941 => x"39",
          5942 => x"08",
          5943 => x"81",
          5944 => x"85",
          5945 => x"87",
          5946 => x"3d",
          5947 => x"3d",
          5948 => x"5b",
          5949 => x"34",
          5950 => x"3d",
          5951 => x"52",
          5952 => x"e8",
          5953 => x"87",
          5954 => x"82",
          5955 => x"82",
          5956 => x"43",
          5957 => x"11",
          5958 => x"58",
          5959 => x"80",
          5960 => x"38",
          5961 => x"3d",
          5962 => x"d5",
          5963 => x"87",
          5964 => x"82",
          5965 => x"82",
          5966 => x"52",
          5967 => x"c9",
          5968 => x"cc",
          5969 => x"87",
          5970 => x"c1",
          5971 => x"7b",
          5972 => x"3f",
          5973 => x"08",
          5974 => x"74",
          5975 => x"3f",
          5976 => x"08",
          5977 => x"cc",
          5978 => x"38",
          5979 => x"51",
          5980 => x"82",
          5981 => x"57",
          5982 => x"08",
          5983 => x"52",
          5984 => x"f3",
          5985 => x"87",
          5986 => x"a6",
          5987 => x"74",
          5988 => x"3f",
          5989 => x"08",
          5990 => x"cc",
          5991 => x"cc",
          5992 => x"2e",
          5993 => x"86",
          5994 => x"81",
          5995 => x"81",
          5996 => x"3d",
          5997 => x"52",
          5998 => x"ca",
          5999 => x"3d",
          6000 => x"11",
          6001 => x"5a",
          6002 => x"2e",
          6003 => x"b9",
          6004 => x"16",
          6005 => x"33",
          6006 => x"73",
          6007 => x"16",
          6008 => x"26",
          6009 => x"75",
          6010 => x"38",
          6011 => x"05",
          6012 => x"6f",
          6013 => x"ff",
          6014 => x"55",
          6015 => x"74",
          6016 => x"38",
          6017 => x"11",
          6018 => x"74",
          6019 => x"39",
          6020 => x"09",
          6021 => x"38",
          6022 => x"11",
          6023 => x"74",
          6024 => x"82",
          6025 => x"70",
          6026 => x"81",
          6027 => x"08",
          6028 => x"5c",
          6029 => x"73",
          6030 => x"38",
          6031 => x"1a",
          6032 => x"55",
          6033 => x"38",
          6034 => x"73",
          6035 => x"38",
          6036 => x"76",
          6037 => x"74",
          6038 => x"33",
          6039 => x"05",
          6040 => x"15",
          6041 => x"ba",
          6042 => x"05",
          6043 => x"ff",
          6044 => x"06",
          6045 => x"57",
          6046 => x"18",
          6047 => x"54",
          6048 => x"70",
          6049 => x"34",
          6050 => x"ee",
          6051 => x"34",
          6052 => x"cc",
          6053 => x"0d",
          6054 => x"0d",
          6055 => x"3d",
          6056 => x"71",
          6057 => x"ec",
          6058 => x"87",
          6059 => x"82",
          6060 => x"82",
          6061 => x"15",
          6062 => x"82",
          6063 => x"15",
          6064 => x"76",
          6065 => x"90",
          6066 => x"81",
          6067 => x"06",
          6068 => x"72",
          6069 => x"56",
          6070 => x"54",
          6071 => x"17",
          6072 => x"78",
          6073 => x"38",
          6074 => x"22",
          6075 => x"59",
          6076 => x"78",
          6077 => x"76",
          6078 => x"51",
          6079 => x"3f",
          6080 => x"08",
          6081 => x"54",
          6082 => x"53",
          6083 => x"3f",
          6084 => x"08",
          6085 => x"38",
          6086 => x"75",
          6087 => x"18",
          6088 => x"31",
          6089 => x"57",
          6090 => x"b1",
          6091 => x"08",
          6092 => x"38",
          6093 => x"51",
          6094 => x"82",
          6095 => x"54",
          6096 => x"08",
          6097 => x"9a",
          6098 => x"cc",
          6099 => x"81",
          6100 => x"87",
          6101 => x"16",
          6102 => x"16",
          6103 => x"2e",
          6104 => x"76",
          6105 => x"dc",
          6106 => x"31",
          6107 => x"18",
          6108 => x"90",
          6109 => x"81",
          6110 => x"06",
          6111 => x"56",
          6112 => x"9a",
          6113 => x"74",
          6114 => x"3f",
          6115 => x"08",
          6116 => x"cc",
          6117 => x"82",
          6118 => x"56",
          6119 => x"52",
          6120 => x"85",
          6121 => x"cc",
          6122 => x"ff",
          6123 => x"81",
          6124 => x"38",
          6125 => x"98",
          6126 => x"a6",
          6127 => x"16",
          6128 => x"39",
          6129 => x"16",
          6130 => x"75",
          6131 => x"53",
          6132 => x"aa",
          6133 => x"79",
          6134 => x"3f",
          6135 => x"08",
          6136 => x"0b",
          6137 => x"82",
          6138 => x"39",
          6139 => x"16",
          6140 => x"bb",
          6141 => x"2a",
          6142 => x"08",
          6143 => x"15",
          6144 => x"15",
          6145 => x"90",
          6146 => x"16",
          6147 => x"33",
          6148 => x"53",
          6149 => x"34",
          6150 => x"06",
          6151 => x"2e",
          6152 => x"9c",
          6153 => x"85",
          6154 => x"16",
          6155 => x"72",
          6156 => x"0c",
          6157 => x"04",
          6158 => x"79",
          6159 => x"75",
          6160 => x"8a",
          6161 => x"89",
          6162 => x"52",
          6163 => x"05",
          6164 => x"3f",
          6165 => x"08",
          6166 => x"cc",
          6167 => x"38",
          6168 => x"7a",
          6169 => x"d8",
          6170 => x"87",
          6171 => x"82",
          6172 => x"80",
          6173 => x"16",
          6174 => x"2b",
          6175 => x"74",
          6176 => x"86",
          6177 => x"84",
          6178 => x"06",
          6179 => x"73",
          6180 => x"38",
          6181 => x"52",
          6182 => x"db",
          6183 => x"cc",
          6184 => x"0c",
          6185 => x"14",
          6186 => x"23",
          6187 => x"51",
          6188 => x"82",
          6189 => x"55",
          6190 => x"09",
          6191 => x"38",
          6192 => x"39",
          6193 => x"84",
          6194 => x"0c",
          6195 => x"82",
          6196 => x"89",
          6197 => x"fc",
          6198 => x"87",
          6199 => x"53",
          6200 => x"e7",
          6201 => x"87",
          6202 => x"38",
          6203 => x"08",
          6204 => x"3d",
          6205 => x"3d",
          6206 => x"89",
          6207 => x"54",
          6208 => x"54",
          6209 => x"82",
          6210 => x"53",
          6211 => x"08",
          6212 => x"74",
          6213 => x"87",
          6214 => x"73",
          6215 => x"3f",
          6216 => x"08",
          6217 => x"39",
          6218 => x"08",
          6219 => x"d3",
          6220 => x"87",
          6221 => x"82",
          6222 => x"84",
          6223 => x"06",
          6224 => x"53",
          6225 => x"87",
          6226 => x"38",
          6227 => x"51",
          6228 => x"72",
          6229 => x"cf",
          6230 => x"87",
          6231 => x"32",
          6232 => x"72",
          6233 => x"70",
          6234 => x"08",
          6235 => x"54",
          6236 => x"87",
          6237 => x"3d",
          6238 => x"3d",
          6239 => x"80",
          6240 => x"70",
          6241 => x"52",
          6242 => x"3f",
          6243 => x"08",
          6244 => x"cc",
          6245 => x"64",
          6246 => x"d6",
          6247 => x"87",
          6248 => x"82",
          6249 => x"a0",
          6250 => x"cb",
          6251 => x"98",
          6252 => x"73",
          6253 => x"38",
          6254 => x"39",
          6255 => x"88",
          6256 => x"75",
          6257 => x"3f",
          6258 => x"cc",
          6259 => x"0d",
          6260 => x"0d",
          6261 => x"5c",
          6262 => x"3d",
          6263 => x"93",
          6264 => x"d7",
          6265 => x"cc",
          6266 => x"87",
          6267 => x"80",
          6268 => x"0c",
          6269 => x"11",
          6270 => x"90",
          6271 => x"56",
          6272 => x"74",
          6273 => x"75",
          6274 => x"e4",
          6275 => x"81",
          6276 => x"5b",
          6277 => x"82",
          6278 => x"75",
          6279 => x"73",
          6280 => x"81",
          6281 => x"82",
          6282 => x"76",
          6283 => x"f0",
          6284 => x"f5",
          6285 => x"cc",
          6286 => x"d1",
          6287 => x"cc",
          6288 => x"ce",
          6289 => x"cc",
          6290 => x"82",
          6291 => x"07",
          6292 => x"05",
          6293 => x"53",
          6294 => x"98",
          6295 => x"26",
          6296 => x"f9",
          6297 => x"08",
          6298 => x"08",
          6299 => x"98",
          6300 => x"81",
          6301 => x"58",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"cc",
          6305 => x"38",
          6306 => x"77",
          6307 => x"5d",
          6308 => x"74",
          6309 => x"81",
          6310 => x"b4",
          6311 => x"bb",
          6312 => x"87",
          6313 => x"ff",
          6314 => x"30",
          6315 => x"1b",
          6316 => x"5b",
          6317 => x"39",
          6318 => x"ff",
          6319 => x"82",
          6320 => x"f0",
          6321 => x"30",
          6322 => x"1b",
          6323 => x"5b",
          6324 => x"83",
          6325 => x"58",
          6326 => x"92",
          6327 => x"0c",
          6328 => x"12",
          6329 => x"33",
          6330 => x"54",
          6331 => x"34",
          6332 => x"cc",
          6333 => x"0d",
          6334 => x"0d",
          6335 => x"fc",
          6336 => x"52",
          6337 => x"3f",
          6338 => x"08",
          6339 => x"cc",
          6340 => x"38",
          6341 => x"56",
          6342 => x"38",
          6343 => x"70",
          6344 => x"81",
          6345 => x"55",
          6346 => x"80",
          6347 => x"38",
          6348 => x"54",
          6349 => x"08",
          6350 => x"38",
          6351 => x"82",
          6352 => x"53",
          6353 => x"52",
          6354 => x"8d",
          6355 => x"cc",
          6356 => x"19",
          6357 => x"c9",
          6358 => x"08",
          6359 => x"ff",
          6360 => x"82",
          6361 => x"ff",
          6362 => x"06",
          6363 => x"56",
          6364 => x"08",
          6365 => x"81",
          6366 => x"82",
          6367 => x"75",
          6368 => x"54",
          6369 => x"08",
          6370 => x"27",
          6371 => x"17",
          6372 => x"87",
          6373 => x"76",
          6374 => x"3f",
          6375 => x"08",
          6376 => x"08",
          6377 => x"90",
          6378 => x"c0",
          6379 => x"90",
          6380 => x"80",
          6381 => x"75",
          6382 => x"75",
          6383 => x"87",
          6384 => x"3d",
          6385 => x"3d",
          6386 => x"a0",
          6387 => x"05",
          6388 => x"51",
          6389 => x"82",
          6390 => x"55",
          6391 => x"08",
          6392 => x"78",
          6393 => x"08",
          6394 => x"70",
          6395 => x"af",
          6396 => x"cc",
          6397 => x"87",
          6398 => x"db",
          6399 => x"fb",
          6400 => x"85",
          6401 => x"06",
          6402 => x"86",
          6403 => x"c7",
          6404 => x"2b",
          6405 => x"24",
          6406 => x"02",
          6407 => x"33",
          6408 => x"58",
          6409 => x"76",
          6410 => x"6b",
          6411 => x"cc",
          6412 => x"87",
          6413 => x"84",
          6414 => x"06",
          6415 => x"73",
          6416 => x"d4",
          6417 => x"82",
          6418 => x"94",
          6419 => x"81",
          6420 => x"5a",
          6421 => x"08",
          6422 => x"8a",
          6423 => x"54",
          6424 => x"82",
          6425 => x"55",
          6426 => x"08",
          6427 => x"82",
          6428 => x"52",
          6429 => x"e6",
          6430 => x"cc",
          6431 => x"87",
          6432 => x"38",
          6433 => x"cf",
          6434 => x"cc",
          6435 => x"88",
          6436 => x"cc",
          6437 => x"38",
          6438 => x"c3",
          6439 => x"cc",
          6440 => x"cc",
          6441 => x"82",
          6442 => x"07",
          6443 => x"55",
          6444 => x"2e",
          6445 => x"80",
          6446 => x"80",
          6447 => x"77",
          6448 => x"3f",
          6449 => x"08",
          6450 => x"38",
          6451 => x"ba",
          6452 => x"87",
          6453 => x"74",
          6454 => x"0c",
          6455 => x"04",
          6456 => x"82",
          6457 => x"c0",
          6458 => x"3d",
          6459 => x"3f",
          6460 => x"08",
          6461 => x"cc",
          6462 => x"38",
          6463 => x"52",
          6464 => x"52",
          6465 => x"3f",
          6466 => x"08",
          6467 => x"cc",
          6468 => x"88",
          6469 => x"39",
          6470 => x"08",
          6471 => x"81",
          6472 => x"38",
          6473 => x"05",
          6474 => x"2a",
          6475 => x"55",
          6476 => x"81",
          6477 => x"5a",
          6478 => x"3d",
          6479 => x"c1",
          6480 => x"87",
          6481 => x"55",
          6482 => x"cc",
          6483 => x"87",
          6484 => x"cc",
          6485 => x"09",
          6486 => x"38",
          6487 => x"87",
          6488 => x"2e",
          6489 => x"86",
          6490 => x"81",
          6491 => x"81",
          6492 => x"87",
          6493 => x"78",
          6494 => x"3f",
          6495 => x"08",
          6496 => x"cc",
          6497 => x"38",
          6498 => x"52",
          6499 => x"ff",
          6500 => x"78",
          6501 => x"b4",
          6502 => x"54",
          6503 => x"15",
          6504 => x"b2",
          6505 => x"ca",
          6506 => x"b6",
          6507 => x"53",
          6508 => x"53",
          6509 => x"3f",
          6510 => x"b4",
          6511 => x"d4",
          6512 => x"b6",
          6513 => x"54",
          6514 => x"d5",
          6515 => x"53",
          6516 => x"11",
          6517 => x"d8",
          6518 => x"81",
          6519 => x"34",
          6520 => x"a5",
          6521 => x"cc",
          6522 => x"87",
          6523 => x"38",
          6524 => x"0a",
          6525 => x"05",
          6526 => x"d1",
          6527 => x"64",
          6528 => x"c9",
          6529 => x"54",
          6530 => x"15",
          6531 => x"81",
          6532 => x"34",
          6533 => x"b8",
          6534 => x"87",
          6535 => x"8b",
          6536 => x"75",
          6537 => x"ff",
          6538 => x"73",
          6539 => x"0c",
          6540 => x"04",
          6541 => x"a9",
          6542 => x"51",
          6543 => x"82",
          6544 => x"ff",
          6545 => x"a9",
          6546 => x"ef",
          6547 => x"cc",
          6548 => x"87",
          6549 => x"d3",
          6550 => x"a9",
          6551 => x"9d",
          6552 => x"58",
          6553 => x"82",
          6554 => x"55",
          6555 => x"08",
          6556 => x"02",
          6557 => x"33",
          6558 => x"54",
          6559 => x"82",
          6560 => x"53",
          6561 => x"52",
          6562 => x"88",
          6563 => x"b4",
          6564 => x"53",
          6565 => x"3d",
          6566 => x"ff",
          6567 => x"aa",
          6568 => x"73",
          6569 => x"3f",
          6570 => x"08",
          6571 => x"cc",
          6572 => x"63",
          6573 => x"81",
          6574 => x"65",
          6575 => x"2e",
          6576 => x"55",
          6577 => x"82",
          6578 => x"84",
          6579 => x"06",
          6580 => x"73",
          6581 => x"3f",
          6582 => x"08",
          6583 => x"cc",
          6584 => x"38",
          6585 => x"53",
          6586 => x"95",
          6587 => x"16",
          6588 => x"88",
          6589 => x"05",
          6590 => x"34",
          6591 => x"70",
          6592 => x"81",
          6593 => x"55",
          6594 => x"74",
          6595 => x"73",
          6596 => x"78",
          6597 => x"83",
          6598 => x"16",
          6599 => x"2a",
          6600 => x"51",
          6601 => x"80",
          6602 => x"38",
          6603 => x"80",
          6604 => x"52",
          6605 => x"bf",
          6606 => x"cc",
          6607 => x"51",
          6608 => x"3f",
          6609 => x"87",
          6610 => x"2e",
          6611 => x"82",
          6612 => x"52",
          6613 => x"b5",
          6614 => x"87",
          6615 => x"80",
          6616 => x"58",
          6617 => x"cc",
          6618 => x"38",
          6619 => x"54",
          6620 => x"09",
          6621 => x"38",
          6622 => x"52",
          6623 => x"b0",
          6624 => x"81",
          6625 => x"34",
          6626 => x"87",
          6627 => x"38",
          6628 => x"cb",
          6629 => x"cc",
          6630 => x"87",
          6631 => x"38",
          6632 => x"b5",
          6633 => x"87",
          6634 => x"74",
          6635 => x"0c",
          6636 => x"04",
          6637 => x"02",
          6638 => x"33",
          6639 => x"80",
          6640 => x"57",
          6641 => x"95",
          6642 => x"52",
          6643 => x"d2",
          6644 => x"87",
          6645 => x"82",
          6646 => x"80",
          6647 => x"5a",
          6648 => x"3d",
          6649 => x"c9",
          6650 => x"87",
          6651 => x"82",
          6652 => x"b8",
          6653 => x"cf",
          6654 => x"a0",
          6655 => x"55",
          6656 => x"75",
          6657 => x"71",
          6658 => x"33",
          6659 => x"74",
          6660 => x"57",
          6661 => x"8b",
          6662 => x"54",
          6663 => x"15",
          6664 => x"ff",
          6665 => x"82",
          6666 => x"55",
          6667 => x"cc",
          6668 => x"0d",
          6669 => x"0d",
          6670 => x"53",
          6671 => x"05",
          6672 => x"51",
          6673 => x"82",
          6674 => x"55",
          6675 => x"08",
          6676 => x"76",
          6677 => x"93",
          6678 => x"51",
          6679 => x"82",
          6680 => x"55",
          6681 => x"08",
          6682 => x"80",
          6683 => x"81",
          6684 => x"86",
          6685 => x"38",
          6686 => x"86",
          6687 => x"90",
          6688 => x"54",
          6689 => x"ff",
          6690 => x"76",
          6691 => x"83",
          6692 => x"51",
          6693 => x"3f",
          6694 => x"08",
          6695 => x"87",
          6696 => x"3d",
          6697 => x"3d",
          6698 => x"5c",
          6699 => x"98",
          6700 => x"52",
          6701 => x"d1",
          6702 => x"87",
          6703 => x"87",
          6704 => x"70",
          6705 => x"08",
          6706 => x"51",
          6707 => x"80",
          6708 => x"38",
          6709 => x"06",
          6710 => x"80",
          6711 => x"38",
          6712 => x"5f",
          6713 => x"3d",
          6714 => x"ff",
          6715 => x"82",
          6716 => x"57",
          6717 => x"08",
          6718 => x"74",
          6719 => x"c3",
          6720 => x"87",
          6721 => x"82",
          6722 => x"bf",
          6723 => x"cc",
          6724 => x"cc",
          6725 => x"59",
          6726 => x"81",
          6727 => x"56",
          6728 => x"33",
          6729 => x"16",
          6730 => x"27",
          6731 => x"56",
          6732 => x"80",
          6733 => x"80",
          6734 => x"ff",
          6735 => x"70",
          6736 => x"56",
          6737 => x"e8",
          6738 => x"76",
          6739 => x"81",
          6740 => x"80",
          6741 => x"57",
          6742 => x"78",
          6743 => x"51",
          6744 => x"2e",
          6745 => x"73",
          6746 => x"38",
          6747 => x"08",
          6748 => x"b1",
          6749 => x"87",
          6750 => x"82",
          6751 => x"a7",
          6752 => x"33",
          6753 => x"c3",
          6754 => x"2e",
          6755 => x"e4",
          6756 => x"2e",
          6757 => x"56",
          6758 => x"05",
          6759 => x"e4",
          6760 => x"cc",
          6761 => x"76",
          6762 => x"0c",
          6763 => x"04",
          6764 => x"82",
          6765 => x"ff",
          6766 => x"9d",
          6767 => x"fb",
          6768 => x"cc",
          6769 => x"cc",
          6770 => x"82",
          6771 => x"83",
          6772 => x"53",
          6773 => x"3d",
          6774 => x"ff",
          6775 => x"73",
          6776 => x"70",
          6777 => x"52",
          6778 => x"9f",
          6779 => x"bc",
          6780 => x"74",
          6781 => x"6d",
          6782 => x"70",
          6783 => x"af",
          6784 => x"87",
          6785 => x"2e",
          6786 => x"70",
          6787 => x"57",
          6788 => x"fe",
          6789 => x"cc",
          6790 => x"8d",
          6791 => x"2b",
          6792 => x"81",
          6793 => x"86",
          6794 => x"cc",
          6795 => x"9f",
          6796 => x"ff",
          6797 => x"54",
          6798 => x"8a",
          6799 => x"70",
          6800 => x"06",
          6801 => x"ff",
          6802 => x"38",
          6803 => x"15",
          6804 => x"80",
          6805 => x"74",
          6806 => x"94",
          6807 => x"8a",
          6808 => x"cc",
          6809 => x"81",
          6810 => x"88",
          6811 => x"26",
          6812 => x"39",
          6813 => x"86",
          6814 => x"81",
          6815 => x"ff",
          6816 => x"38",
          6817 => x"54",
          6818 => x"81",
          6819 => x"81",
          6820 => x"78",
          6821 => x"5a",
          6822 => x"6d",
          6823 => x"81",
          6824 => x"57",
          6825 => x"9f",
          6826 => x"38",
          6827 => x"54",
          6828 => x"81",
          6829 => x"b1",
          6830 => x"2e",
          6831 => x"a7",
          6832 => x"15",
          6833 => x"54",
          6834 => x"09",
          6835 => x"38",
          6836 => x"76",
          6837 => x"41",
          6838 => x"52",
          6839 => x"52",
          6840 => x"b4",
          6841 => x"cc",
          6842 => x"87",
          6843 => x"f7",
          6844 => x"74",
          6845 => x"e6",
          6846 => x"cc",
          6847 => x"87",
          6848 => x"38",
          6849 => x"38",
          6850 => x"74",
          6851 => x"39",
          6852 => x"08",
          6853 => x"81",
          6854 => x"38",
          6855 => x"74",
          6856 => x"38",
          6857 => x"51",
          6858 => x"3f",
          6859 => x"08",
          6860 => x"cc",
          6861 => x"a0",
          6862 => x"cc",
          6863 => x"51",
          6864 => x"3f",
          6865 => x"0b",
          6866 => x"8b",
          6867 => x"67",
          6868 => x"a8",
          6869 => x"81",
          6870 => x"34",
          6871 => x"ad",
          6872 => x"87",
          6873 => x"73",
          6874 => x"87",
          6875 => x"3d",
          6876 => x"3d",
          6877 => x"02",
          6878 => x"cb",
          6879 => x"3d",
          6880 => x"72",
          6881 => x"5a",
          6882 => x"82",
          6883 => x"58",
          6884 => x"08",
          6885 => x"91",
          6886 => x"77",
          6887 => x"7c",
          6888 => x"38",
          6889 => x"59",
          6890 => x"90",
          6891 => x"81",
          6892 => x"06",
          6893 => x"73",
          6894 => x"54",
          6895 => x"82",
          6896 => x"39",
          6897 => x"8b",
          6898 => x"11",
          6899 => x"2b",
          6900 => x"54",
          6901 => x"ff",
          6902 => x"ff",
          6903 => x"70",
          6904 => x"07",
          6905 => x"87",
          6906 => x"8c",
          6907 => x"40",
          6908 => x"55",
          6909 => x"88",
          6910 => x"08",
          6911 => x"38",
          6912 => x"77",
          6913 => x"56",
          6914 => x"51",
          6915 => x"3f",
          6916 => x"55",
          6917 => x"08",
          6918 => x"38",
          6919 => x"87",
          6920 => x"2e",
          6921 => x"82",
          6922 => x"ff",
          6923 => x"38",
          6924 => x"08",
          6925 => x"16",
          6926 => x"2e",
          6927 => x"87",
          6928 => x"74",
          6929 => x"74",
          6930 => x"81",
          6931 => x"38",
          6932 => x"ff",
          6933 => x"2e",
          6934 => x"7b",
          6935 => x"80",
          6936 => x"81",
          6937 => x"81",
          6938 => x"06",
          6939 => x"56",
          6940 => x"52",
          6941 => x"af",
          6942 => x"87",
          6943 => x"82",
          6944 => x"80",
          6945 => x"81",
          6946 => x"56",
          6947 => x"d3",
          6948 => x"ff",
          6949 => x"7c",
          6950 => x"55",
          6951 => x"b3",
          6952 => x"1b",
          6953 => x"1b",
          6954 => x"33",
          6955 => x"54",
          6956 => x"34",
          6957 => x"fe",
          6958 => x"08",
          6959 => x"74",
          6960 => x"75",
          6961 => x"16",
          6962 => x"33",
          6963 => x"73",
          6964 => x"77",
          6965 => x"87",
          6966 => x"3d",
          6967 => x"3d",
          6968 => x"02",
          6969 => x"eb",
          6970 => x"3d",
          6971 => x"59",
          6972 => x"8b",
          6973 => x"82",
          6974 => x"24",
          6975 => x"82",
          6976 => x"84",
          6977 => x"f0",
          6978 => x"51",
          6979 => x"2e",
          6980 => x"75",
          6981 => x"cc",
          6982 => x"06",
          6983 => x"7e",
          6984 => x"d1",
          6985 => x"cc",
          6986 => x"06",
          6987 => x"56",
          6988 => x"74",
          6989 => x"76",
          6990 => x"81",
          6991 => x"8a",
          6992 => x"b2",
          6993 => x"fc",
          6994 => x"52",
          6995 => x"a4",
          6996 => x"87",
          6997 => x"38",
          6998 => x"80",
          6999 => x"74",
          7000 => x"26",
          7001 => x"15",
          7002 => x"74",
          7003 => x"38",
          7004 => x"80",
          7005 => x"84",
          7006 => x"92",
          7007 => x"80",
          7008 => x"38",
          7009 => x"06",
          7010 => x"2e",
          7011 => x"56",
          7012 => x"78",
          7013 => x"89",
          7014 => x"2b",
          7015 => x"43",
          7016 => x"38",
          7017 => x"30",
          7018 => x"77",
          7019 => x"91",
          7020 => x"c2",
          7021 => x"f8",
          7022 => x"52",
          7023 => x"a4",
          7024 => x"56",
          7025 => x"08",
          7026 => x"77",
          7027 => x"77",
          7028 => x"cc",
          7029 => x"45",
          7030 => x"bf",
          7031 => x"8e",
          7032 => x"26",
          7033 => x"74",
          7034 => x"48",
          7035 => x"75",
          7036 => x"38",
          7037 => x"81",
          7038 => x"fa",
          7039 => x"2a",
          7040 => x"56",
          7041 => x"2e",
          7042 => x"87",
          7043 => x"82",
          7044 => x"38",
          7045 => x"55",
          7046 => x"83",
          7047 => x"81",
          7048 => x"56",
          7049 => x"80",
          7050 => x"38",
          7051 => x"83",
          7052 => x"06",
          7053 => x"78",
          7054 => x"91",
          7055 => x"0b",
          7056 => x"22",
          7057 => x"80",
          7058 => x"74",
          7059 => x"38",
          7060 => x"56",
          7061 => x"17",
          7062 => x"57",
          7063 => x"2e",
          7064 => x"75",
          7065 => x"79",
          7066 => x"ff",
          7067 => x"82",
          7068 => x"84",
          7069 => x"05",
          7070 => x"5e",
          7071 => x"80",
          7072 => x"cc",
          7073 => x"8a",
          7074 => x"fd",
          7075 => x"75",
          7076 => x"38",
          7077 => x"78",
          7078 => x"8c",
          7079 => x"0b",
          7080 => x"22",
          7081 => x"80",
          7082 => x"74",
          7083 => x"38",
          7084 => x"56",
          7085 => x"17",
          7086 => x"57",
          7087 => x"2e",
          7088 => x"75",
          7089 => x"79",
          7090 => x"ff",
          7091 => x"82",
          7092 => x"10",
          7093 => x"82",
          7094 => x"9f",
          7095 => x"38",
          7096 => x"87",
          7097 => x"82",
          7098 => x"05",
          7099 => x"2a",
          7100 => x"56",
          7101 => x"17",
          7102 => x"81",
          7103 => x"60",
          7104 => x"65",
          7105 => x"12",
          7106 => x"30",
          7107 => x"74",
          7108 => x"59",
          7109 => x"7d",
          7110 => x"81",
          7111 => x"76",
          7112 => x"41",
          7113 => x"76",
          7114 => x"90",
          7115 => x"62",
          7116 => x"51",
          7117 => x"26",
          7118 => x"75",
          7119 => x"31",
          7120 => x"65",
          7121 => x"ff",
          7122 => x"82",
          7123 => x"58",
          7124 => x"09",
          7125 => x"38",
          7126 => x"08",
          7127 => x"26",
          7128 => x"78",
          7129 => x"79",
          7130 => x"78",
          7131 => x"86",
          7132 => x"82",
          7133 => x"06",
          7134 => x"83",
          7135 => x"82",
          7136 => x"27",
          7137 => x"8f",
          7138 => x"55",
          7139 => x"26",
          7140 => x"59",
          7141 => x"62",
          7142 => x"74",
          7143 => x"38",
          7144 => x"88",
          7145 => x"cc",
          7146 => x"26",
          7147 => x"86",
          7148 => x"1a",
          7149 => x"79",
          7150 => x"38",
          7151 => x"80",
          7152 => x"2e",
          7153 => x"83",
          7154 => x"9f",
          7155 => x"8b",
          7156 => x"06",
          7157 => x"74",
          7158 => x"84",
          7159 => x"52",
          7160 => x"a2",
          7161 => x"53",
          7162 => x"52",
          7163 => x"a2",
          7164 => x"80",
          7165 => x"51",
          7166 => x"3f",
          7167 => x"34",
          7168 => x"ff",
          7169 => x"1b",
          7170 => x"a3",
          7171 => x"90",
          7172 => x"83",
          7173 => x"70",
          7174 => x"80",
          7175 => x"55",
          7176 => x"ff",
          7177 => x"66",
          7178 => x"ff",
          7179 => x"38",
          7180 => x"ff",
          7181 => x"1b",
          7182 => x"f3",
          7183 => x"74",
          7184 => x"51",
          7185 => x"3f",
          7186 => x"1c",
          7187 => x"98",
          7188 => x"a0",
          7189 => x"ff",
          7190 => x"51",
          7191 => x"3f",
          7192 => x"1b",
          7193 => x"e5",
          7194 => x"2e",
          7195 => x"80",
          7196 => x"88",
          7197 => x"80",
          7198 => x"ff",
          7199 => x"7c",
          7200 => x"51",
          7201 => x"3f",
          7202 => x"1b",
          7203 => x"bd",
          7204 => x"b0",
          7205 => x"a0",
          7206 => x"52",
          7207 => x"ff",
          7208 => x"ff",
          7209 => x"c0",
          7210 => x"0b",
          7211 => x"34",
          7212 => x"80",
          7213 => x"c7",
          7214 => x"39",
          7215 => x"0a",
          7216 => x"51",
          7217 => x"3f",
          7218 => x"ff",
          7219 => x"1b",
          7220 => x"db",
          7221 => x"0b",
          7222 => x"a9",
          7223 => x"34",
          7224 => x"80",
          7225 => x"1b",
          7226 => x"90",
          7227 => x"d5",
          7228 => x"1b",
          7229 => x"ff",
          7230 => x"81",
          7231 => x"7a",
          7232 => x"ff",
          7233 => x"81",
          7234 => x"cc",
          7235 => x"38",
          7236 => x"09",
          7237 => x"ee",
          7238 => x"60",
          7239 => x"7a",
          7240 => x"ff",
          7241 => x"84",
          7242 => x"52",
          7243 => x"9f",
          7244 => x"8b",
          7245 => x"52",
          7246 => x"9f",
          7247 => x"8a",
          7248 => x"52",
          7249 => x"51",
          7250 => x"3f",
          7251 => x"83",
          7252 => x"ff",
          7253 => x"82",
          7254 => x"1b",
          7255 => x"ed",
          7256 => x"d5",
          7257 => x"ff",
          7258 => x"75",
          7259 => x"05",
          7260 => x"7e",
          7261 => x"e6",
          7262 => x"60",
          7263 => x"52",
          7264 => x"9a",
          7265 => x"53",
          7266 => x"51",
          7267 => x"3f",
          7268 => x"58",
          7269 => x"09",
          7270 => x"38",
          7271 => x"51",
          7272 => x"3f",
          7273 => x"1b",
          7274 => x"a1",
          7275 => x"52",
          7276 => x"91",
          7277 => x"ff",
          7278 => x"81",
          7279 => x"f8",
          7280 => x"7a",
          7281 => x"85",
          7282 => x"61",
          7283 => x"26",
          7284 => x"57",
          7285 => x"53",
          7286 => x"51",
          7287 => x"3f",
          7288 => x"08",
          7289 => x"84",
          7290 => x"87",
          7291 => x"7a",
          7292 => x"ab",
          7293 => x"75",
          7294 => x"56",
          7295 => x"81",
          7296 => x"80",
          7297 => x"38",
          7298 => x"83",
          7299 => x"63",
          7300 => x"74",
          7301 => x"38",
          7302 => x"54",
          7303 => x"52",
          7304 => x"99",
          7305 => x"87",
          7306 => x"c1",
          7307 => x"75",
          7308 => x"56",
          7309 => x"8c",
          7310 => x"2e",
          7311 => x"56",
          7312 => x"ff",
          7313 => x"84",
          7314 => x"2e",
          7315 => x"56",
          7316 => x"58",
          7317 => x"38",
          7318 => x"77",
          7319 => x"ff",
          7320 => x"82",
          7321 => x"78",
          7322 => x"c3",
          7323 => x"1b",
          7324 => x"34",
          7325 => x"16",
          7326 => x"82",
          7327 => x"83",
          7328 => x"84",
          7329 => x"67",
          7330 => x"fd",
          7331 => x"51",
          7332 => x"3f",
          7333 => x"16",
          7334 => x"cc",
          7335 => x"bf",
          7336 => x"86",
          7337 => x"87",
          7338 => x"16",
          7339 => x"83",
          7340 => x"ff",
          7341 => x"66",
          7342 => x"1b",
          7343 => x"8d",
          7344 => x"77",
          7345 => x"7e",
          7346 => x"92",
          7347 => x"82",
          7348 => x"a2",
          7349 => x"80",
          7350 => x"ff",
          7351 => x"81",
          7352 => x"cc",
          7353 => x"89",
          7354 => x"8a",
          7355 => x"86",
          7356 => x"cc",
          7357 => x"82",
          7358 => x"99",
          7359 => x"f5",
          7360 => x"60",
          7361 => x"79",
          7362 => x"5a",
          7363 => x"78",
          7364 => x"8d",
          7365 => x"55",
          7366 => x"fc",
          7367 => x"51",
          7368 => x"7a",
          7369 => x"81",
          7370 => x"8c",
          7371 => x"74",
          7372 => x"38",
          7373 => x"81",
          7374 => x"81",
          7375 => x"8a",
          7376 => x"06",
          7377 => x"76",
          7378 => x"76",
          7379 => x"55",
          7380 => x"cc",
          7381 => x"0d",
          7382 => x"0d",
          7383 => x"05",
          7384 => x"59",
          7385 => x"2e",
          7386 => x"87",
          7387 => x"76",
          7388 => x"84",
          7389 => x"80",
          7390 => x"38",
          7391 => x"77",
          7392 => x"56",
          7393 => x"34",
          7394 => x"bb",
          7395 => x"38",
          7396 => x"05",
          7397 => x"8c",
          7398 => x"08",
          7399 => x"3f",
          7400 => x"70",
          7401 => x"07",
          7402 => x"30",
          7403 => x"56",
          7404 => x"0c",
          7405 => x"18",
          7406 => x"0d",
          7407 => x"0d",
          7408 => x"08",
          7409 => x"75",
          7410 => x"89",
          7411 => x"54",
          7412 => x"16",
          7413 => x"51",
          7414 => x"82",
          7415 => x"91",
          7416 => x"08",
          7417 => x"81",
          7418 => x"88",
          7419 => x"83",
          7420 => x"74",
          7421 => x"0c",
          7422 => x"04",
          7423 => x"75",
          7424 => x"53",
          7425 => x"51",
          7426 => x"3f",
          7427 => x"85",
          7428 => x"ea",
          7429 => x"80",
          7430 => x"6a",
          7431 => x"70",
          7432 => x"d8",
          7433 => x"72",
          7434 => x"3f",
          7435 => x"8d",
          7436 => x"0d",
          7437 => x"ff",
          7438 => x"00",
          7439 => x"ff",
          7440 => x"ff",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"00",
          7471 => x"00",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"00",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"00",
          7480 => x"00",
          7481 => x"00",
          7482 => x"00",
          7483 => x"00",
          7484 => x"00",
          7485 => x"00",
          7486 => x"00",
          7487 => x"00",
          7488 => x"69",
          7489 => x"00",
          7490 => x"69",
          7491 => x"6c",
          7492 => x"69",
          7493 => x"00",
          7494 => x"6c",
          7495 => x"00",
          7496 => x"65",
          7497 => x"00",
          7498 => x"63",
          7499 => x"72",
          7500 => x"63",
          7501 => x"00",
          7502 => x"64",
          7503 => x"00",
          7504 => x"64",
          7505 => x"00",
          7506 => x"65",
          7507 => x"65",
          7508 => x"65",
          7509 => x"69",
          7510 => x"69",
          7511 => x"66",
          7512 => x"66",
          7513 => x"61",
          7514 => x"00",
          7515 => x"6d",
          7516 => x"65",
          7517 => x"72",
          7518 => x"65",
          7519 => x"00",
          7520 => x"6e",
          7521 => x"00",
          7522 => x"65",
          7523 => x"00",
          7524 => x"62",
          7525 => x"63",
          7526 => x"62",
          7527 => x"63",
          7528 => x"69",
          7529 => x"00",
          7530 => x"64",
          7531 => x"69",
          7532 => x"45",
          7533 => x"72",
          7534 => x"6e",
          7535 => x"6e",
          7536 => x"65",
          7537 => x"72",
          7538 => x"00",
          7539 => x"69",
          7540 => x"6e",
          7541 => x"72",
          7542 => x"79",
          7543 => x"00",
          7544 => x"6f",
          7545 => x"6c",
          7546 => x"6f",
          7547 => x"2e",
          7548 => x"6f",
          7549 => x"74",
          7550 => x"6f",
          7551 => x"2e",
          7552 => x"6e",
          7553 => x"69",
          7554 => x"69",
          7555 => x"61",
          7556 => x"0a",
          7557 => x"63",
          7558 => x"73",
          7559 => x"6e",
          7560 => x"2e",
          7561 => x"69",
          7562 => x"61",
          7563 => x"61",
          7564 => x"65",
          7565 => x"74",
          7566 => x"00",
          7567 => x"69",
          7568 => x"68",
          7569 => x"6c",
          7570 => x"6e",
          7571 => x"69",
          7572 => x"00",
          7573 => x"44",
          7574 => x"20",
          7575 => x"74",
          7576 => x"72",
          7577 => x"63",
          7578 => x"2e",
          7579 => x"72",
          7580 => x"20",
          7581 => x"62",
          7582 => x"69",
          7583 => x"6e",
          7584 => x"69",
          7585 => x"00",
          7586 => x"69",
          7587 => x"6e",
          7588 => x"65",
          7589 => x"6c",
          7590 => x"0a",
          7591 => x"6f",
          7592 => x"6d",
          7593 => x"69",
          7594 => x"20",
          7595 => x"65",
          7596 => x"74",
          7597 => x"66",
          7598 => x"64",
          7599 => x"20",
          7600 => x"6b",
          7601 => x"00",
          7602 => x"6f",
          7603 => x"74",
          7604 => x"6f",
          7605 => x"64",
          7606 => x"00",
          7607 => x"69",
          7608 => x"75",
          7609 => x"6f",
          7610 => x"61",
          7611 => x"6e",
          7612 => x"6e",
          7613 => x"6c",
          7614 => x"0a",
          7615 => x"69",
          7616 => x"69",
          7617 => x"6f",
          7618 => x"64",
          7619 => x"00",
          7620 => x"6e",
          7621 => x"66",
          7622 => x"65",
          7623 => x"6d",
          7624 => x"72",
          7625 => x"00",
          7626 => x"6f",
          7627 => x"61",
          7628 => x"6f",
          7629 => x"20",
          7630 => x"65",
          7631 => x"00",
          7632 => x"61",
          7633 => x"65",
          7634 => x"73",
          7635 => x"63",
          7636 => x"65",
          7637 => x"0a",
          7638 => x"75",
          7639 => x"73",
          7640 => x"00",
          7641 => x"6e",
          7642 => x"77",
          7643 => x"72",
          7644 => x"2e",
          7645 => x"25",
          7646 => x"62",
          7647 => x"73",
          7648 => x"20",
          7649 => x"25",
          7650 => x"62",
          7651 => x"73",
          7652 => x"63",
          7653 => x"00",
          7654 => x"65",
          7655 => x"00",
          7656 => x"30",
          7657 => x"00",
          7658 => x"20",
          7659 => x"30",
          7660 => x"00",
          7661 => x"20",
          7662 => x"20",
          7663 => x"00",
          7664 => x"30",
          7665 => x"00",
          7666 => x"20",
          7667 => x"7c",
          7668 => x"0d",
          7669 => x"50",
          7670 => x"00",
          7671 => x"2a",
          7672 => x"73",
          7673 => x"00",
          7674 => x"32",
          7675 => x"2f",
          7676 => x"30",
          7677 => x"31",
          7678 => x"00",
          7679 => x"5a",
          7680 => x"20",
          7681 => x"20",
          7682 => x"78",
          7683 => x"73",
          7684 => x"20",
          7685 => x"0a",
          7686 => x"50",
          7687 => x"20",
          7688 => x"65",
          7689 => x"70",
          7690 => x"61",
          7691 => x"65",
          7692 => x"00",
          7693 => x"69",
          7694 => x"20",
          7695 => x"65",
          7696 => x"70",
          7697 => x"00",
          7698 => x"53",
          7699 => x"6e",
          7700 => x"72",
          7701 => x"0a",
          7702 => x"4f",
          7703 => x"20",
          7704 => x"69",
          7705 => x"72",
          7706 => x"74",
          7707 => x"4f",
          7708 => x"20",
          7709 => x"69",
          7710 => x"72",
          7711 => x"74",
          7712 => x"41",
          7713 => x"20",
          7714 => x"69",
          7715 => x"72",
          7716 => x"74",
          7717 => x"41",
          7718 => x"20",
          7719 => x"69",
          7720 => x"72",
          7721 => x"74",
          7722 => x"41",
          7723 => x"20",
          7724 => x"69",
          7725 => x"72",
          7726 => x"74",
          7727 => x"41",
          7728 => x"20",
          7729 => x"69",
          7730 => x"72",
          7731 => x"74",
          7732 => x"65",
          7733 => x"6e",
          7734 => x"70",
          7735 => x"6d",
          7736 => x"2e",
          7737 => x"00",
          7738 => x"6e",
          7739 => x"69",
          7740 => x"74",
          7741 => x"72",
          7742 => x"0a",
          7743 => x"75",
          7744 => x"78",
          7745 => x"62",
          7746 => x"00",
          7747 => x"70",
          7748 => x"2e",
          7749 => x"00",
          7750 => x"3a",
          7751 => x"61",
          7752 => x"64",
          7753 => x"20",
          7754 => x"74",
          7755 => x"69",
          7756 => x"73",
          7757 => x"61",
          7758 => x"30",
          7759 => x"6c",
          7760 => x"65",
          7761 => x"69",
          7762 => x"61",
          7763 => x"6c",
          7764 => x"0a",
          7765 => x"20",
          7766 => x"61",
          7767 => x"69",
          7768 => x"69",
          7769 => x"00",
          7770 => x"6e",
          7771 => x"61",
          7772 => x"65",
          7773 => x"00",
          7774 => x"61",
          7775 => x"64",
          7776 => x"20",
          7777 => x"74",
          7778 => x"69",
          7779 => x"0a",
          7780 => x"63",
          7781 => x"0a",
          7782 => x"75",
          7783 => x"6c",
          7784 => x"69",
          7785 => x"2e",
          7786 => x"00",
          7787 => x"6f",
          7788 => x"6e",
          7789 => x"2e",
          7790 => x"6f",
          7791 => x"72",
          7792 => x"2e",
          7793 => x"00",
          7794 => x"30",
          7795 => x"28",
          7796 => x"78",
          7797 => x"25",
          7798 => x"78",
          7799 => x"38",
          7800 => x"00",
          7801 => x"75",
          7802 => x"4d",
          7803 => x"72",
          7804 => x"00",
          7805 => x"43",
          7806 => x"6c",
          7807 => x"2e",
          7808 => x"30",
          7809 => x"25",
          7810 => x"2d",
          7811 => x"3f",
          7812 => x"00",
          7813 => x"30",
          7814 => x"25",
          7815 => x"2d",
          7816 => x"30",
          7817 => x"25",
          7818 => x"2d",
          7819 => x"69",
          7820 => x"6c",
          7821 => x"20",
          7822 => x"65",
          7823 => x"70",
          7824 => x"00",
          7825 => x"6e",
          7826 => x"69",
          7827 => x"69",
          7828 => x"72",
          7829 => x"74",
          7830 => x"00",
          7831 => x"69",
          7832 => x"6c",
          7833 => x"75",
          7834 => x"20",
          7835 => x"6f",
          7836 => x"6e",
          7837 => x"69",
          7838 => x"75",
          7839 => x"20",
          7840 => x"6f",
          7841 => x"78",
          7842 => x"74",
          7843 => x"20",
          7844 => x"65",
          7845 => x"25",
          7846 => x"20",
          7847 => x"0a",
          7848 => x"61",
          7849 => x"6e",
          7850 => x"6f",
          7851 => x"40",
          7852 => x"38",
          7853 => x"2e",
          7854 => x"00",
          7855 => x"61",
          7856 => x"72",
          7857 => x"72",
          7858 => x"20",
          7859 => x"65",
          7860 => x"64",
          7861 => x"00",
          7862 => x"65",
          7863 => x"72",
          7864 => x"67",
          7865 => x"70",
          7866 => x"61",
          7867 => x"6e",
          7868 => x"0a",
          7869 => x"6f",
          7870 => x"72",
          7871 => x"6f",
          7872 => x"67",
          7873 => x"0a",
          7874 => x"50",
          7875 => x"69",
          7876 => x"64",
          7877 => x"73",
          7878 => x"2e",
          7879 => x"00",
          7880 => x"64",
          7881 => x"73",
          7882 => x"00",
          7883 => x"64",
          7884 => x"73",
          7885 => x"61",
          7886 => x"6f",
          7887 => x"6e",
          7888 => x"00",
          7889 => x"75",
          7890 => x"6e",
          7891 => x"2e",
          7892 => x"6e",
          7893 => x"69",
          7894 => x"69",
          7895 => x"72",
          7896 => x"74",
          7897 => x"2e",
          7898 => x"64",
          7899 => x"2f",
          7900 => x"25",
          7901 => x"64",
          7902 => x"2e",
          7903 => x"64",
          7904 => x"6f",
          7905 => x"6f",
          7906 => x"67",
          7907 => x"74",
          7908 => x"00",
          7909 => x"28",
          7910 => x"6d",
          7911 => x"43",
          7912 => x"6e",
          7913 => x"29",
          7914 => x"0a",
          7915 => x"69",
          7916 => x"20",
          7917 => x"6c",
          7918 => x"6e",
          7919 => x"3a",
          7920 => x"20",
          7921 => x"42",
          7922 => x"52",
          7923 => x"20",
          7924 => x"38",
          7925 => x"30",
          7926 => x"2e",
          7927 => x"20",
          7928 => x"44",
          7929 => x"20",
          7930 => x"20",
          7931 => x"38",
          7932 => x"30",
          7933 => x"2e",
          7934 => x"20",
          7935 => x"4e",
          7936 => x"42",
          7937 => x"20",
          7938 => x"38",
          7939 => x"30",
          7940 => x"2e",
          7941 => x"20",
          7942 => x"52",
          7943 => x"20",
          7944 => x"20",
          7945 => x"38",
          7946 => x"30",
          7947 => x"2e",
          7948 => x"20",
          7949 => x"41",
          7950 => x"20",
          7951 => x"20",
          7952 => x"38",
          7953 => x"30",
          7954 => x"2e",
          7955 => x"20",
          7956 => x"44",
          7957 => x"52",
          7958 => x"20",
          7959 => x"76",
          7960 => x"73",
          7961 => x"30",
          7962 => x"2e",
          7963 => x"20",
          7964 => x"49",
          7965 => x"31",
          7966 => x"20",
          7967 => x"6d",
          7968 => x"20",
          7969 => x"30",
          7970 => x"2e",
          7971 => x"20",
          7972 => x"4e",
          7973 => x"43",
          7974 => x"20",
          7975 => x"61",
          7976 => x"6c",
          7977 => x"30",
          7978 => x"2e",
          7979 => x"20",
          7980 => x"49",
          7981 => x"4f",
          7982 => x"42",
          7983 => x"00",
          7984 => x"20",
          7985 => x"42",
          7986 => x"43",
          7987 => x"20",
          7988 => x"4f",
          7989 => x"0a",
          7990 => x"20",
          7991 => x"53",
          7992 => x"00",
          7993 => x"20",
          7994 => x"50",
          7995 => x"00",
          7996 => x"64",
          7997 => x"73",
          7998 => x"3a",
          7999 => x"20",
          8000 => x"50",
          8001 => x"65",
          8002 => x"20",
          8003 => x"74",
          8004 => x"41",
          8005 => x"65",
          8006 => x"3d",
          8007 => x"38",
          8008 => x"00",
          8009 => x"20",
          8010 => x"50",
          8011 => x"65",
          8012 => x"79",
          8013 => x"61",
          8014 => x"41",
          8015 => x"65",
          8016 => x"3d",
          8017 => x"38",
          8018 => x"00",
          8019 => x"20",
          8020 => x"74",
          8021 => x"20",
          8022 => x"72",
          8023 => x"64",
          8024 => x"73",
          8025 => x"20",
          8026 => x"3d",
          8027 => x"38",
          8028 => x"00",
          8029 => x"69",
          8030 => x"0a",
          8031 => x"20",
          8032 => x"50",
          8033 => x"64",
          8034 => x"20",
          8035 => x"20",
          8036 => x"20",
          8037 => x"20",
          8038 => x"3d",
          8039 => x"34",
          8040 => x"00",
          8041 => x"20",
          8042 => x"79",
          8043 => x"6d",
          8044 => x"6f",
          8045 => x"46",
          8046 => x"20",
          8047 => x"20",
          8048 => x"3d",
          8049 => x"2e",
          8050 => x"64",
          8051 => x"0a",
          8052 => x"20",
          8053 => x"44",
          8054 => x"20",
          8055 => x"63",
          8056 => x"72",
          8057 => x"20",
          8058 => x"20",
          8059 => x"3d",
          8060 => x"2e",
          8061 => x"64",
          8062 => x"0a",
          8063 => x"20",
          8064 => x"69",
          8065 => x"6f",
          8066 => x"53",
          8067 => x"4d",
          8068 => x"6f",
          8069 => x"46",
          8070 => x"3d",
          8071 => x"2e",
          8072 => x"64",
          8073 => x"0a",
          8074 => x"6d",
          8075 => x"00",
          8076 => x"65",
          8077 => x"6d",
          8078 => x"6c",
          8079 => x"00",
          8080 => x"56",
          8081 => x"56",
          8082 => x"6e",
          8083 => x"6e",
          8084 => x"77",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"5b",
          8152 => x"5b",
          8153 => x"5b",
          8154 => x"5b",
          8155 => x"5b",
          8156 => x"5b",
          8157 => x"5b",
          8158 => x"30",
          8159 => x"5b",
          8160 => x"5b",
          8161 => x"5b",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"69",
          8174 => x"72",
          8175 => x"69",
          8176 => x"00",
          8177 => x"00",
          8178 => x"30",
          8179 => x"20",
          8180 => x"00",
          8181 => x"61",
          8182 => x"64",
          8183 => x"20",
          8184 => x"65",
          8185 => x"68",
          8186 => x"69",
          8187 => x"72",
          8188 => x"69",
          8189 => x"74",
          8190 => x"4f",
          8191 => x"00",
          8192 => x"61",
          8193 => x"74",
          8194 => x"65",
          8195 => x"72",
          8196 => x"65",
          8197 => x"73",
          8198 => x"79",
          8199 => x"6c",
          8200 => x"64",
          8201 => x"62",
          8202 => x"67",
          8203 => x"00",
          8204 => x"44",
          8205 => x"2a",
          8206 => x"3b",
          8207 => x"3f",
          8208 => x"7f",
          8209 => x"41",
          8210 => x"41",
          8211 => x"00",
          8212 => x"fe",
          8213 => x"44",
          8214 => x"2e",
          8215 => x"4f",
          8216 => x"4d",
          8217 => x"20",
          8218 => x"54",
          8219 => x"20",
          8220 => x"4f",
          8221 => x"4d",
          8222 => x"20",
          8223 => x"54",
          8224 => x"20",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"9a",
          8230 => x"41",
          8231 => x"45",
          8232 => x"49",
          8233 => x"92",
          8234 => x"4f",
          8235 => x"99",
          8236 => x"9d",
          8237 => x"49",
          8238 => x"a5",
          8239 => x"a9",
          8240 => x"ad",
          8241 => x"b1",
          8242 => x"b5",
          8243 => x"b9",
          8244 => x"bd",
          8245 => x"c1",
          8246 => x"c5",
          8247 => x"c9",
          8248 => x"cd",
          8249 => x"d1",
          8250 => x"d5",
          8251 => x"d9",
          8252 => x"dd",
          8253 => x"e1",
          8254 => x"e5",
          8255 => x"e9",
          8256 => x"ed",
          8257 => x"f1",
          8258 => x"f5",
          8259 => x"f9",
          8260 => x"fd",
          8261 => x"2e",
          8262 => x"5b",
          8263 => x"22",
          8264 => x"3e",
          8265 => x"00",
          8266 => x"01",
          8267 => x"10",
          8268 => x"00",
          8269 => x"00",
          8270 => x"01",
          8271 => x"04",
          8272 => x"10",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"02",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"04",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"14",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"2b",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"30",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"3c",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"3d",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"3f",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"40",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"41",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"42",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"43",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"50",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"51",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"54",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"55",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"79",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"78",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"82",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"83",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"85",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"87",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"8c",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"8d",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"8e",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"8f",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"01",
          8385 => x"00",
          8386 => x"01",
          8387 => x"81",
          8388 => x"00",
          8389 => x"7f",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"f5",
          8395 => x"f5",
          8396 => x"f5",
          8397 => x"00",
          8398 => x"01",
          8399 => x"01",
          8400 => x"01",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"99",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"fd",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"b4",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"b6",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"f2",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b4",
           272 => x"0b",
           273 => x"0b",
           274 => x"d4",
           275 => x"0b",
           276 => x"0b",
           277 => x"f4",
           278 => x"0b",
           279 => x"0b",
           280 => x"94",
           281 => x"0b",
           282 => x"0b",
           283 => x"b4",
           284 => x"0b",
           285 => x"0b",
           286 => x"d4",
           287 => x"0b",
           288 => x"0b",
           289 => x"f4",
           290 => x"0b",
           291 => x"0b",
           292 => x"92",
           293 => x"0b",
           294 => x"0b",
           295 => x"b1",
           296 => x"0b",
           297 => x"0b",
           298 => x"d1",
           299 => x"0b",
           300 => x"0b",
           301 => x"f1",
           302 => x"0b",
           303 => x"0b",
           304 => x"91",
           305 => x"0b",
           306 => x"0b",
           307 => x"b1",
           308 => x"0b",
           309 => x"0b",
           310 => x"d1",
           311 => x"0b",
           312 => x"0b",
           313 => x"f1",
           314 => x"0b",
           315 => x"0b",
           316 => x"91",
           317 => x"0b",
           318 => x"0b",
           319 => x"b1",
           320 => x"0b",
           321 => x"0b",
           322 => x"d1",
           323 => x"0b",
           324 => x"0b",
           325 => x"f1",
           326 => x"0b",
           327 => x"0b",
           328 => x"91",
           329 => x"0b",
           330 => x"0b",
           331 => x"b1",
           332 => x"0b",
           333 => x"0b",
           334 => x"d1",
           335 => x"0b",
           336 => x"0b",
           337 => x"f1",
           338 => x"0b",
           339 => x"0b",
           340 => x"90",
           341 => x"0b",
           342 => x"0b",
           343 => x"ae",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"80",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"80",
           395 => x"82",
           396 => x"82",
           397 => x"82",
           398 => x"80",
           399 => x"82",
           400 => x"82",
           401 => x"82",
           402 => x"80",
           403 => x"82",
           404 => x"82",
           405 => x"82",
           406 => x"80",
           407 => x"82",
           408 => x"82",
           409 => x"82",
           410 => x"80",
           411 => x"82",
           412 => x"82",
           413 => x"82",
           414 => x"80",
           415 => x"82",
           416 => x"82",
           417 => x"82",
           418 => x"80",
           419 => x"82",
           420 => x"82",
           421 => x"82",
           422 => x"80",
           423 => x"82",
           424 => x"82",
           425 => x"82",
           426 => x"80",
           427 => x"82",
           428 => x"82",
           429 => x"82",
           430 => x"80",
           431 => x"82",
           432 => x"82",
           433 => x"82",
           434 => x"80",
           435 => x"82",
           436 => x"82",
           437 => x"82",
           438 => x"80",
           439 => x"82",
           440 => x"82",
           441 => x"82",
           442 => x"80",
           443 => x"82",
           444 => x"82",
           445 => x"82",
           446 => x"b8",
           447 => x"87",
           448 => x"a0",
           449 => x"87",
           450 => x"ca",
           451 => x"d8",
           452 => x"90",
           453 => x"d8",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"04",
           565 => x"0c",
           566 => x"2d",
           567 => x"08",
           568 => x"04",
           569 => x"0c",
           570 => x"2d",
           571 => x"08",
           572 => x"04",
           573 => x"0c",
           574 => x"2d",
           575 => x"08",
           576 => x"04",
           577 => x"0c",
           578 => x"82",
           579 => x"82",
           580 => x"82",
           581 => x"ba",
           582 => x"87",
           583 => x"a0",
           584 => x"87",
           585 => x"8d",
           586 => x"d8",
           587 => x"90",
           588 => x"d8",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"00",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"53",
           601 => x"00",
           602 => x"06",
           603 => x"09",
           604 => x"05",
           605 => x"2b",
           606 => x"06",
           607 => x"04",
           608 => x"72",
           609 => x"05",
           610 => x"05",
           611 => x"72",
           612 => x"53",
           613 => x"51",
           614 => x"04",
           615 => x"70",
           616 => x"27",
           617 => x"71",
           618 => x"53",
           619 => x"0b",
           620 => x"8c",
           621 => x"ad",
           622 => x"87",
           623 => x"82",
           624 => x"fe",
           625 => x"87",
           626 => x"05",
           627 => x"d8",
           628 => x"0c",
           629 => x"08",
           630 => x"52",
           631 => x"87",
           632 => x"05",
           633 => x"82",
           634 => x"fc",
           635 => x"81",
           636 => x"51",
           637 => x"83",
           638 => x"82",
           639 => x"fc",
           640 => x"05",
           641 => x"08",
           642 => x"82",
           643 => x"fc",
           644 => x"87",
           645 => x"05",
           646 => x"82",
           647 => x"51",
           648 => x"82",
           649 => x"04",
           650 => x"08",
           651 => x"d8",
           652 => x"0d",
           653 => x"08",
           654 => x"82",
           655 => x"fc",
           656 => x"87",
           657 => x"05",
           658 => x"33",
           659 => x"08",
           660 => x"81",
           661 => x"d8",
           662 => x"0c",
           663 => x"08",
           664 => x"53",
           665 => x"34",
           666 => x"08",
           667 => x"81",
           668 => x"d8",
           669 => x"0c",
           670 => x"06",
           671 => x"2e",
           672 => x"be",
           673 => x"d8",
           674 => x"08",
           675 => x"cc",
           676 => x"3d",
           677 => x"d8",
           678 => x"87",
           679 => x"82",
           680 => x"fd",
           681 => x"87",
           682 => x"05",
           683 => x"d8",
           684 => x"0c",
           685 => x"08",
           686 => x"82",
           687 => x"f8",
           688 => x"87",
           689 => x"05",
           690 => x"80",
           691 => x"87",
           692 => x"05",
           693 => x"82",
           694 => x"90",
           695 => x"87",
           696 => x"05",
           697 => x"82",
           698 => x"90",
           699 => x"87",
           700 => x"05",
           701 => x"ba",
           702 => x"d8",
           703 => x"08",
           704 => x"82",
           705 => x"f8",
           706 => x"05",
           707 => x"08",
           708 => x"82",
           709 => x"fc",
           710 => x"52",
           711 => x"82",
           712 => x"fc",
           713 => x"05",
           714 => x"08",
           715 => x"ff",
           716 => x"87",
           717 => x"05",
           718 => x"87",
           719 => x"85",
           720 => x"87",
           721 => x"82",
           722 => x"02",
           723 => x"0c",
           724 => x"82",
           725 => x"90",
           726 => x"2e",
           727 => x"82",
           728 => x"8c",
           729 => x"71",
           730 => x"d8",
           731 => x"08",
           732 => x"87",
           733 => x"05",
           734 => x"d8",
           735 => x"08",
           736 => x"81",
           737 => x"54",
           738 => x"71",
           739 => x"80",
           740 => x"87",
           741 => x"05",
           742 => x"33",
           743 => x"08",
           744 => x"81",
           745 => x"d8",
           746 => x"0c",
           747 => x"06",
           748 => x"8d",
           749 => x"82",
           750 => x"fc",
           751 => x"9b",
           752 => x"d8",
           753 => x"08",
           754 => x"87",
           755 => x"05",
           756 => x"d8",
           757 => x"08",
           758 => x"38",
           759 => x"82",
           760 => x"90",
           761 => x"2e",
           762 => x"82",
           763 => x"88",
           764 => x"33",
           765 => x"8d",
           766 => x"82",
           767 => x"fc",
           768 => x"d7",
           769 => x"d8",
           770 => x"08",
           771 => x"87",
           772 => x"05",
           773 => x"d8",
           774 => x"08",
           775 => x"52",
           776 => x"81",
           777 => x"d8",
           778 => x"0c",
           779 => x"87",
           780 => x"05",
           781 => x"82",
           782 => x"8c",
           783 => x"33",
           784 => x"70",
           785 => x"08",
           786 => x"53",
           787 => x"53",
           788 => x"0b",
           789 => x"08",
           790 => x"82",
           791 => x"fc",
           792 => x"87",
           793 => x"3d",
           794 => x"d8",
           795 => x"87",
           796 => x"82",
           797 => x"fe",
           798 => x"87",
           799 => x"05",
           800 => x"d8",
           801 => x"0c",
           802 => x"08",
           803 => x"80",
           804 => x"38",
           805 => x"08",
           806 => x"81",
           807 => x"d8",
           808 => x"0c",
           809 => x"08",
           810 => x"ff",
           811 => x"d8",
           812 => x"0c",
           813 => x"08",
           814 => x"80",
           815 => x"82",
           816 => x"8c",
           817 => x"70",
           818 => x"08",
           819 => x"52",
           820 => x"34",
           821 => x"08",
           822 => x"81",
           823 => x"d8",
           824 => x"0c",
           825 => x"82",
           826 => x"88",
           827 => x"82",
           828 => x"51",
           829 => x"82",
           830 => x"04",
           831 => x"79",
           832 => x"56",
           833 => x"80",
           834 => x"38",
           835 => x"08",
           836 => x"3f",
           837 => x"08",
           838 => x"85",
           839 => x"80",
           840 => x"33",
           841 => x"2e",
           842 => x"86",
           843 => x"55",
           844 => x"57",
           845 => x"82",
           846 => x"70",
           847 => x"f8",
           848 => x"87",
           849 => x"74",
           850 => x"51",
           851 => x"82",
           852 => x"8b",
           853 => x"33",
           854 => x"2e",
           855 => x"81",
           856 => x"ff",
           857 => x"99",
           858 => x"38",
           859 => x"82",
           860 => x"89",
           861 => x"ff",
           862 => x"52",
           863 => x"81",
           864 => x"84",
           865 => x"c4",
           866 => x"08",
           867 => x"ac",
           868 => x"39",
           869 => x"51",
           870 => x"81",
           871 => x"80",
           872 => x"eb",
           873 => x"eb",
           874 => x"f0",
           875 => x"39",
           876 => x"51",
           877 => x"81",
           878 => x"80",
           879 => x"ec",
           880 => x"cf",
           881 => x"bc",
           882 => x"39",
           883 => x"51",
           884 => x"81",
           885 => x"bb",
           886 => x"88",
           887 => x"81",
           888 => x"af",
           889 => x"c8",
           890 => x"81",
           891 => x"a3",
           892 => x"fc",
           893 => x"81",
           894 => x"97",
           895 => x"a8",
           896 => x"81",
           897 => x"8b",
           898 => x"d8",
           899 => x"81",
           900 => x"b0",
           901 => x"3d",
           902 => x"3d",
           903 => x"56",
           904 => x"e7",
           905 => x"74",
           906 => x"e8",
           907 => x"39",
           908 => x"74",
           909 => x"b6",
           910 => x"cc",
           911 => x"51",
           912 => x"3f",
           913 => x"08",
           914 => x"75",
           915 => x"f4",
           916 => x"3f",
           917 => x"04",
           918 => x"66",
           919 => x"80",
           920 => x"5b",
           921 => x"78",
           922 => x"07",
           923 => x"57",
           924 => x"56",
           925 => x"26",
           926 => x"56",
           927 => x"70",
           928 => x"51",
           929 => x"74",
           930 => x"81",
           931 => x"8c",
           932 => x"56",
           933 => x"3f",
           934 => x"08",
           935 => x"cc",
           936 => x"82",
           937 => x"87",
           938 => x"0c",
           939 => x"08",
           940 => x"d4",
           941 => x"80",
           942 => x"75",
           943 => x"bf",
           944 => x"cc",
           945 => x"87",
           946 => x"38",
           947 => x"80",
           948 => x"74",
           949 => x"59",
           950 => x"96",
           951 => x"51",
           952 => x"3f",
           953 => x"78",
           954 => x"7b",
           955 => x"2a",
           956 => x"57",
           957 => x"80",
           958 => x"81",
           959 => x"87",
           960 => x"08",
           961 => x"fe",
           962 => x"56",
           963 => x"cc",
           964 => x"0d",
           965 => x"0d",
           966 => x"05",
           967 => x"57",
           968 => x"80",
           969 => x"79",
           970 => x"3f",
           971 => x"08",
           972 => x"80",
           973 => x"75",
           974 => x"38",
           975 => x"55",
           976 => x"87",
           977 => x"52",
           978 => x"2d",
           979 => x"08",
           980 => x"77",
           981 => x"87",
           982 => x"3d",
           983 => x"3d",
           984 => x"63",
           985 => x"80",
           986 => x"73",
           987 => x"41",
           988 => x"5e",
           989 => x"52",
           990 => x"51",
           991 => x"81",
           992 => x"ad",
           993 => x"55",
           994 => x"80",
           995 => x"90",
           996 => x"7b",
           997 => x"38",
           998 => x"74",
           999 => x"7a",
          1000 => x"72",
          1001 => x"ef",
          1002 => x"db",
          1003 => x"81",
          1004 => x"ac",
          1005 => x"15",
          1006 => x"74",
          1007 => x"7a",
          1008 => x"72",
          1009 => x"ef",
          1010 => x"bb",
          1011 => x"81",
          1012 => x"ac",
          1013 => x"15",
          1014 => x"74",
          1015 => x"7a",
          1016 => x"72",
          1017 => x"ef",
          1018 => x"9b",
          1019 => x"81",
          1020 => x"ac",
          1021 => x"15",
          1022 => x"ab",
          1023 => x"88",
          1024 => x"cc",
          1025 => x"3f",
          1026 => x"79",
          1027 => x"74",
          1028 => x"55",
          1029 => x"72",
          1030 => x"38",
          1031 => x"53",
          1032 => x"83",
          1033 => x"75",
          1034 => x"81",
          1035 => x"53",
          1036 => x"8b",
          1037 => x"fe",
          1038 => x"73",
          1039 => x"a0",
          1040 => x"3f",
          1041 => x"c2",
          1042 => x"d0",
          1043 => x"3f",
          1044 => x"1c",
          1045 => x"9a",
          1046 => x"cc",
          1047 => x"70",
          1048 => x"57",
          1049 => x"09",
          1050 => x"38",
          1051 => x"82",
          1052 => x"98",
          1053 => x"2c",
          1054 => x"70",
          1055 => x"32",
          1056 => x"72",
          1057 => x"07",
          1058 => x"58",
          1059 => x"57",
          1060 => x"d8",
          1061 => x"2e",
          1062 => x"85",
          1063 => x"8c",
          1064 => x"53",
          1065 => x"fd",
          1066 => x"53",
          1067 => x"cc",
          1068 => x"0d",
          1069 => x"0d",
          1070 => x"33",
          1071 => x"53",
          1072 => x"52",
          1073 => x"3f",
          1074 => x"22",
          1075 => x"3f",
          1076 => x"54",
          1077 => x"53",
          1078 => x"33",
          1079 => x"fc",
          1080 => x"3f",
          1081 => x"84",
          1082 => x"3f",
          1083 => x"04",
          1084 => x"87",
          1085 => x"08",
          1086 => x"3f",
          1087 => x"90",
          1088 => x"98",
          1089 => x"3f",
          1090 => x"84",
          1091 => x"2a",
          1092 => x"51",
          1093 => x"2e",
          1094 => x"51",
          1095 => x"81",
          1096 => x"9c",
          1097 => x"51",
          1098 => x"72",
          1099 => x"81",
          1100 => x"71",
          1101 => x"38",
          1102 => x"d4",
          1103 => x"c8",
          1104 => x"3f",
          1105 => x"c8",
          1106 => x"2a",
          1107 => x"51",
          1108 => x"2e",
          1109 => x"51",
          1110 => x"81",
          1111 => x"9c",
          1112 => x"51",
          1113 => x"72",
          1114 => x"81",
          1115 => x"71",
          1116 => x"38",
          1117 => x"98",
          1118 => x"ec",
          1119 => x"3f",
          1120 => x"8c",
          1121 => x"2a",
          1122 => x"51",
          1123 => x"2e",
          1124 => x"51",
          1125 => x"81",
          1126 => x"9b",
          1127 => x"51",
          1128 => x"72",
          1129 => x"81",
          1130 => x"71",
          1131 => x"38",
          1132 => x"dc",
          1133 => x"94",
          1134 => x"3f",
          1135 => x"d0",
          1136 => x"2a",
          1137 => x"51",
          1138 => x"2e",
          1139 => x"51",
          1140 => x"81",
          1141 => x"9b",
          1142 => x"51",
          1143 => x"72",
          1144 => x"81",
          1145 => x"71",
          1146 => x"38",
          1147 => x"a0",
          1148 => x"bc",
          1149 => x"3f",
          1150 => x"94",
          1151 => x"3f",
          1152 => x"04",
          1153 => x"77",
          1154 => x"a3",
          1155 => x"55",
          1156 => x"52",
          1157 => x"d6",
          1158 => x"82",
          1159 => x"54",
          1160 => x"81",
          1161 => x"fc",
          1162 => x"ac",
          1163 => x"ea",
          1164 => x"cc",
          1165 => x"82",
          1166 => x"07",
          1167 => x"71",
          1168 => x"54",
          1169 => x"82",
          1170 => x"0b",
          1171 => x"c8",
          1172 => x"81",
          1173 => x"06",
          1174 => x"9e",
          1175 => x"52",
          1176 => x"c1",
          1177 => x"87",
          1178 => x"2e",
          1179 => x"87",
          1180 => x"a7",
          1181 => x"39",
          1182 => x"51",
          1183 => x"3f",
          1184 => x"0b",
          1185 => x"34",
          1186 => x"82",
          1187 => x"73",
          1188 => x"81",
          1189 => x"81",
          1190 => x"74",
          1191 => x"b9",
          1192 => x"0b",
          1193 => x"0c",
          1194 => x"04",
          1195 => x"80",
          1196 => x"9e",
          1197 => x"5d",
          1198 => x"51",
          1199 => x"3f",
          1200 => x"08",
          1201 => x"59",
          1202 => x"09",
          1203 => x"38",
          1204 => x"52",
          1205 => x"52",
          1206 => x"3f",
          1207 => x"52",
          1208 => x"51",
          1209 => x"3f",
          1210 => x"08",
          1211 => x"38",
          1212 => x"51",
          1213 => x"81",
          1214 => x"81",
          1215 => x"a6",
          1216 => x"3d",
          1217 => x"80",
          1218 => x"51",
          1219 => x"b4",
          1220 => x"05",
          1221 => x"3f",
          1222 => x"08",
          1223 => x"90",
          1224 => x"78",
          1225 => x"89",
          1226 => x"80",
          1227 => x"d9",
          1228 => x"2e",
          1229 => x"78",
          1230 => x"38",
          1231 => x"81",
          1232 => x"82",
          1233 => x"78",
          1234 => x"af",
          1235 => x"39",
          1236 => x"82",
          1237 => x"94",
          1238 => x"38",
          1239 => x"78",
          1240 => x"fa",
          1241 => x"24",
          1242 => x"b0",
          1243 => x"38",
          1244 => x"84",
          1245 => x"b8",
          1246 => x"2e",
          1247 => x"78",
          1248 => x"86",
          1249 => x"a8",
          1250 => x"d5",
          1251 => x"38",
          1252 => x"24",
          1253 => x"80",
          1254 => x"c1",
          1255 => x"d0",
          1256 => x"78",
          1257 => x"89",
          1258 => x"80",
          1259 => x"94",
          1260 => x"39",
          1261 => x"2e",
          1262 => x"78",
          1263 => x"8c",
          1264 => x"ec",
          1265 => x"82",
          1266 => x"38",
          1267 => x"24",
          1268 => x"80",
          1269 => x"db",
          1270 => x"f9",
          1271 => x"38",
          1272 => x"78",
          1273 => x"8d",
          1274 => x"81",
          1275 => x"ba",
          1276 => x"39",
          1277 => x"80",
          1278 => x"84",
          1279 => x"fc",
          1280 => x"cc",
          1281 => x"81",
          1282 => x"8f",
          1283 => x"3d",
          1284 => x"53",
          1285 => x"51",
          1286 => x"82",
          1287 => x"80",
          1288 => x"81",
          1289 => x"38",
          1290 => x"80",
          1291 => x"52",
          1292 => x"05",
          1293 => x"d2",
          1294 => x"87",
          1295 => x"ff",
          1296 => x"8d",
          1297 => x"e8",
          1298 => x"3f",
          1299 => x"ab",
          1300 => x"f8",
          1301 => x"39",
          1302 => x"80",
          1303 => x"84",
          1304 => x"98",
          1305 => x"cc",
          1306 => x"fd",
          1307 => x"53",
          1308 => x"80",
          1309 => x"51",
          1310 => x"3f",
          1311 => x"08",
          1312 => x"90",
          1313 => x"39",
          1314 => x"80",
          1315 => x"84",
          1316 => x"e8",
          1317 => x"cc",
          1318 => x"87",
          1319 => x"26",
          1320 => x"b4",
          1321 => x"11",
          1322 => x"05",
          1323 => x"3f",
          1324 => x"08",
          1325 => x"87",
          1326 => x"63",
          1327 => x"98",
          1328 => x"a8",
          1329 => x"80",
          1330 => x"53",
          1331 => x"84",
          1332 => x"88",
          1333 => x"81",
          1334 => x"82",
          1335 => x"81",
          1336 => x"f2",
          1337 => x"bb",
          1338 => x"fc",
          1339 => x"3d",
          1340 => x"51",
          1341 => x"82",
          1342 => x"b5",
          1343 => x"05",
          1344 => x"9f",
          1345 => x"82",
          1346 => x"52",
          1347 => x"c8",
          1348 => x"39",
          1349 => x"84",
          1350 => x"e3",
          1351 => x"cc",
          1352 => x"ff",
          1353 => x"5b",
          1354 => x"82",
          1355 => x"b5",
          1356 => x"05",
          1357 => x"eb",
          1358 => x"cc",
          1359 => x"ff",
          1360 => x"59",
          1361 => x"82",
          1362 => x"82",
          1363 => x"80",
          1364 => x"82",
          1365 => x"81",
          1366 => x"78",
          1367 => x"7a",
          1368 => x"3f",
          1369 => x"08",
          1370 => x"8f",
          1371 => x"cc",
          1372 => x"83",
          1373 => x"39",
          1374 => x"80",
          1375 => x"84",
          1376 => x"f8",
          1377 => x"cc",
          1378 => x"fa",
          1379 => x"3d",
          1380 => x"53",
          1381 => x"51",
          1382 => x"82",
          1383 => x"80",
          1384 => x"38",
          1385 => x"f8",
          1386 => x"84",
          1387 => x"cc",
          1388 => x"cc",
          1389 => x"82",
          1390 => x"42",
          1391 => x"51",
          1392 => x"63",
          1393 => x"79",
          1394 => x"e9",
          1395 => x"78",
          1396 => x"05",
          1397 => x"7a",
          1398 => x"81",
          1399 => x"3d",
          1400 => x"53",
          1401 => x"51",
          1402 => x"82",
          1403 => x"80",
          1404 => x"38",
          1405 => x"fc",
          1406 => x"84",
          1407 => x"fc",
          1408 => x"cc",
          1409 => x"f9",
          1410 => x"3d",
          1411 => x"53",
          1412 => x"51",
          1413 => x"82",
          1414 => x"80",
          1415 => x"38",
          1416 => x"51",
          1417 => x"63",
          1418 => x"27",
          1419 => x"61",
          1420 => x"81",
          1421 => x"79",
          1422 => x"05",
          1423 => x"b4",
          1424 => x"11",
          1425 => x"05",
          1426 => x"3f",
          1427 => x"08",
          1428 => x"a7",
          1429 => x"fe",
          1430 => x"ff",
          1431 => x"a7",
          1432 => x"87",
          1433 => x"2e",
          1434 => x"b4",
          1435 => x"11",
          1436 => x"05",
          1437 => x"3f",
          1438 => x"08",
          1439 => x"fb",
          1440 => x"b8",
          1441 => x"3f",
          1442 => x"63",
          1443 => x"61",
          1444 => x"33",
          1445 => x"78",
          1446 => x"38",
          1447 => x"54",
          1448 => x"79",
          1449 => x"c8",
          1450 => x"3f",
          1451 => x"81",
          1452 => x"d6",
          1453 => x"e4",
          1454 => x"39",
          1455 => x"80",
          1456 => x"84",
          1457 => x"b4",
          1458 => x"cc",
          1459 => x"38",
          1460 => x"33",
          1461 => x"2e",
          1462 => x"85",
          1463 => x"80",
          1464 => x"86",
          1465 => x"78",
          1466 => x"38",
          1467 => x"08",
          1468 => x"82",
          1469 => x"59",
          1470 => x"88",
          1471 => x"80",
          1472 => x"39",
          1473 => x"33",
          1474 => x"2e",
          1475 => x"86",
          1476 => x"9a",
          1477 => x"b6",
          1478 => x"80",
          1479 => x"82",
          1480 => x"44",
          1481 => x"86",
          1482 => x"80",
          1483 => x"3d",
          1484 => x"53",
          1485 => x"51",
          1486 => x"82",
          1487 => x"80",
          1488 => x"86",
          1489 => x"78",
          1490 => x"38",
          1491 => x"08",
          1492 => x"39",
          1493 => x"33",
          1494 => x"2e",
          1495 => x"85",
          1496 => x"bb",
          1497 => x"ba",
          1498 => x"80",
          1499 => x"82",
          1500 => x"43",
          1501 => x"86",
          1502 => x"78",
          1503 => x"38",
          1504 => x"08",
          1505 => x"82",
          1506 => x"59",
          1507 => x"88",
          1508 => x"94",
          1509 => x"39",
          1510 => x"08",
          1511 => x"b4",
          1512 => x"11",
          1513 => x"05",
          1514 => x"3f",
          1515 => x"08",
          1516 => x"38",
          1517 => x"5c",
          1518 => x"83",
          1519 => x"7a",
          1520 => x"30",
          1521 => x"9f",
          1522 => x"06",
          1523 => x"5a",
          1524 => x"88",
          1525 => x"2e",
          1526 => x"42",
          1527 => x"51",
          1528 => x"a0",
          1529 => x"61",
          1530 => x"63",
          1531 => x"3f",
          1532 => x"51",
          1533 => x"f6",
          1534 => x"3d",
          1535 => x"53",
          1536 => x"51",
          1537 => x"82",
          1538 => x"80",
          1539 => x"38",
          1540 => x"fc",
          1541 => x"84",
          1542 => x"e0",
          1543 => x"cc",
          1544 => x"a4",
          1545 => x"02",
          1546 => x"33",
          1547 => x"81",
          1548 => x"3d",
          1549 => x"53",
          1550 => x"51",
          1551 => x"82",
          1552 => x"e1",
          1553 => x"39",
          1554 => x"54",
          1555 => x"80",
          1556 => x"3f",
          1557 => x"79",
          1558 => x"3f",
          1559 => x"33",
          1560 => x"2e",
          1561 => x"9f",
          1562 => x"38",
          1563 => x"fc",
          1564 => x"84",
          1565 => x"84",
          1566 => x"cc",
          1567 => x"91",
          1568 => x"02",
          1569 => x"33",
          1570 => x"81",
          1571 => x"b8",
          1572 => x"8c",
          1573 => x"3f",
          1574 => x"b4",
          1575 => x"11",
          1576 => x"05",
          1577 => x"3f",
          1578 => x"08",
          1579 => x"cb",
          1580 => x"fe",
          1581 => x"ff",
          1582 => x"a4",
          1583 => x"87",
          1584 => x"2e",
          1585 => x"59",
          1586 => x"22",
          1587 => x"05",
          1588 => x"41",
          1589 => x"f0",
          1590 => x"84",
          1591 => x"8e",
          1592 => x"cc",
          1593 => x"f4",
          1594 => x"70",
          1595 => x"81",
          1596 => x"a0",
          1597 => x"f8",
          1598 => x"a0",
          1599 => x"45",
          1600 => x"78",
          1601 => x"f3",
          1602 => x"26",
          1603 => x"82",
          1604 => x"39",
          1605 => x"f0",
          1606 => x"84",
          1607 => x"ce",
          1608 => x"cc",
          1609 => x"92",
          1610 => x"02",
          1611 => x"79",
          1612 => x"5b",
          1613 => x"ff",
          1614 => x"f4",
          1615 => x"e3",
          1616 => x"39",
          1617 => x"f4",
          1618 => x"84",
          1619 => x"9e",
          1620 => x"cc",
          1621 => x"f3",
          1622 => x"3d",
          1623 => x"53",
          1624 => x"51",
          1625 => x"82",
          1626 => x"80",
          1627 => x"60",
          1628 => x"59",
          1629 => x"41",
          1630 => x"f0",
          1631 => x"84",
          1632 => x"ea",
          1633 => x"cc",
          1634 => x"f2",
          1635 => x"70",
          1636 => x"81",
          1637 => x"9e",
          1638 => x"f8",
          1639 => x"9f",
          1640 => x"45",
          1641 => x"78",
          1642 => x"cf",
          1643 => x"27",
          1644 => x"3d",
          1645 => x"53",
          1646 => x"51",
          1647 => x"82",
          1648 => x"80",
          1649 => x"60",
          1650 => x"59",
          1651 => x"41",
          1652 => x"81",
          1653 => x"98",
          1654 => x"b2",
          1655 => x"ac",
          1656 => x"3f",
          1657 => x"a7",
          1658 => x"39",
          1659 => x"51",
          1660 => x"a2",
          1661 => x"3f",
          1662 => x"81",
          1663 => x"98",
          1664 => x"80",
          1665 => x"c0",
          1666 => x"84",
          1667 => x"87",
          1668 => x"0c",
          1669 => x"81",
          1670 => x"98",
          1671 => x"80",
          1672 => x"c0",
          1673 => x"8c",
          1674 => x"87",
          1675 => x"0c",
          1676 => x"b4",
          1677 => x"11",
          1678 => x"05",
          1679 => x"3f",
          1680 => x"08",
          1681 => x"b3",
          1682 => x"81",
          1683 => x"9d",
          1684 => x"59",
          1685 => x"3d",
          1686 => x"53",
          1687 => x"51",
          1688 => x"82",
          1689 => x"80",
          1690 => x"38",
          1691 => x"f5",
          1692 => x"93",
          1693 => x"78",
          1694 => x"cc",
          1695 => x"f0",
          1696 => x"87",
          1697 => x"81",
          1698 => x"9c",
          1699 => x"eb",
          1700 => x"d8",
          1701 => x"3f",
          1702 => x"f0",
          1703 => x"f5",
          1704 => x"ff",
          1705 => x"ff",
          1706 => x"e8",
          1707 => x"39",
          1708 => x"33",
          1709 => x"2e",
          1710 => x"7d",
          1711 => x"78",
          1712 => x"ce",
          1713 => x"ff",
          1714 => x"83",
          1715 => x"87",
          1716 => x"81",
          1717 => x"2e",
          1718 => x"82",
          1719 => x"7b",
          1720 => x"38",
          1721 => x"7b",
          1722 => x"38",
          1723 => x"81",
          1724 => x"7a",
          1725 => x"8c",
          1726 => x"81",
          1727 => x"b4",
          1728 => x"05",
          1729 => x"3f",
          1730 => x"f6",
          1731 => x"3d",
          1732 => x"51",
          1733 => x"a9",
          1734 => x"81",
          1735 => x"80",
          1736 => x"a0",
          1737 => x"ff",
          1738 => x"9b",
          1739 => x"39",
          1740 => x"53",
          1741 => x"52",
          1742 => x"b0",
          1743 => x"dd",
          1744 => x"f0",
          1745 => x"dc",
          1746 => x"64",
          1747 => x"82",
          1748 => x"82",
          1749 => x"b4",
          1750 => x"05",
          1751 => x"3f",
          1752 => x"08",
          1753 => x"08",
          1754 => x"70",
          1755 => x"25",
          1756 => x"5f",
          1757 => x"83",
          1758 => x"81",
          1759 => x"06",
          1760 => x"2e",
          1761 => x"1c",
          1762 => x"06",
          1763 => x"fe",
          1764 => x"81",
          1765 => x"32",
          1766 => x"8a",
          1767 => x"2e",
          1768 => x"ee",
          1769 => x"f6",
          1770 => x"db",
          1771 => x"39",
          1772 => x"80",
          1773 => x"dc",
          1774 => x"94",
          1775 => x"54",
          1776 => x"80",
          1777 => x"b4",
          1778 => x"87",
          1779 => x"2b",
          1780 => x"53",
          1781 => x"52",
          1782 => x"92",
          1783 => x"87",
          1784 => x"75",
          1785 => x"94",
          1786 => x"54",
          1787 => x"80",
          1788 => x"b3",
          1789 => x"87",
          1790 => x"2b",
          1791 => x"53",
          1792 => x"52",
          1793 => x"e6",
          1794 => x"87",
          1795 => x"75",
          1796 => x"83",
          1797 => x"94",
          1798 => x"80",
          1799 => x"c0",
          1800 => x"bd",
          1801 => x"9e",
          1802 => x"c0",
          1803 => x"9e",
          1804 => x"94",
          1805 => x"3f",
          1806 => x"51",
          1807 => x"81",
          1808 => x"93",
          1809 => x"ed",
          1810 => x"3f",
          1811 => x"e5",
          1812 => x"3f",
          1813 => x"3d",
          1814 => x"83",
          1815 => x"2b",
          1816 => x"3f",
          1817 => x"08",
          1818 => x"72",
          1819 => x"54",
          1820 => x"25",
          1821 => x"82",
          1822 => x"84",
          1823 => x"fc",
          1824 => x"70",
          1825 => x"80",
          1826 => x"72",
          1827 => x"8a",
          1828 => x"51",
          1829 => x"09",
          1830 => x"38",
          1831 => x"f1",
          1832 => x"51",
          1833 => x"09",
          1834 => x"38",
          1835 => x"81",
          1836 => x"73",
          1837 => x"81",
          1838 => x"84",
          1839 => x"52",
          1840 => x"52",
          1841 => x"2e",
          1842 => x"54",
          1843 => x"9d",
          1844 => x"38",
          1845 => x"12",
          1846 => x"33",
          1847 => x"a0",
          1848 => x"81",
          1849 => x"2e",
          1850 => x"ea",
          1851 => x"33",
          1852 => x"a0",
          1853 => x"06",
          1854 => x"54",
          1855 => x"70",
          1856 => x"25",
          1857 => x"51",
          1858 => x"2e",
          1859 => x"72",
          1860 => x"54",
          1861 => x"0c",
          1862 => x"82",
          1863 => x"86",
          1864 => x"fc",
          1865 => x"53",
          1866 => x"2e",
          1867 => x"3d",
          1868 => x"72",
          1869 => x"3f",
          1870 => x"08",
          1871 => x"53",
          1872 => x"53",
          1873 => x"cc",
          1874 => x"0d",
          1875 => x"0d",
          1876 => x"33",
          1877 => x"53",
          1878 => x"8b",
          1879 => x"38",
          1880 => x"ff",
          1881 => x"52",
          1882 => x"81",
          1883 => x"13",
          1884 => x"52",
          1885 => x"80",
          1886 => x"13",
          1887 => x"52",
          1888 => x"80",
          1889 => x"13",
          1890 => x"52",
          1891 => x"80",
          1892 => x"13",
          1893 => x"52",
          1894 => x"26",
          1895 => x"8a",
          1896 => x"87",
          1897 => x"e7",
          1898 => x"38",
          1899 => x"c0",
          1900 => x"72",
          1901 => x"98",
          1902 => x"13",
          1903 => x"98",
          1904 => x"13",
          1905 => x"98",
          1906 => x"13",
          1907 => x"98",
          1908 => x"13",
          1909 => x"98",
          1910 => x"13",
          1911 => x"98",
          1912 => x"87",
          1913 => x"0c",
          1914 => x"98",
          1915 => x"0b",
          1916 => x"9c",
          1917 => x"71",
          1918 => x"0c",
          1919 => x"04",
          1920 => x"7f",
          1921 => x"98",
          1922 => x"7d",
          1923 => x"98",
          1924 => x"7d",
          1925 => x"c0",
          1926 => x"5a",
          1927 => x"34",
          1928 => x"b4",
          1929 => x"83",
          1930 => x"c0",
          1931 => x"5a",
          1932 => x"34",
          1933 => x"ac",
          1934 => x"85",
          1935 => x"c0",
          1936 => x"5a",
          1937 => x"34",
          1938 => x"a4",
          1939 => x"88",
          1940 => x"c0",
          1941 => x"5a",
          1942 => x"23",
          1943 => x"79",
          1944 => x"06",
          1945 => x"ff",
          1946 => x"86",
          1947 => x"85",
          1948 => x"84",
          1949 => x"83",
          1950 => x"82",
          1951 => x"7d",
          1952 => x"06",
          1953 => x"e8",
          1954 => x"3f",
          1955 => x"04",
          1956 => x"02",
          1957 => x"70",
          1958 => x"2a",
          1959 => x"70",
          1960 => x"34",
          1961 => x"04",
          1962 => x"77",
          1963 => x"33",
          1964 => x"06",
          1965 => x"87",
          1966 => x"51",
          1967 => x"86",
          1968 => x"94",
          1969 => x"08",
          1970 => x"70",
          1971 => x"54",
          1972 => x"2e",
          1973 => x"91",
          1974 => x"06",
          1975 => x"d7",
          1976 => x"32",
          1977 => x"51",
          1978 => x"2e",
          1979 => x"93",
          1980 => x"06",
          1981 => x"ff",
          1982 => x"81",
          1983 => x"87",
          1984 => x"52",
          1985 => x"86",
          1986 => x"94",
          1987 => x"72",
          1988 => x"87",
          1989 => x"3d",
          1990 => x"3d",
          1991 => x"05",
          1992 => x"ec",
          1993 => x"ff",
          1994 => x"56",
          1995 => x"84",
          1996 => x"2e",
          1997 => x"c0",
          1998 => x"70",
          1999 => x"2a",
          2000 => x"53",
          2001 => x"80",
          2002 => x"71",
          2003 => x"81",
          2004 => x"70",
          2005 => x"81",
          2006 => x"06",
          2007 => x"80",
          2008 => x"71",
          2009 => x"81",
          2010 => x"70",
          2011 => x"73",
          2012 => x"51",
          2013 => x"80",
          2014 => x"2e",
          2015 => x"c0",
          2016 => x"75",
          2017 => x"3d",
          2018 => x"3d",
          2019 => x"80",
          2020 => x"81",
          2021 => x"53",
          2022 => x"2e",
          2023 => x"71",
          2024 => x"81",
          2025 => x"ec",
          2026 => x"ff",
          2027 => x"55",
          2028 => x"94",
          2029 => x"80",
          2030 => x"87",
          2031 => x"51",
          2032 => x"96",
          2033 => x"06",
          2034 => x"70",
          2035 => x"38",
          2036 => x"70",
          2037 => x"51",
          2038 => x"72",
          2039 => x"81",
          2040 => x"70",
          2041 => x"38",
          2042 => x"70",
          2043 => x"51",
          2044 => x"38",
          2045 => x"06",
          2046 => x"94",
          2047 => x"80",
          2048 => x"87",
          2049 => x"52",
          2050 => x"81",
          2051 => x"70",
          2052 => x"53",
          2053 => x"ff",
          2054 => x"82",
          2055 => x"89",
          2056 => x"fe",
          2057 => x"85",
          2058 => x"81",
          2059 => x"52",
          2060 => x"84",
          2061 => x"2e",
          2062 => x"c0",
          2063 => x"70",
          2064 => x"2a",
          2065 => x"51",
          2066 => x"80",
          2067 => x"71",
          2068 => x"51",
          2069 => x"80",
          2070 => x"2e",
          2071 => x"c0",
          2072 => x"71",
          2073 => x"ff",
          2074 => x"cc",
          2075 => x"3d",
          2076 => x"3d",
          2077 => x"ec",
          2078 => x"ff",
          2079 => x"87",
          2080 => x"52",
          2081 => x"86",
          2082 => x"94",
          2083 => x"08",
          2084 => x"70",
          2085 => x"51",
          2086 => x"70",
          2087 => x"38",
          2088 => x"06",
          2089 => x"94",
          2090 => x"80",
          2091 => x"87",
          2092 => x"52",
          2093 => x"98",
          2094 => x"2c",
          2095 => x"71",
          2096 => x"0c",
          2097 => x"04",
          2098 => x"87",
          2099 => x"08",
          2100 => x"8a",
          2101 => x"70",
          2102 => x"b4",
          2103 => x"9e",
          2104 => x"85",
          2105 => x"c0",
          2106 => x"82",
          2107 => x"87",
          2108 => x"08",
          2109 => x"0c",
          2110 => x"98",
          2111 => x"fc",
          2112 => x"9e",
          2113 => x"86",
          2114 => x"c0",
          2115 => x"82",
          2116 => x"87",
          2117 => x"08",
          2118 => x"0c",
          2119 => x"b0",
          2120 => x"8c",
          2121 => x"9e",
          2122 => x"86",
          2123 => x"c0",
          2124 => x"82",
          2125 => x"87",
          2126 => x"08",
          2127 => x"0c",
          2128 => x"c0",
          2129 => x"9c",
          2130 => x"9e",
          2131 => x"86",
          2132 => x"c0",
          2133 => x"51",
          2134 => x"a4",
          2135 => x"9e",
          2136 => x"86",
          2137 => x"c0",
          2138 => x"82",
          2139 => x"87",
          2140 => x"08",
          2141 => x"0c",
          2142 => x"86",
          2143 => x"0b",
          2144 => x"90",
          2145 => x"80",
          2146 => x"52",
          2147 => x"2e",
          2148 => x"52",
          2149 => x"b5",
          2150 => x"87",
          2151 => x"08",
          2152 => x"0a",
          2153 => x"52",
          2154 => x"83",
          2155 => x"71",
          2156 => x"34",
          2157 => x"c0",
          2158 => x"70",
          2159 => x"06",
          2160 => x"70",
          2161 => x"38",
          2162 => x"82",
          2163 => x"80",
          2164 => x"9e",
          2165 => x"88",
          2166 => x"51",
          2167 => x"80",
          2168 => x"81",
          2169 => x"86",
          2170 => x"0b",
          2171 => x"90",
          2172 => x"80",
          2173 => x"52",
          2174 => x"2e",
          2175 => x"52",
          2176 => x"b9",
          2177 => x"87",
          2178 => x"08",
          2179 => x"80",
          2180 => x"52",
          2181 => x"83",
          2182 => x"71",
          2183 => x"34",
          2184 => x"c0",
          2185 => x"70",
          2186 => x"06",
          2187 => x"70",
          2188 => x"38",
          2189 => x"82",
          2190 => x"80",
          2191 => x"9e",
          2192 => x"82",
          2193 => x"51",
          2194 => x"80",
          2195 => x"81",
          2196 => x"86",
          2197 => x"0b",
          2198 => x"90",
          2199 => x"80",
          2200 => x"52",
          2201 => x"2e",
          2202 => x"52",
          2203 => x"bd",
          2204 => x"87",
          2205 => x"08",
          2206 => x"80",
          2207 => x"52",
          2208 => x"83",
          2209 => x"71",
          2210 => x"34",
          2211 => x"c0",
          2212 => x"70",
          2213 => x"51",
          2214 => x"80",
          2215 => x"81",
          2216 => x"86",
          2217 => x"c0",
          2218 => x"70",
          2219 => x"70",
          2220 => x"51",
          2221 => x"86",
          2222 => x"0b",
          2223 => x"90",
          2224 => x"80",
          2225 => x"52",
          2226 => x"83",
          2227 => x"71",
          2228 => x"34",
          2229 => x"90",
          2230 => x"f0",
          2231 => x"2a",
          2232 => x"70",
          2233 => x"34",
          2234 => x"c0",
          2235 => x"70",
          2236 => x"52",
          2237 => x"2e",
          2238 => x"52",
          2239 => x"c3",
          2240 => x"9e",
          2241 => x"87",
          2242 => x"70",
          2243 => x"34",
          2244 => x"04",
          2245 => x"81",
          2246 => x"86",
          2247 => x"86",
          2248 => x"73",
          2249 => x"38",
          2250 => x"51",
          2251 => x"81",
          2252 => x"85",
          2253 => x"86",
          2254 => x"73",
          2255 => x"38",
          2256 => x"08",
          2257 => x"08",
          2258 => x"81",
          2259 => x"8b",
          2260 => x"86",
          2261 => x"73",
          2262 => x"38",
          2263 => x"08",
          2264 => x"08",
          2265 => x"81",
          2266 => x"8b",
          2267 => x"86",
          2268 => x"73",
          2269 => x"38",
          2270 => x"08",
          2271 => x"08",
          2272 => x"81",
          2273 => x"8a",
          2274 => x"86",
          2275 => x"73",
          2276 => x"38",
          2277 => x"08",
          2278 => x"08",
          2279 => x"81",
          2280 => x"8a",
          2281 => x"86",
          2282 => x"73",
          2283 => x"38",
          2284 => x"08",
          2285 => x"08",
          2286 => x"81",
          2287 => x"8a",
          2288 => x"86",
          2289 => x"73",
          2290 => x"38",
          2291 => x"33",
          2292 => x"cc",
          2293 => x"3f",
          2294 => x"33",
          2295 => x"2e",
          2296 => x"86",
          2297 => x"81",
          2298 => x"8a",
          2299 => x"86",
          2300 => x"73",
          2301 => x"38",
          2302 => x"33",
          2303 => x"8c",
          2304 => x"3f",
          2305 => x"33",
          2306 => x"2e",
          2307 => x"f9",
          2308 => x"8f",
          2309 => x"b7",
          2310 => x"80",
          2311 => x"81",
          2312 => x"83",
          2313 => x"86",
          2314 => x"73",
          2315 => x"38",
          2316 => x"51",
          2317 => x"82",
          2318 => x"54",
          2319 => x"88",
          2320 => x"d8",
          2321 => x"3f",
          2322 => x"33",
          2323 => x"2e",
          2324 => x"f9",
          2325 => x"cb",
          2326 => x"f0",
          2327 => x"3f",
          2328 => x"08",
          2329 => x"fc",
          2330 => x"3f",
          2331 => x"08",
          2332 => x"a4",
          2333 => x"3f",
          2334 => x"08",
          2335 => x"cc",
          2336 => x"3f",
          2337 => x"51",
          2338 => x"82",
          2339 => x"52",
          2340 => x"51",
          2341 => x"82",
          2342 => x"56",
          2343 => x"52",
          2344 => x"ca",
          2345 => x"cc",
          2346 => x"c0",
          2347 => x"31",
          2348 => x"87",
          2349 => x"81",
          2350 => x"88",
          2351 => x"86",
          2352 => x"73",
          2353 => x"38",
          2354 => x"08",
          2355 => x"c0",
          2356 => x"a2",
          2357 => x"87",
          2358 => x"84",
          2359 => x"71",
          2360 => x"82",
          2361 => x"52",
          2362 => x"51",
          2363 => x"82",
          2364 => x"54",
          2365 => x"a8",
          2366 => x"b0",
          2367 => x"84",
          2368 => x"51",
          2369 => x"82",
          2370 => x"bd",
          2371 => x"76",
          2372 => x"54",
          2373 => x"08",
          2374 => x"fc",
          2375 => x"3f",
          2376 => x"51",
          2377 => x"87",
          2378 => x"fe",
          2379 => x"92",
          2380 => x"05",
          2381 => x"26",
          2382 => x"84",
          2383 => x"94",
          2384 => x"08",
          2385 => x"a8",
          2386 => x"81",
          2387 => x"97",
          2388 => x"b8",
          2389 => x"81",
          2390 => x"8b",
          2391 => x"c4",
          2392 => x"81",
          2393 => x"81",
          2394 => x"3d",
          2395 => x"88",
          2396 => x"ff",
          2397 => x"c0",
          2398 => x"08",
          2399 => x"72",
          2400 => x"07",
          2401 => x"c8",
          2402 => x"83",
          2403 => x"ff",
          2404 => x"c0",
          2405 => x"08",
          2406 => x"0c",
          2407 => x"0c",
          2408 => x"82",
          2409 => x"06",
          2410 => x"c8",
          2411 => x"51",
          2412 => x"04",
          2413 => x"c0",
          2414 => x"04",
          2415 => x"08",
          2416 => x"84",
          2417 => x"3d",
          2418 => x"05",
          2419 => x"8a",
          2420 => x"06",
          2421 => x"51",
          2422 => x"9e",
          2423 => x"71",
          2424 => x"38",
          2425 => x"82",
          2426 => x"81",
          2427 => x"dc",
          2428 => x"82",
          2429 => x"52",
          2430 => x"85",
          2431 => x"71",
          2432 => x"0d",
          2433 => x"0d",
          2434 => x"33",
          2435 => x"08",
          2436 => x"d4",
          2437 => x"ff",
          2438 => x"82",
          2439 => x"84",
          2440 => x"fd",
          2441 => x"54",
          2442 => x"81",
          2443 => x"53",
          2444 => x"8e",
          2445 => x"ff",
          2446 => x"14",
          2447 => x"3f",
          2448 => x"3d",
          2449 => x"3d",
          2450 => x"9e",
          2451 => x"82",
          2452 => x"56",
          2453 => x"70",
          2454 => x"53",
          2455 => x"2e",
          2456 => x"81",
          2457 => x"81",
          2458 => x"da",
          2459 => x"74",
          2460 => x"0c",
          2461 => x"04",
          2462 => x"66",
          2463 => x"78",
          2464 => x"5a",
          2465 => x"80",
          2466 => x"38",
          2467 => x"09",
          2468 => x"de",
          2469 => x"7a",
          2470 => x"5c",
          2471 => x"5b",
          2472 => x"09",
          2473 => x"38",
          2474 => x"39",
          2475 => x"09",
          2476 => x"38",
          2477 => x"70",
          2478 => x"33",
          2479 => x"2e",
          2480 => x"92",
          2481 => x"19",
          2482 => x"70",
          2483 => x"33",
          2484 => x"53",
          2485 => x"16",
          2486 => x"26",
          2487 => x"88",
          2488 => x"05",
          2489 => x"05",
          2490 => x"05",
          2491 => x"5b",
          2492 => x"80",
          2493 => x"30",
          2494 => x"80",
          2495 => x"cc",
          2496 => x"70",
          2497 => x"25",
          2498 => x"54",
          2499 => x"53",
          2500 => x"8c",
          2501 => x"07",
          2502 => x"05",
          2503 => x"5a",
          2504 => x"83",
          2505 => x"54",
          2506 => x"27",
          2507 => x"16",
          2508 => x"06",
          2509 => x"80",
          2510 => x"aa",
          2511 => x"cf",
          2512 => x"73",
          2513 => x"81",
          2514 => x"80",
          2515 => x"38",
          2516 => x"2e",
          2517 => x"81",
          2518 => x"80",
          2519 => x"8a",
          2520 => x"39",
          2521 => x"2e",
          2522 => x"73",
          2523 => x"8a",
          2524 => x"d3",
          2525 => x"80",
          2526 => x"80",
          2527 => x"ee",
          2528 => x"39",
          2529 => x"71",
          2530 => x"53",
          2531 => x"54",
          2532 => x"2e",
          2533 => x"15",
          2534 => x"33",
          2535 => x"72",
          2536 => x"81",
          2537 => x"39",
          2538 => x"56",
          2539 => x"27",
          2540 => x"51",
          2541 => x"75",
          2542 => x"72",
          2543 => x"38",
          2544 => x"df",
          2545 => x"16",
          2546 => x"7b",
          2547 => x"38",
          2548 => x"f2",
          2549 => x"77",
          2550 => x"12",
          2551 => x"53",
          2552 => x"5c",
          2553 => x"5c",
          2554 => x"5c",
          2555 => x"5c",
          2556 => x"51",
          2557 => x"fd",
          2558 => x"82",
          2559 => x"06",
          2560 => x"80",
          2561 => x"77",
          2562 => x"53",
          2563 => x"18",
          2564 => x"72",
          2565 => x"c4",
          2566 => x"70",
          2567 => x"25",
          2568 => x"55",
          2569 => x"8d",
          2570 => x"2e",
          2571 => x"30",
          2572 => x"5b",
          2573 => x"8f",
          2574 => x"7b",
          2575 => x"9d",
          2576 => x"87",
          2577 => x"ff",
          2578 => x"75",
          2579 => x"9e",
          2580 => x"cc",
          2581 => x"74",
          2582 => x"a7",
          2583 => x"80",
          2584 => x"38",
          2585 => x"72",
          2586 => x"54",
          2587 => x"72",
          2588 => x"05",
          2589 => x"17",
          2590 => x"77",
          2591 => x"51",
          2592 => x"9f",
          2593 => x"72",
          2594 => x"79",
          2595 => x"81",
          2596 => x"72",
          2597 => x"38",
          2598 => x"05",
          2599 => x"ad",
          2600 => x"17",
          2601 => x"81",
          2602 => x"b0",
          2603 => x"38",
          2604 => x"81",
          2605 => x"06",
          2606 => x"9f",
          2607 => x"55",
          2608 => x"97",
          2609 => x"f9",
          2610 => x"81",
          2611 => x"8b",
          2612 => x"16",
          2613 => x"73",
          2614 => x"96",
          2615 => x"e0",
          2616 => x"17",
          2617 => x"33",
          2618 => x"f9",
          2619 => x"f2",
          2620 => x"16",
          2621 => x"7b",
          2622 => x"38",
          2623 => x"c6",
          2624 => x"96",
          2625 => x"fd",
          2626 => x"3d",
          2627 => x"05",
          2628 => x"52",
          2629 => x"e0",
          2630 => x"0d",
          2631 => x"0d",
          2632 => x"dc",
          2633 => x"88",
          2634 => x"51",
          2635 => x"82",
          2636 => x"53",
          2637 => x"80",
          2638 => x"dc",
          2639 => x"0d",
          2640 => x"0d",
          2641 => x"08",
          2642 => x"d4",
          2643 => x"88",
          2644 => x"52",
          2645 => x"3f",
          2646 => x"d4",
          2647 => x"0d",
          2648 => x"0d",
          2649 => x"9e",
          2650 => x"56",
          2651 => x"80",
          2652 => x"2e",
          2653 => x"82",
          2654 => x"52",
          2655 => x"87",
          2656 => x"ff",
          2657 => x"80",
          2658 => x"38",
          2659 => x"b9",
          2660 => x"32",
          2661 => x"80",
          2662 => x"52",
          2663 => x"8b",
          2664 => x"2e",
          2665 => x"14",
          2666 => x"9f",
          2667 => x"38",
          2668 => x"73",
          2669 => x"38",
          2670 => x"72",
          2671 => x"14",
          2672 => x"f8",
          2673 => x"af",
          2674 => x"52",
          2675 => x"8a",
          2676 => x"3f",
          2677 => x"82",
          2678 => x"87",
          2679 => x"fe",
          2680 => x"9e",
          2681 => x"82",
          2682 => x"77",
          2683 => x"53",
          2684 => x"72",
          2685 => x"0c",
          2686 => x"04",
          2687 => x"7a",
          2688 => x"80",
          2689 => x"58",
          2690 => x"33",
          2691 => x"a0",
          2692 => x"06",
          2693 => x"13",
          2694 => x"39",
          2695 => x"09",
          2696 => x"38",
          2697 => x"11",
          2698 => x"08",
          2699 => x"54",
          2700 => x"2e",
          2701 => x"80",
          2702 => x"08",
          2703 => x"0c",
          2704 => x"33",
          2705 => x"80",
          2706 => x"38",
          2707 => x"80",
          2708 => x"38",
          2709 => x"57",
          2710 => x"0c",
          2711 => x"33",
          2712 => x"39",
          2713 => x"74",
          2714 => x"38",
          2715 => x"80",
          2716 => x"89",
          2717 => x"38",
          2718 => x"d0",
          2719 => x"55",
          2720 => x"80",
          2721 => x"39",
          2722 => x"d9",
          2723 => x"80",
          2724 => x"27",
          2725 => x"80",
          2726 => x"89",
          2727 => x"70",
          2728 => x"55",
          2729 => x"70",
          2730 => x"55",
          2731 => x"27",
          2732 => x"14",
          2733 => x"06",
          2734 => x"74",
          2735 => x"73",
          2736 => x"38",
          2737 => x"14",
          2738 => x"05",
          2739 => x"08",
          2740 => x"54",
          2741 => x"39",
          2742 => x"84",
          2743 => x"55",
          2744 => x"81",
          2745 => x"87",
          2746 => x"3d",
          2747 => x"3d",
          2748 => x"5a",
          2749 => x"7a",
          2750 => x"08",
          2751 => x"53",
          2752 => x"09",
          2753 => x"38",
          2754 => x"0c",
          2755 => x"ad",
          2756 => x"06",
          2757 => x"76",
          2758 => x"0c",
          2759 => x"33",
          2760 => x"73",
          2761 => x"81",
          2762 => x"38",
          2763 => x"05",
          2764 => x"08",
          2765 => x"53",
          2766 => x"2e",
          2767 => x"57",
          2768 => x"2e",
          2769 => x"39",
          2770 => x"13",
          2771 => x"08",
          2772 => x"53",
          2773 => x"55",
          2774 => x"80",
          2775 => x"14",
          2776 => x"88",
          2777 => x"27",
          2778 => x"eb",
          2779 => x"53",
          2780 => x"89",
          2781 => x"38",
          2782 => x"55",
          2783 => x"8a",
          2784 => x"a0",
          2785 => x"c2",
          2786 => x"74",
          2787 => x"e0",
          2788 => x"ff",
          2789 => x"d0",
          2790 => x"ff",
          2791 => x"90",
          2792 => x"38",
          2793 => x"81",
          2794 => x"53",
          2795 => x"ca",
          2796 => x"27",
          2797 => x"77",
          2798 => x"08",
          2799 => x"0c",
          2800 => x"33",
          2801 => x"ff",
          2802 => x"80",
          2803 => x"74",
          2804 => x"79",
          2805 => x"74",
          2806 => x"0c",
          2807 => x"04",
          2808 => x"76",
          2809 => x"98",
          2810 => x"2b",
          2811 => x"72",
          2812 => x"82",
          2813 => x"51",
          2814 => x"80",
          2815 => x"d8",
          2816 => x"53",
          2817 => x"9c",
          2818 => x"d4",
          2819 => x"02",
          2820 => x"05",
          2821 => x"52",
          2822 => x"72",
          2823 => x"06",
          2824 => x"53",
          2825 => x"cc",
          2826 => x"0d",
          2827 => x"0d",
          2828 => x"05",
          2829 => x"71",
          2830 => x"53",
          2831 => x"9f",
          2832 => x"f3",
          2833 => x"51",
          2834 => x"88",
          2835 => x"3f",
          2836 => x"05",
          2837 => x"34",
          2838 => x"06",
          2839 => x"76",
          2840 => x"3f",
          2841 => x"86",
          2842 => x"f6",
          2843 => x"02",
          2844 => x"05",
          2845 => x"05",
          2846 => x"82",
          2847 => x"70",
          2848 => x"86",
          2849 => x"08",
          2850 => x"5a",
          2851 => x"80",
          2852 => x"74",
          2853 => x"3f",
          2854 => x"33",
          2855 => x"82",
          2856 => x"81",
          2857 => x"58",
          2858 => x"84",
          2859 => x"cc",
          2860 => x"82",
          2861 => x"70",
          2862 => x"86",
          2863 => x"08",
          2864 => x"74",
          2865 => x"38",
          2866 => x"52",
          2867 => x"bb",
          2868 => x"87",
          2869 => x"05",
          2870 => x"87",
          2871 => x"81",
          2872 => x"93",
          2873 => x"38",
          2874 => x"87",
          2875 => x"80",
          2876 => x"82",
          2877 => x"56",
          2878 => x"ac",
          2879 => x"9c",
          2880 => x"a4",
          2881 => x"fc",
          2882 => x"53",
          2883 => x"51",
          2884 => x"3f",
          2885 => x"08",
          2886 => x"81",
          2887 => x"82",
          2888 => x"51",
          2889 => x"3f",
          2890 => x"04",
          2891 => x"82",
          2892 => x"93",
          2893 => x"52",
          2894 => x"89",
          2895 => x"9c",
          2896 => x"73",
          2897 => x"84",
          2898 => x"73",
          2899 => x"38",
          2900 => x"87",
          2901 => x"87",
          2902 => x"71",
          2903 => x"38",
          2904 => x"dd",
          2905 => x"87",
          2906 => x"9c",
          2907 => x"0b",
          2908 => x"0c",
          2909 => x"04",
          2910 => x"81",
          2911 => x"82",
          2912 => x"51",
          2913 => x"3f",
          2914 => x"08",
          2915 => x"82",
          2916 => x"53",
          2917 => x"88",
          2918 => x"56",
          2919 => x"3f",
          2920 => x"08",
          2921 => x"38",
          2922 => x"b8",
          2923 => x"87",
          2924 => x"80",
          2925 => x"cc",
          2926 => x"38",
          2927 => x"08",
          2928 => x"17",
          2929 => x"74",
          2930 => x"76",
          2931 => x"81",
          2932 => x"57",
          2933 => x"74",
          2934 => x"81",
          2935 => x"38",
          2936 => x"04",
          2937 => x"aa",
          2938 => x"3d",
          2939 => x"81",
          2940 => x"80",
          2941 => x"a0",
          2942 => x"e1",
          2943 => x"87",
          2944 => x"94",
          2945 => x"82",
          2946 => x"54",
          2947 => x"52",
          2948 => x"52",
          2949 => x"e8",
          2950 => x"cc",
          2951 => x"a5",
          2952 => x"ff",
          2953 => x"82",
          2954 => x"81",
          2955 => x"80",
          2956 => x"cc",
          2957 => x"38",
          2958 => x"08",
          2959 => x"17",
          2960 => x"74",
          2961 => x"70",
          2962 => x"07",
          2963 => x"55",
          2964 => x"2e",
          2965 => x"ff",
          2966 => x"87",
          2967 => x"11",
          2968 => x"80",
          2969 => x"82",
          2970 => x"80",
          2971 => x"81",
          2972 => x"ef",
          2973 => x"77",
          2974 => x"06",
          2975 => x"52",
          2976 => x"b7",
          2977 => x"51",
          2978 => x"3f",
          2979 => x"54",
          2980 => x"08",
          2981 => x"58",
          2982 => x"cc",
          2983 => x"0d",
          2984 => x"0d",
          2985 => x"5c",
          2986 => x"57",
          2987 => x"73",
          2988 => x"81",
          2989 => x"78",
          2990 => x"56",
          2991 => x"98",
          2992 => x"70",
          2993 => x"33",
          2994 => x"73",
          2995 => x"81",
          2996 => x"75",
          2997 => x"38",
          2998 => x"88",
          2999 => x"a8",
          3000 => x"52",
          3001 => x"d2",
          3002 => x"cc",
          3003 => x"52",
          3004 => x"ff",
          3005 => x"82",
          3006 => x"80",
          3007 => x"15",
          3008 => x"81",
          3009 => x"74",
          3010 => x"38",
          3011 => x"e8",
          3012 => x"81",
          3013 => x"3d",
          3014 => x"f8",
          3015 => x"dc",
          3016 => x"cc",
          3017 => x"9a",
          3018 => x"53",
          3019 => x"51",
          3020 => x"82",
          3021 => x"81",
          3022 => x"74",
          3023 => x"54",
          3024 => x"14",
          3025 => x"06",
          3026 => x"74",
          3027 => x"38",
          3028 => x"82",
          3029 => x"8c",
          3030 => x"d3",
          3031 => x"3d",
          3032 => x"08",
          3033 => x"59",
          3034 => x"0b",
          3035 => x"82",
          3036 => x"82",
          3037 => x"55",
          3038 => x"ca",
          3039 => x"87",
          3040 => x"55",
          3041 => x"81",
          3042 => x"2e",
          3043 => x"81",
          3044 => x"55",
          3045 => x"2e",
          3046 => x"a8",
          3047 => x"3f",
          3048 => x"08",
          3049 => x"0c",
          3050 => x"08",
          3051 => x"91",
          3052 => x"76",
          3053 => x"cc",
          3054 => x"cb",
          3055 => x"87",
          3056 => x"2e",
          3057 => x"80",
          3058 => x"bb",
          3059 => x"39",
          3060 => x"08",
          3061 => x"a0",
          3062 => x"f8",
          3063 => x"70",
          3064 => x"86",
          3065 => x"87",
          3066 => x"82",
          3067 => x"74",
          3068 => x"06",
          3069 => x"82",
          3070 => x"51",
          3071 => x"3f",
          3072 => x"08",
          3073 => x"82",
          3074 => x"25",
          3075 => x"87",
          3076 => x"05",
          3077 => x"55",
          3078 => x"80",
          3079 => x"ff",
          3080 => x"51",
          3081 => x"81",
          3082 => x"ff",
          3083 => x"93",
          3084 => x"38",
          3085 => x"ff",
          3086 => x"06",
          3087 => x"86",
          3088 => x"87",
          3089 => x"8c",
          3090 => x"a0",
          3091 => x"84",
          3092 => x"3f",
          3093 => x"e0",
          3094 => x"87",
          3095 => x"2b",
          3096 => x"51",
          3097 => x"2e",
          3098 => x"81",
          3099 => x"9e",
          3100 => x"98",
          3101 => x"2c",
          3102 => x"33",
          3103 => x"70",
          3104 => x"98",
          3105 => x"84",
          3106 => x"d4",
          3107 => x"15",
          3108 => x"51",
          3109 => x"59",
          3110 => x"58",
          3111 => x"78",
          3112 => x"38",
          3113 => x"b4",
          3114 => x"80",
          3115 => x"ff",
          3116 => x"98",
          3117 => x"80",
          3118 => x"ce",
          3119 => x"74",
          3120 => x"f6",
          3121 => x"87",
          3122 => x"ff",
          3123 => x"80",
          3124 => x"74",
          3125 => x"34",
          3126 => x"39",
          3127 => x"0a",
          3128 => x"0a",
          3129 => x"2c",
          3130 => x"06",
          3131 => x"73",
          3132 => x"38",
          3133 => x"52",
          3134 => x"e4",
          3135 => x"cc",
          3136 => x"06",
          3137 => x"38",
          3138 => x"56",
          3139 => x"80",
          3140 => x"1c",
          3141 => x"9e",
          3142 => x"98",
          3143 => x"2c",
          3144 => x"33",
          3145 => x"70",
          3146 => x"10",
          3147 => x"2b",
          3148 => x"11",
          3149 => x"51",
          3150 => x"51",
          3151 => x"2e",
          3152 => x"fe",
          3153 => x"fc",
          3154 => x"7d",
          3155 => x"82",
          3156 => x"80",
          3157 => x"e0",
          3158 => x"75",
          3159 => x"34",
          3160 => x"e0",
          3161 => x"3d",
          3162 => x"0c",
          3163 => x"95",
          3164 => x"38",
          3165 => x"81",
          3166 => x"54",
          3167 => x"82",
          3168 => x"54",
          3169 => x"fd",
          3170 => x"9e",
          3171 => x"73",
          3172 => x"38",
          3173 => x"70",
          3174 => x"55",
          3175 => x"9e",
          3176 => x"54",
          3177 => x"15",
          3178 => x"80",
          3179 => x"ff",
          3180 => x"98",
          3181 => x"ec",
          3182 => x"55",
          3183 => x"9e",
          3184 => x"11",
          3185 => x"82",
          3186 => x"73",
          3187 => x"3d",
          3188 => x"82",
          3189 => x"54",
          3190 => x"89",
          3191 => x"54",
          3192 => x"e8",
          3193 => x"ec",
          3194 => x"80",
          3195 => x"ff",
          3196 => x"98",
          3197 => x"e8",
          3198 => x"56",
          3199 => x"25",
          3200 => x"1a",
          3201 => x"54",
          3202 => x"74",
          3203 => x"29",
          3204 => x"05",
          3205 => x"82",
          3206 => x"56",
          3207 => x"75",
          3208 => x"82",
          3209 => x"70",
          3210 => x"98",
          3211 => x"e8",
          3212 => x"56",
          3213 => x"25",
          3214 => x"88",
          3215 => x"3f",
          3216 => x"0a",
          3217 => x"0a",
          3218 => x"2c",
          3219 => x"33",
          3220 => x"73",
          3221 => x"38",
          3222 => x"83",
          3223 => x"0b",
          3224 => x"82",
          3225 => x"80",
          3226 => x"b8",
          3227 => x"3f",
          3228 => x"82",
          3229 => x"70",
          3230 => x"55",
          3231 => x"2e",
          3232 => x"82",
          3233 => x"ff",
          3234 => x"82",
          3235 => x"ff",
          3236 => x"82",
          3237 => x"88",
          3238 => x"3f",
          3239 => x"33",
          3240 => x"70",
          3241 => x"9e",
          3242 => x"51",
          3243 => x"74",
          3244 => x"74",
          3245 => x"14",
          3246 => x"73",
          3247 => x"86",
          3248 => x"80",
          3249 => x"80",
          3250 => x"98",
          3251 => x"e8",
          3252 => x"55",
          3253 => x"db",
          3254 => x"e5",
          3255 => x"9e",
          3256 => x"98",
          3257 => x"2c",
          3258 => x"33",
          3259 => x"57",
          3260 => x"fa",
          3261 => x"51",
          3262 => x"74",
          3263 => x"29",
          3264 => x"05",
          3265 => x"82",
          3266 => x"58",
          3267 => x"75",
          3268 => x"fa",
          3269 => x"9e",
          3270 => x"05",
          3271 => x"34",
          3272 => x"a2",
          3273 => x"e8",
          3274 => x"f6",
          3275 => x"87",
          3276 => x"ff",
          3277 => x"96",
          3278 => x"e8",
          3279 => x"80",
          3280 => x"81",
          3281 => x"79",
          3282 => x"3f",
          3283 => x"7a",
          3284 => x"82",
          3285 => x"80",
          3286 => x"e8",
          3287 => x"87",
          3288 => x"3d",
          3289 => x"9e",
          3290 => x"73",
          3291 => x"e4",
          3292 => x"e4",
          3293 => x"9e",
          3294 => x"05",
          3295 => x"9e",
          3296 => x"81",
          3297 => x"e3",
          3298 => x"ec",
          3299 => x"e8",
          3300 => x"73",
          3301 => x"bc",
          3302 => x"54",
          3303 => x"e8",
          3304 => x"2b",
          3305 => x"75",
          3306 => x"56",
          3307 => x"74",
          3308 => x"74",
          3309 => x"14",
          3310 => x"73",
          3311 => x"86",
          3312 => x"80",
          3313 => x"80",
          3314 => x"98",
          3315 => x"e8",
          3316 => x"55",
          3317 => x"db",
          3318 => x"e3",
          3319 => x"9e",
          3320 => x"98",
          3321 => x"2c",
          3322 => x"33",
          3323 => x"57",
          3324 => x"f8",
          3325 => x"51",
          3326 => x"74",
          3327 => x"29",
          3328 => x"05",
          3329 => x"82",
          3330 => x"58",
          3331 => x"75",
          3332 => x"f8",
          3333 => x"9e",
          3334 => x"81",
          3335 => x"9e",
          3336 => x"56",
          3337 => x"27",
          3338 => x"81",
          3339 => x"82",
          3340 => x"74",
          3341 => x"52",
          3342 => x"3f",
          3343 => x"33",
          3344 => x"06",
          3345 => x"33",
          3346 => x"75",
          3347 => x"38",
          3348 => x"82",
          3349 => x"80",
          3350 => x"b8",
          3351 => x"3f",
          3352 => x"9e",
          3353 => x"0b",
          3354 => x"34",
          3355 => x"7a",
          3356 => x"87",
          3357 => x"74",
          3358 => x"38",
          3359 => x"aa",
          3360 => x"87",
          3361 => x"9e",
          3362 => x"87",
          3363 => x"ff",
          3364 => x"53",
          3365 => x"51",
          3366 => x"3f",
          3367 => x"c0",
          3368 => x"29",
          3369 => x"05",
          3370 => x"56",
          3371 => x"2e",
          3372 => x"51",
          3373 => x"3f",
          3374 => x"08",
          3375 => x"34",
          3376 => x"08",
          3377 => x"81",
          3378 => x"52",
          3379 => x"ab",
          3380 => x"1b",
          3381 => x"39",
          3382 => x"74",
          3383 => x"f4",
          3384 => x"ff",
          3385 => x"99",
          3386 => x"2e",
          3387 => x"ae",
          3388 => x"cc",
          3389 => x"80",
          3390 => x"74",
          3391 => x"ba",
          3392 => x"cc",
          3393 => x"e8",
          3394 => x"cc",
          3395 => x"06",
          3396 => x"74",
          3397 => x"ff",
          3398 => x"80",
          3399 => x"84",
          3400 => x"d0",
          3401 => x"56",
          3402 => x"2e",
          3403 => x"51",
          3404 => x"3f",
          3405 => x"08",
          3406 => x"34",
          3407 => x"08",
          3408 => x"81",
          3409 => x"52",
          3410 => x"aa",
          3411 => x"1b",
          3412 => x"ff",
          3413 => x"39",
          3414 => x"e8",
          3415 => x"34",
          3416 => x"53",
          3417 => x"33",
          3418 => x"ed",
          3419 => x"e4",
          3420 => x"ec",
          3421 => x"ff",
          3422 => x"e8",
          3423 => x"54",
          3424 => x"f5",
          3425 => x"14",
          3426 => x"9e",
          3427 => x"1a",
          3428 => x"54",
          3429 => x"f5",
          3430 => x"9e",
          3431 => x"73",
          3432 => x"b0",
          3433 => x"e0",
          3434 => x"9e",
          3435 => x"05",
          3436 => x"9e",
          3437 => x"9c",
          3438 => x"0d",
          3439 => x"79",
          3440 => x"9f",
          3441 => x"70",
          3442 => x"9f",
          3443 => x"74",
          3444 => x"75",
          3445 => x"59",
          3446 => x"54",
          3447 => x"87",
          3448 => x"32",
          3449 => x"87",
          3450 => x"3d",
          3451 => x"3d",
          3452 => x"58",
          3453 => x"76",
          3454 => x"38",
          3455 => x"f5",
          3456 => x"cc",
          3457 => x"12",
          3458 => x"2e",
          3459 => x"51",
          3460 => x"71",
          3461 => x"08",
          3462 => x"52",
          3463 => x"80",
          3464 => x"52",
          3465 => x"80",
          3466 => x"13",
          3467 => x"a0",
          3468 => x"71",
          3469 => x"55",
          3470 => x"72",
          3471 => x"38",
          3472 => x"9f",
          3473 => x"10",
          3474 => x"72",
          3475 => x"9f",
          3476 => x"06",
          3477 => x"75",
          3478 => x"1a",
          3479 => x"5a",
          3480 => x"54",
          3481 => x"74",
          3482 => x"52",
          3483 => x"cc",
          3484 => x"0d",
          3485 => x"0d",
          3486 => x"80",
          3487 => x"30",
          3488 => x"80",
          3489 => x"2b",
          3490 => x"75",
          3491 => x"52",
          3492 => x"80",
          3493 => x"70",
          3494 => x"2b",
          3495 => x"78",
          3496 => x"52",
          3497 => x"81",
          3498 => x"30",
          3499 => x"82",
          3500 => x"31",
          3501 => x"5c",
          3502 => x"7a",
          3503 => x"30",
          3504 => x"10",
          3505 => x"7e",
          3506 => x"81",
          3507 => x"70",
          3508 => x"30",
          3509 => x"06",
          3510 => x"82",
          3511 => x"51",
          3512 => x"41",
          3513 => x"51",
          3514 => x"52",
          3515 => x"54",
          3516 => x"0d",
          3517 => x"0d",
          3518 => x"54",
          3519 => x"54",
          3520 => x"82",
          3521 => x"73",
          3522 => x"31",
          3523 => x"0c",
          3524 => x"0d",
          3525 => x"0d",
          3526 => x"55",
          3527 => x"80",
          3528 => x"75",
          3529 => x"3f",
          3530 => x"08",
          3531 => x"53",
          3532 => x"8d",
          3533 => x"fe",
          3534 => x"82",
          3535 => x"31",
          3536 => x"72",
          3537 => x"c8",
          3538 => x"72",
          3539 => x"c0",
          3540 => x"75",
          3541 => x"72",
          3542 => x"2b",
          3543 => x"53",
          3544 => x"77",
          3545 => x"73",
          3546 => x"2a",
          3547 => x"78",
          3548 => x"31",
          3549 => x"2c",
          3550 => x"7a",
          3551 => x"71",
          3552 => x"5a",
          3553 => x"51",
          3554 => x"72",
          3555 => x"52",
          3556 => x"cc",
          3557 => x"0d",
          3558 => x"0d",
          3559 => x"0b",
          3560 => x"0c",
          3561 => x"82",
          3562 => x"a0",
          3563 => x"52",
          3564 => x"51",
          3565 => x"3f",
          3566 => x"08",
          3567 => x"77",
          3568 => x"57",
          3569 => x"34",
          3570 => x"08",
          3571 => x"15",
          3572 => x"15",
          3573 => x"c4",
          3574 => x"86",
          3575 => x"87",
          3576 => x"87",
          3577 => x"87",
          3578 => x"05",
          3579 => x"07",
          3580 => x"ff",
          3581 => x"2a",
          3582 => x"56",
          3583 => x"34",
          3584 => x"34",
          3585 => x"22",
          3586 => x"82",
          3587 => x"05",
          3588 => x"55",
          3589 => x"15",
          3590 => x"15",
          3591 => x"0d",
          3592 => x"0d",
          3593 => x"51",
          3594 => x"8f",
          3595 => x"83",
          3596 => x"70",
          3597 => x"06",
          3598 => x"70",
          3599 => x"0c",
          3600 => x"04",
          3601 => x"02",
          3602 => x"02",
          3603 => x"05",
          3604 => x"82",
          3605 => x"71",
          3606 => x"11",
          3607 => x"73",
          3608 => x"81",
          3609 => x"88",
          3610 => x"a4",
          3611 => x"22",
          3612 => x"ff",
          3613 => x"88",
          3614 => x"52",
          3615 => x"5b",
          3616 => x"55",
          3617 => x"70",
          3618 => x"82",
          3619 => x"14",
          3620 => x"52",
          3621 => x"15",
          3622 => x"15",
          3623 => x"c4",
          3624 => x"70",
          3625 => x"33",
          3626 => x"07",
          3627 => x"8f",
          3628 => x"51",
          3629 => x"71",
          3630 => x"ff",
          3631 => x"88",
          3632 => x"51",
          3633 => x"34",
          3634 => x"06",
          3635 => x"12",
          3636 => x"c4",
          3637 => x"71",
          3638 => x"81",
          3639 => x"3d",
          3640 => x"3d",
          3641 => x"c4",
          3642 => x"05",
          3643 => x"70",
          3644 => x"11",
          3645 => x"87",
          3646 => x"8b",
          3647 => x"2b",
          3648 => x"59",
          3649 => x"72",
          3650 => x"33",
          3651 => x"71",
          3652 => x"70",
          3653 => x"56",
          3654 => x"84",
          3655 => x"85",
          3656 => x"87",
          3657 => x"14",
          3658 => x"85",
          3659 => x"8b",
          3660 => x"2b",
          3661 => x"57",
          3662 => x"86",
          3663 => x"13",
          3664 => x"2b",
          3665 => x"2a",
          3666 => x"52",
          3667 => x"34",
          3668 => x"34",
          3669 => x"08",
          3670 => x"81",
          3671 => x"88",
          3672 => x"81",
          3673 => x"70",
          3674 => x"51",
          3675 => x"71",
          3676 => x"81",
          3677 => x"3d",
          3678 => x"3d",
          3679 => x"05",
          3680 => x"c4",
          3681 => x"2b",
          3682 => x"33",
          3683 => x"71",
          3684 => x"70",
          3685 => x"70",
          3686 => x"33",
          3687 => x"71",
          3688 => x"53",
          3689 => x"52",
          3690 => x"53",
          3691 => x"25",
          3692 => x"72",
          3693 => x"3f",
          3694 => x"08",
          3695 => x"33",
          3696 => x"71",
          3697 => x"83",
          3698 => x"11",
          3699 => x"12",
          3700 => x"2b",
          3701 => x"2b",
          3702 => x"06",
          3703 => x"51",
          3704 => x"53",
          3705 => x"88",
          3706 => x"72",
          3707 => x"73",
          3708 => x"82",
          3709 => x"70",
          3710 => x"81",
          3711 => x"8b",
          3712 => x"2b",
          3713 => x"57",
          3714 => x"70",
          3715 => x"33",
          3716 => x"07",
          3717 => x"ff",
          3718 => x"2a",
          3719 => x"58",
          3720 => x"34",
          3721 => x"34",
          3722 => x"04",
          3723 => x"82",
          3724 => x"02",
          3725 => x"05",
          3726 => x"2b",
          3727 => x"11",
          3728 => x"33",
          3729 => x"71",
          3730 => x"59",
          3731 => x"56",
          3732 => x"71",
          3733 => x"33",
          3734 => x"07",
          3735 => x"a2",
          3736 => x"07",
          3737 => x"53",
          3738 => x"53",
          3739 => x"70",
          3740 => x"82",
          3741 => x"70",
          3742 => x"81",
          3743 => x"8b",
          3744 => x"2b",
          3745 => x"57",
          3746 => x"82",
          3747 => x"13",
          3748 => x"2b",
          3749 => x"2a",
          3750 => x"52",
          3751 => x"34",
          3752 => x"34",
          3753 => x"08",
          3754 => x"33",
          3755 => x"71",
          3756 => x"82",
          3757 => x"52",
          3758 => x"0d",
          3759 => x"0d",
          3760 => x"c4",
          3761 => x"2a",
          3762 => x"ff",
          3763 => x"57",
          3764 => x"3f",
          3765 => x"08",
          3766 => x"71",
          3767 => x"33",
          3768 => x"71",
          3769 => x"83",
          3770 => x"11",
          3771 => x"12",
          3772 => x"2b",
          3773 => x"07",
          3774 => x"51",
          3775 => x"55",
          3776 => x"80",
          3777 => x"82",
          3778 => x"75",
          3779 => x"3f",
          3780 => x"84",
          3781 => x"15",
          3782 => x"2b",
          3783 => x"07",
          3784 => x"88",
          3785 => x"55",
          3786 => x"86",
          3787 => x"81",
          3788 => x"75",
          3789 => x"82",
          3790 => x"70",
          3791 => x"33",
          3792 => x"71",
          3793 => x"70",
          3794 => x"57",
          3795 => x"72",
          3796 => x"73",
          3797 => x"82",
          3798 => x"18",
          3799 => x"86",
          3800 => x"0b",
          3801 => x"82",
          3802 => x"53",
          3803 => x"34",
          3804 => x"34",
          3805 => x"08",
          3806 => x"81",
          3807 => x"88",
          3808 => x"82",
          3809 => x"70",
          3810 => x"51",
          3811 => x"74",
          3812 => x"81",
          3813 => x"3d",
          3814 => x"3d",
          3815 => x"82",
          3816 => x"84",
          3817 => x"3f",
          3818 => x"86",
          3819 => x"fe",
          3820 => x"3d",
          3821 => x"3d",
          3822 => x"52",
          3823 => x"3f",
          3824 => x"08",
          3825 => x"06",
          3826 => x"08",
          3827 => x"85",
          3828 => x"88",
          3829 => x"5f",
          3830 => x"5a",
          3831 => x"59",
          3832 => x"80",
          3833 => x"88",
          3834 => x"33",
          3835 => x"71",
          3836 => x"70",
          3837 => x"06",
          3838 => x"83",
          3839 => x"70",
          3840 => x"53",
          3841 => x"55",
          3842 => x"8a",
          3843 => x"2e",
          3844 => x"78",
          3845 => x"15",
          3846 => x"33",
          3847 => x"07",
          3848 => x"c2",
          3849 => x"ff",
          3850 => x"38",
          3851 => x"56",
          3852 => x"2b",
          3853 => x"08",
          3854 => x"81",
          3855 => x"88",
          3856 => x"81",
          3857 => x"51",
          3858 => x"5c",
          3859 => x"2e",
          3860 => x"55",
          3861 => x"78",
          3862 => x"38",
          3863 => x"80",
          3864 => x"38",
          3865 => x"09",
          3866 => x"38",
          3867 => x"f2",
          3868 => x"39",
          3869 => x"53",
          3870 => x"51",
          3871 => x"82",
          3872 => x"70",
          3873 => x"33",
          3874 => x"71",
          3875 => x"83",
          3876 => x"5a",
          3877 => x"05",
          3878 => x"83",
          3879 => x"70",
          3880 => x"59",
          3881 => x"84",
          3882 => x"81",
          3883 => x"76",
          3884 => x"82",
          3885 => x"75",
          3886 => x"11",
          3887 => x"11",
          3888 => x"33",
          3889 => x"07",
          3890 => x"53",
          3891 => x"5a",
          3892 => x"86",
          3893 => x"87",
          3894 => x"87",
          3895 => x"1c",
          3896 => x"85",
          3897 => x"8b",
          3898 => x"2b",
          3899 => x"5a",
          3900 => x"54",
          3901 => x"34",
          3902 => x"34",
          3903 => x"08",
          3904 => x"1d",
          3905 => x"85",
          3906 => x"88",
          3907 => x"88",
          3908 => x"5f",
          3909 => x"73",
          3910 => x"75",
          3911 => x"82",
          3912 => x"1b",
          3913 => x"73",
          3914 => x"0c",
          3915 => x"04",
          3916 => x"74",
          3917 => x"c4",
          3918 => x"f4",
          3919 => x"53",
          3920 => x"8b",
          3921 => x"fc",
          3922 => x"87",
          3923 => x"72",
          3924 => x"0c",
          3925 => x"04",
          3926 => x"02",
          3927 => x"51",
          3928 => x"72",
          3929 => x"82",
          3930 => x"33",
          3931 => x"87",
          3932 => x"3d",
          3933 => x"3d",
          3934 => x"05",
          3935 => x"05",
          3936 => x"56",
          3937 => x"72",
          3938 => x"e0",
          3939 => x"2b",
          3940 => x"8c",
          3941 => x"88",
          3942 => x"2e",
          3943 => x"88",
          3944 => x"0c",
          3945 => x"8c",
          3946 => x"71",
          3947 => x"87",
          3948 => x"0c",
          3949 => x"08",
          3950 => x"51",
          3951 => x"2e",
          3952 => x"c0",
          3953 => x"51",
          3954 => x"71",
          3955 => x"80",
          3956 => x"92",
          3957 => x"98",
          3958 => x"70",
          3959 => x"38",
          3960 => x"c8",
          3961 => x"87",
          3962 => x"51",
          3963 => x"cc",
          3964 => x"0d",
          3965 => x"0d",
          3966 => x"02",
          3967 => x"05",
          3968 => x"58",
          3969 => x"52",
          3970 => x"3f",
          3971 => x"08",
          3972 => x"54",
          3973 => x"be",
          3974 => x"75",
          3975 => x"c0",
          3976 => x"87",
          3977 => x"12",
          3978 => x"84",
          3979 => x"40",
          3980 => x"85",
          3981 => x"98",
          3982 => x"7d",
          3983 => x"0c",
          3984 => x"85",
          3985 => x"06",
          3986 => x"71",
          3987 => x"38",
          3988 => x"71",
          3989 => x"05",
          3990 => x"19",
          3991 => x"a2",
          3992 => x"71",
          3993 => x"38",
          3994 => x"83",
          3995 => x"38",
          3996 => x"8a",
          3997 => x"98",
          3998 => x"71",
          3999 => x"c0",
          4000 => x"52",
          4001 => x"87",
          4002 => x"80",
          4003 => x"81",
          4004 => x"c0",
          4005 => x"53",
          4006 => x"82",
          4007 => x"71",
          4008 => x"1a",
          4009 => x"84",
          4010 => x"19",
          4011 => x"06",
          4012 => x"79",
          4013 => x"38",
          4014 => x"80",
          4015 => x"87",
          4016 => x"26",
          4017 => x"73",
          4018 => x"06",
          4019 => x"2e",
          4020 => x"52",
          4021 => x"82",
          4022 => x"8f",
          4023 => x"f3",
          4024 => x"62",
          4025 => x"05",
          4026 => x"57",
          4027 => x"83",
          4028 => x"52",
          4029 => x"3f",
          4030 => x"08",
          4031 => x"54",
          4032 => x"2e",
          4033 => x"81",
          4034 => x"74",
          4035 => x"c0",
          4036 => x"87",
          4037 => x"12",
          4038 => x"84",
          4039 => x"5f",
          4040 => x"0b",
          4041 => x"8c",
          4042 => x"0c",
          4043 => x"80",
          4044 => x"70",
          4045 => x"81",
          4046 => x"54",
          4047 => x"8c",
          4048 => x"81",
          4049 => x"7c",
          4050 => x"58",
          4051 => x"70",
          4052 => x"52",
          4053 => x"8a",
          4054 => x"98",
          4055 => x"71",
          4056 => x"c0",
          4057 => x"52",
          4058 => x"87",
          4059 => x"80",
          4060 => x"81",
          4061 => x"c0",
          4062 => x"53",
          4063 => x"82",
          4064 => x"71",
          4065 => x"19",
          4066 => x"81",
          4067 => x"ff",
          4068 => x"19",
          4069 => x"78",
          4070 => x"38",
          4071 => x"80",
          4072 => x"87",
          4073 => x"26",
          4074 => x"73",
          4075 => x"06",
          4076 => x"2e",
          4077 => x"52",
          4078 => x"82",
          4079 => x"8f",
          4080 => x"fa",
          4081 => x"02",
          4082 => x"05",
          4083 => x"05",
          4084 => x"71",
          4085 => x"57",
          4086 => x"82",
          4087 => x"81",
          4088 => x"54",
          4089 => x"38",
          4090 => x"c0",
          4091 => x"81",
          4092 => x"2e",
          4093 => x"71",
          4094 => x"38",
          4095 => x"87",
          4096 => x"11",
          4097 => x"80",
          4098 => x"80",
          4099 => x"83",
          4100 => x"38",
          4101 => x"72",
          4102 => x"2a",
          4103 => x"51",
          4104 => x"80",
          4105 => x"87",
          4106 => x"08",
          4107 => x"38",
          4108 => x"8c",
          4109 => x"96",
          4110 => x"0c",
          4111 => x"8c",
          4112 => x"08",
          4113 => x"51",
          4114 => x"38",
          4115 => x"56",
          4116 => x"80",
          4117 => x"85",
          4118 => x"77",
          4119 => x"83",
          4120 => x"75",
          4121 => x"87",
          4122 => x"3d",
          4123 => x"3d",
          4124 => x"11",
          4125 => x"71",
          4126 => x"82",
          4127 => x"53",
          4128 => x"0d",
          4129 => x"0d",
          4130 => x"33",
          4131 => x"71",
          4132 => x"88",
          4133 => x"14",
          4134 => x"07",
          4135 => x"33",
          4136 => x"87",
          4137 => x"53",
          4138 => x"52",
          4139 => x"04",
          4140 => x"73",
          4141 => x"92",
          4142 => x"52",
          4143 => x"81",
          4144 => x"70",
          4145 => x"70",
          4146 => x"3d",
          4147 => x"3d",
          4148 => x"52",
          4149 => x"70",
          4150 => x"34",
          4151 => x"51",
          4152 => x"81",
          4153 => x"70",
          4154 => x"70",
          4155 => x"05",
          4156 => x"88",
          4157 => x"72",
          4158 => x"0d",
          4159 => x"0d",
          4160 => x"54",
          4161 => x"80",
          4162 => x"71",
          4163 => x"53",
          4164 => x"81",
          4165 => x"ff",
          4166 => x"39",
          4167 => x"04",
          4168 => x"75",
          4169 => x"52",
          4170 => x"70",
          4171 => x"34",
          4172 => x"70",
          4173 => x"3d",
          4174 => x"3d",
          4175 => x"79",
          4176 => x"74",
          4177 => x"56",
          4178 => x"81",
          4179 => x"71",
          4180 => x"16",
          4181 => x"52",
          4182 => x"86",
          4183 => x"2e",
          4184 => x"82",
          4185 => x"86",
          4186 => x"fe",
          4187 => x"76",
          4188 => x"39",
          4189 => x"8a",
          4190 => x"51",
          4191 => x"71",
          4192 => x"33",
          4193 => x"0c",
          4194 => x"04",
          4195 => x"87",
          4196 => x"80",
          4197 => x"cc",
          4198 => x"3d",
          4199 => x"80",
          4200 => x"33",
          4201 => x"7a",
          4202 => x"38",
          4203 => x"16",
          4204 => x"16",
          4205 => x"17",
          4206 => x"fa",
          4207 => x"87",
          4208 => x"2e",
          4209 => x"b7",
          4210 => x"cc",
          4211 => x"34",
          4212 => x"70",
          4213 => x"31",
          4214 => x"59",
          4215 => x"77",
          4216 => x"82",
          4217 => x"74",
          4218 => x"81",
          4219 => x"81",
          4220 => x"53",
          4221 => x"16",
          4222 => x"e3",
          4223 => x"81",
          4224 => x"87",
          4225 => x"3d",
          4226 => x"3d",
          4227 => x"56",
          4228 => x"74",
          4229 => x"2e",
          4230 => x"51",
          4231 => x"82",
          4232 => x"57",
          4233 => x"08",
          4234 => x"54",
          4235 => x"16",
          4236 => x"33",
          4237 => x"3f",
          4238 => x"08",
          4239 => x"38",
          4240 => x"57",
          4241 => x"0c",
          4242 => x"cc",
          4243 => x"0d",
          4244 => x"0d",
          4245 => x"57",
          4246 => x"82",
          4247 => x"58",
          4248 => x"08",
          4249 => x"76",
          4250 => x"83",
          4251 => x"06",
          4252 => x"84",
          4253 => x"78",
          4254 => x"81",
          4255 => x"38",
          4256 => x"82",
          4257 => x"52",
          4258 => x"52",
          4259 => x"3f",
          4260 => x"52",
          4261 => x"51",
          4262 => x"84",
          4263 => x"d2",
          4264 => x"fc",
          4265 => x"8a",
          4266 => x"52",
          4267 => x"51",
          4268 => x"90",
          4269 => x"84",
          4270 => x"fc",
          4271 => x"17",
          4272 => x"a0",
          4273 => x"86",
          4274 => x"08",
          4275 => x"b0",
          4276 => x"55",
          4277 => x"81",
          4278 => x"f8",
          4279 => x"84",
          4280 => x"53",
          4281 => x"17",
          4282 => x"d7",
          4283 => x"cc",
          4284 => x"83",
          4285 => x"77",
          4286 => x"0c",
          4287 => x"04",
          4288 => x"77",
          4289 => x"12",
          4290 => x"55",
          4291 => x"56",
          4292 => x"8d",
          4293 => x"22",
          4294 => x"ac",
          4295 => x"57",
          4296 => x"87",
          4297 => x"3d",
          4298 => x"3d",
          4299 => x"70",
          4300 => x"57",
          4301 => x"81",
          4302 => x"98",
          4303 => x"81",
          4304 => x"74",
          4305 => x"72",
          4306 => x"f5",
          4307 => x"24",
          4308 => x"81",
          4309 => x"81",
          4310 => x"83",
          4311 => x"38",
          4312 => x"76",
          4313 => x"70",
          4314 => x"16",
          4315 => x"74",
          4316 => x"96",
          4317 => x"cc",
          4318 => x"38",
          4319 => x"06",
          4320 => x"33",
          4321 => x"89",
          4322 => x"08",
          4323 => x"54",
          4324 => x"fc",
          4325 => x"87",
          4326 => x"fe",
          4327 => x"ff",
          4328 => x"11",
          4329 => x"2b",
          4330 => x"81",
          4331 => x"2a",
          4332 => x"51",
          4333 => x"e2",
          4334 => x"ff",
          4335 => x"da",
          4336 => x"2a",
          4337 => x"05",
          4338 => x"fc",
          4339 => x"87",
          4340 => x"c6",
          4341 => x"83",
          4342 => x"05",
          4343 => x"f9",
          4344 => x"87",
          4345 => x"ff",
          4346 => x"ae",
          4347 => x"2a",
          4348 => x"05",
          4349 => x"fc",
          4350 => x"87",
          4351 => x"38",
          4352 => x"83",
          4353 => x"05",
          4354 => x"f8",
          4355 => x"87",
          4356 => x"0a",
          4357 => x"39",
          4358 => x"82",
          4359 => x"89",
          4360 => x"f8",
          4361 => x"7c",
          4362 => x"56",
          4363 => x"77",
          4364 => x"38",
          4365 => x"08",
          4366 => x"38",
          4367 => x"72",
          4368 => x"9d",
          4369 => x"24",
          4370 => x"81",
          4371 => x"82",
          4372 => x"83",
          4373 => x"38",
          4374 => x"76",
          4375 => x"70",
          4376 => x"18",
          4377 => x"76",
          4378 => x"9e",
          4379 => x"cc",
          4380 => x"87",
          4381 => x"d9",
          4382 => x"ff",
          4383 => x"05",
          4384 => x"81",
          4385 => x"54",
          4386 => x"80",
          4387 => x"77",
          4388 => x"f0",
          4389 => x"8f",
          4390 => x"51",
          4391 => x"34",
          4392 => x"17",
          4393 => x"2a",
          4394 => x"05",
          4395 => x"fa",
          4396 => x"87",
          4397 => x"82",
          4398 => x"81",
          4399 => x"83",
          4400 => x"b4",
          4401 => x"2a",
          4402 => x"8f",
          4403 => x"2a",
          4404 => x"f0",
          4405 => x"06",
          4406 => x"72",
          4407 => x"ec",
          4408 => x"2a",
          4409 => x"05",
          4410 => x"fa",
          4411 => x"87",
          4412 => x"82",
          4413 => x"80",
          4414 => x"83",
          4415 => x"52",
          4416 => x"fe",
          4417 => x"b4",
          4418 => x"a4",
          4419 => x"76",
          4420 => x"17",
          4421 => x"75",
          4422 => x"3f",
          4423 => x"08",
          4424 => x"cc",
          4425 => x"77",
          4426 => x"77",
          4427 => x"fc",
          4428 => x"b4",
          4429 => x"51",
          4430 => x"c9",
          4431 => x"cc",
          4432 => x"06",
          4433 => x"72",
          4434 => x"3f",
          4435 => x"17",
          4436 => x"87",
          4437 => x"3d",
          4438 => x"3d",
          4439 => x"7e",
          4440 => x"56",
          4441 => x"75",
          4442 => x"74",
          4443 => x"27",
          4444 => x"80",
          4445 => x"ff",
          4446 => x"75",
          4447 => x"3f",
          4448 => x"08",
          4449 => x"cc",
          4450 => x"38",
          4451 => x"54",
          4452 => x"81",
          4453 => x"39",
          4454 => x"08",
          4455 => x"39",
          4456 => x"51",
          4457 => x"82",
          4458 => x"58",
          4459 => x"08",
          4460 => x"c7",
          4461 => x"cc",
          4462 => x"d2",
          4463 => x"cc",
          4464 => x"cf",
          4465 => x"74",
          4466 => x"fc",
          4467 => x"87",
          4468 => x"38",
          4469 => x"fe",
          4470 => x"08",
          4471 => x"74",
          4472 => x"38",
          4473 => x"17",
          4474 => x"33",
          4475 => x"73",
          4476 => x"77",
          4477 => x"26",
          4478 => x"80",
          4479 => x"87",
          4480 => x"3d",
          4481 => x"3d",
          4482 => x"71",
          4483 => x"5b",
          4484 => x"8c",
          4485 => x"77",
          4486 => x"38",
          4487 => x"78",
          4488 => x"81",
          4489 => x"79",
          4490 => x"f9",
          4491 => x"55",
          4492 => x"cc",
          4493 => x"e0",
          4494 => x"cc",
          4495 => x"87",
          4496 => x"2e",
          4497 => x"98",
          4498 => x"87",
          4499 => x"82",
          4500 => x"58",
          4501 => x"70",
          4502 => x"80",
          4503 => x"38",
          4504 => x"09",
          4505 => x"e2",
          4506 => x"56",
          4507 => x"76",
          4508 => x"82",
          4509 => x"7a",
          4510 => x"3f",
          4511 => x"87",
          4512 => x"2e",
          4513 => x"86",
          4514 => x"cc",
          4515 => x"87",
          4516 => x"70",
          4517 => x"07",
          4518 => x"7c",
          4519 => x"cc",
          4520 => x"51",
          4521 => x"81",
          4522 => x"87",
          4523 => x"2e",
          4524 => x"17",
          4525 => x"74",
          4526 => x"73",
          4527 => x"27",
          4528 => x"58",
          4529 => x"80",
          4530 => x"56",
          4531 => x"98",
          4532 => x"26",
          4533 => x"56",
          4534 => x"81",
          4535 => x"52",
          4536 => x"c6",
          4537 => x"cc",
          4538 => x"b8",
          4539 => x"82",
          4540 => x"81",
          4541 => x"06",
          4542 => x"87",
          4543 => x"82",
          4544 => x"09",
          4545 => x"72",
          4546 => x"70",
          4547 => x"51",
          4548 => x"80",
          4549 => x"78",
          4550 => x"06",
          4551 => x"73",
          4552 => x"39",
          4553 => x"52",
          4554 => x"f7",
          4555 => x"cc",
          4556 => x"cc",
          4557 => x"82",
          4558 => x"07",
          4559 => x"55",
          4560 => x"2e",
          4561 => x"80",
          4562 => x"75",
          4563 => x"76",
          4564 => x"3f",
          4565 => x"08",
          4566 => x"38",
          4567 => x"0c",
          4568 => x"fe",
          4569 => x"08",
          4570 => x"74",
          4571 => x"ff",
          4572 => x"0c",
          4573 => x"81",
          4574 => x"84",
          4575 => x"39",
          4576 => x"81",
          4577 => x"8c",
          4578 => x"8c",
          4579 => x"cc",
          4580 => x"39",
          4581 => x"55",
          4582 => x"cc",
          4583 => x"0d",
          4584 => x"0d",
          4585 => x"55",
          4586 => x"82",
          4587 => x"58",
          4588 => x"87",
          4589 => x"d8",
          4590 => x"74",
          4591 => x"3f",
          4592 => x"08",
          4593 => x"08",
          4594 => x"59",
          4595 => x"77",
          4596 => x"70",
          4597 => x"c8",
          4598 => x"84",
          4599 => x"56",
          4600 => x"58",
          4601 => x"97",
          4602 => x"75",
          4603 => x"52",
          4604 => x"51",
          4605 => x"82",
          4606 => x"80",
          4607 => x"8a",
          4608 => x"32",
          4609 => x"72",
          4610 => x"2a",
          4611 => x"56",
          4612 => x"cc",
          4613 => x"0d",
          4614 => x"0d",
          4615 => x"08",
          4616 => x"74",
          4617 => x"26",
          4618 => x"74",
          4619 => x"72",
          4620 => x"74",
          4621 => x"88",
          4622 => x"73",
          4623 => x"33",
          4624 => x"27",
          4625 => x"16",
          4626 => x"9b",
          4627 => x"2a",
          4628 => x"88",
          4629 => x"58",
          4630 => x"80",
          4631 => x"16",
          4632 => x"0c",
          4633 => x"8a",
          4634 => x"89",
          4635 => x"72",
          4636 => x"38",
          4637 => x"51",
          4638 => x"82",
          4639 => x"54",
          4640 => x"08",
          4641 => x"38",
          4642 => x"87",
          4643 => x"8b",
          4644 => x"08",
          4645 => x"08",
          4646 => x"82",
          4647 => x"74",
          4648 => x"cb",
          4649 => x"75",
          4650 => x"3f",
          4651 => x"08",
          4652 => x"73",
          4653 => x"98",
          4654 => x"82",
          4655 => x"2e",
          4656 => x"39",
          4657 => x"39",
          4658 => x"13",
          4659 => x"74",
          4660 => x"16",
          4661 => x"18",
          4662 => x"77",
          4663 => x"0c",
          4664 => x"04",
          4665 => x"7a",
          4666 => x"12",
          4667 => x"59",
          4668 => x"80",
          4669 => x"86",
          4670 => x"98",
          4671 => x"14",
          4672 => x"55",
          4673 => x"81",
          4674 => x"83",
          4675 => x"77",
          4676 => x"81",
          4677 => x"0c",
          4678 => x"55",
          4679 => x"76",
          4680 => x"17",
          4681 => x"74",
          4682 => x"9b",
          4683 => x"39",
          4684 => x"ff",
          4685 => x"2a",
          4686 => x"81",
          4687 => x"52",
          4688 => x"e6",
          4689 => x"cc",
          4690 => x"55",
          4691 => x"87",
          4692 => x"80",
          4693 => x"55",
          4694 => x"08",
          4695 => x"f4",
          4696 => x"08",
          4697 => x"08",
          4698 => x"38",
          4699 => x"77",
          4700 => x"84",
          4701 => x"39",
          4702 => x"52",
          4703 => x"86",
          4704 => x"cc",
          4705 => x"55",
          4706 => x"08",
          4707 => x"c4",
          4708 => x"82",
          4709 => x"81",
          4710 => x"81",
          4711 => x"cc",
          4712 => x"b0",
          4713 => x"cc",
          4714 => x"51",
          4715 => x"82",
          4716 => x"a0",
          4717 => x"15",
          4718 => x"75",
          4719 => x"3f",
          4720 => x"08",
          4721 => x"76",
          4722 => x"77",
          4723 => x"9c",
          4724 => x"55",
          4725 => x"cc",
          4726 => x"0d",
          4727 => x"0d",
          4728 => x"08",
          4729 => x"80",
          4730 => x"fc",
          4731 => x"87",
          4732 => x"82",
          4733 => x"80",
          4734 => x"87",
          4735 => x"98",
          4736 => x"78",
          4737 => x"3f",
          4738 => x"08",
          4739 => x"cc",
          4740 => x"38",
          4741 => x"08",
          4742 => x"70",
          4743 => x"58",
          4744 => x"2e",
          4745 => x"83",
          4746 => x"82",
          4747 => x"55",
          4748 => x"81",
          4749 => x"07",
          4750 => x"2e",
          4751 => x"16",
          4752 => x"2e",
          4753 => x"88",
          4754 => x"82",
          4755 => x"56",
          4756 => x"51",
          4757 => x"82",
          4758 => x"54",
          4759 => x"08",
          4760 => x"9b",
          4761 => x"2e",
          4762 => x"83",
          4763 => x"73",
          4764 => x"0c",
          4765 => x"04",
          4766 => x"76",
          4767 => x"54",
          4768 => x"82",
          4769 => x"83",
          4770 => x"76",
          4771 => x"53",
          4772 => x"2e",
          4773 => x"90",
          4774 => x"51",
          4775 => x"82",
          4776 => x"90",
          4777 => x"53",
          4778 => x"cc",
          4779 => x"0d",
          4780 => x"0d",
          4781 => x"83",
          4782 => x"54",
          4783 => x"55",
          4784 => x"3f",
          4785 => x"51",
          4786 => x"2e",
          4787 => x"8b",
          4788 => x"2a",
          4789 => x"51",
          4790 => x"86",
          4791 => x"f7",
          4792 => x"7d",
          4793 => x"75",
          4794 => x"98",
          4795 => x"2e",
          4796 => x"98",
          4797 => x"78",
          4798 => x"3f",
          4799 => x"08",
          4800 => x"cc",
          4801 => x"38",
          4802 => x"70",
          4803 => x"73",
          4804 => x"58",
          4805 => x"8b",
          4806 => x"bf",
          4807 => x"ff",
          4808 => x"53",
          4809 => x"34",
          4810 => x"08",
          4811 => x"e5",
          4812 => x"81",
          4813 => x"2e",
          4814 => x"70",
          4815 => x"57",
          4816 => x"9e",
          4817 => x"2e",
          4818 => x"87",
          4819 => x"df",
          4820 => x"72",
          4821 => x"81",
          4822 => x"76",
          4823 => x"2e",
          4824 => x"52",
          4825 => x"fc",
          4826 => x"cc",
          4827 => x"87",
          4828 => x"38",
          4829 => x"fe",
          4830 => x"39",
          4831 => x"16",
          4832 => x"87",
          4833 => x"3d",
          4834 => x"3d",
          4835 => x"08",
          4836 => x"52",
          4837 => x"c5",
          4838 => x"cc",
          4839 => x"87",
          4840 => x"38",
          4841 => x"52",
          4842 => x"de",
          4843 => x"cc",
          4844 => x"87",
          4845 => x"38",
          4846 => x"87",
          4847 => x"9c",
          4848 => x"ea",
          4849 => x"53",
          4850 => x"9c",
          4851 => x"ea",
          4852 => x"0b",
          4853 => x"74",
          4854 => x"0c",
          4855 => x"04",
          4856 => x"75",
          4857 => x"12",
          4858 => x"53",
          4859 => x"9a",
          4860 => x"cc",
          4861 => x"9c",
          4862 => x"e5",
          4863 => x"0b",
          4864 => x"85",
          4865 => x"fa",
          4866 => x"7a",
          4867 => x"0b",
          4868 => x"98",
          4869 => x"2e",
          4870 => x"80",
          4871 => x"55",
          4872 => x"17",
          4873 => x"33",
          4874 => x"51",
          4875 => x"2e",
          4876 => x"85",
          4877 => x"06",
          4878 => x"e5",
          4879 => x"2e",
          4880 => x"8b",
          4881 => x"70",
          4882 => x"34",
          4883 => x"71",
          4884 => x"05",
          4885 => x"15",
          4886 => x"27",
          4887 => x"15",
          4888 => x"80",
          4889 => x"34",
          4890 => x"52",
          4891 => x"88",
          4892 => x"17",
          4893 => x"52",
          4894 => x"3f",
          4895 => x"08",
          4896 => x"12",
          4897 => x"3f",
          4898 => x"08",
          4899 => x"98",
          4900 => x"da",
          4901 => x"cc",
          4902 => x"23",
          4903 => x"04",
          4904 => x"7f",
          4905 => x"5b",
          4906 => x"33",
          4907 => x"73",
          4908 => x"38",
          4909 => x"80",
          4910 => x"38",
          4911 => x"8c",
          4912 => x"08",
          4913 => x"aa",
          4914 => x"41",
          4915 => x"33",
          4916 => x"73",
          4917 => x"81",
          4918 => x"81",
          4919 => x"dc",
          4920 => x"70",
          4921 => x"07",
          4922 => x"73",
          4923 => x"88",
          4924 => x"70",
          4925 => x"73",
          4926 => x"38",
          4927 => x"ab",
          4928 => x"52",
          4929 => x"91",
          4930 => x"cc",
          4931 => x"98",
          4932 => x"61",
          4933 => x"5a",
          4934 => x"a0",
          4935 => x"e7",
          4936 => x"70",
          4937 => x"79",
          4938 => x"73",
          4939 => x"81",
          4940 => x"38",
          4941 => x"33",
          4942 => x"ae",
          4943 => x"70",
          4944 => x"82",
          4945 => x"51",
          4946 => x"54",
          4947 => x"79",
          4948 => x"74",
          4949 => x"57",
          4950 => x"af",
          4951 => x"70",
          4952 => x"51",
          4953 => x"dc",
          4954 => x"73",
          4955 => x"38",
          4956 => x"82",
          4957 => x"19",
          4958 => x"54",
          4959 => x"82",
          4960 => x"54",
          4961 => x"78",
          4962 => x"81",
          4963 => x"54",
          4964 => x"81",
          4965 => x"af",
          4966 => x"77",
          4967 => x"70",
          4968 => x"25",
          4969 => x"07",
          4970 => x"51",
          4971 => x"2e",
          4972 => x"39",
          4973 => x"80",
          4974 => x"33",
          4975 => x"73",
          4976 => x"81",
          4977 => x"81",
          4978 => x"dc",
          4979 => x"70",
          4980 => x"07",
          4981 => x"73",
          4982 => x"b5",
          4983 => x"2e",
          4984 => x"83",
          4985 => x"76",
          4986 => x"07",
          4987 => x"2e",
          4988 => x"8b",
          4989 => x"77",
          4990 => x"30",
          4991 => x"71",
          4992 => x"53",
          4993 => x"55",
          4994 => x"38",
          4995 => x"5c",
          4996 => x"75",
          4997 => x"73",
          4998 => x"38",
          4999 => x"06",
          5000 => x"11",
          5001 => x"75",
          5002 => x"3f",
          5003 => x"08",
          5004 => x"38",
          5005 => x"33",
          5006 => x"54",
          5007 => x"e6",
          5008 => x"87",
          5009 => x"2e",
          5010 => x"ff",
          5011 => x"74",
          5012 => x"38",
          5013 => x"75",
          5014 => x"17",
          5015 => x"57",
          5016 => x"a7",
          5017 => x"82",
          5018 => x"e5",
          5019 => x"87",
          5020 => x"38",
          5021 => x"54",
          5022 => x"89",
          5023 => x"70",
          5024 => x"57",
          5025 => x"54",
          5026 => x"81",
          5027 => x"f7",
          5028 => x"7e",
          5029 => x"2e",
          5030 => x"33",
          5031 => x"e5",
          5032 => x"06",
          5033 => x"7a",
          5034 => x"a0",
          5035 => x"38",
          5036 => x"55",
          5037 => x"84",
          5038 => x"39",
          5039 => x"8b",
          5040 => x"7b",
          5041 => x"7a",
          5042 => x"3f",
          5043 => x"08",
          5044 => x"cc",
          5045 => x"38",
          5046 => x"52",
          5047 => x"aa",
          5048 => x"cc",
          5049 => x"87",
          5050 => x"c2",
          5051 => x"08",
          5052 => x"55",
          5053 => x"ff",
          5054 => x"15",
          5055 => x"54",
          5056 => x"34",
          5057 => x"70",
          5058 => x"81",
          5059 => x"58",
          5060 => x"8b",
          5061 => x"74",
          5062 => x"3f",
          5063 => x"08",
          5064 => x"38",
          5065 => x"51",
          5066 => x"ff",
          5067 => x"ab",
          5068 => x"55",
          5069 => x"bb",
          5070 => x"2e",
          5071 => x"80",
          5072 => x"85",
          5073 => x"06",
          5074 => x"58",
          5075 => x"80",
          5076 => x"75",
          5077 => x"73",
          5078 => x"b5",
          5079 => x"0b",
          5080 => x"80",
          5081 => x"39",
          5082 => x"54",
          5083 => x"85",
          5084 => x"75",
          5085 => x"81",
          5086 => x"73",
          5087 => x"1b",
          5088 => x"2a",
          5089 => x"51",
          5090 => x"80",
          5091 => x"90",
          5092 => x"ff",
          5093 => x"05",
          5094 => x"f5",
          5095 => x"87",
          5096 => x"1c",
          5097 => x"39",
          5098 => x"cc",
          5099 => x"0d",
          5100 => x"0d",
          5101 => x"7b",
          5102 => x"73",
          5103 => x"55",
          5104 => x"2e",
          5105 => x"75",
          5106 => x"57",
          5107 => x"26",
          5108 => x"ba",
          5109 => x"70",
          5110 => x"ba",
          5111 => x"06",
          5112 => x"73",
          5113 => x"70",
          5114 => x"51",
          5115 => x"89",
          5116 => x"82",
          5117 => x"ff",
          5118 => x"56",
          5119 => x"2e",
          5120 => x"80",
          5121 => x"84",
          5122 => x"08",
          5123 => x"76",
          5124 => x"58",
          5125 => x"81",
          5126 => x"ff",
          5127 => x"53",
          5128 => x"26",
          5129 => x"13",
          5130 => x"06",
          5131 => x"9f",
          5132 => x"99",
          5133 => x"e0",
          5134 => x"ff",
          5135 => x"72",
          5136 => x"2a",
          5137 => x"72",
          5138 => x"06",
          5139 => x"ff",
          5140 => x"30",
          5141 => x"70",
          5142 => x"07",
          5143 => x"9f",
          5144 => x"54",
          5145 => x"80",
          5146 => x"81",
          5147 => x"59",
          5148 => x"25",
          5149 => x"8b",
          5150 => x"24",
          5151 => x"76",
          5152 => x"78",
          5153 => x"82",
          5154 => x"51",
          5155 => x"cc",
          5156 => x"0d",
          5157 => x"0d",
          5158 => x"0b",
          5159 => x"ff",
          5160 => x"0c",
          5161 => x"51",
          5162 => x"84",
          5163 => x"cc",
          5164 => x"38",
          5165 => x"51",
          5166 => x"82",
          5167 => x"83",
          5168 => x"54",
          5169 => x"82",
          5170 => x"09",
          5171 => x"e3",
          5172 => x"b4",
          5173 => x"57",
          5174 => x"2e",
          5175 => x"83",
          5176 => x"74",
          5177 => x"70",
          5178 => x"25",
          5179 => x"51",
          5180 => x"38",
          5181 => x"2e",
          5182 => x"b5",
          5183 => x"82",
          5184 => x"80",
          5185 => x"e0",
          5186 => x"87",
          5187 => x"82",
          5188 => x"80",
          5189 => x"85",
          5190 => x"c8",
          5191 => x"16",
          5192 => x"3f",
          5193 => x"08",
          5194 => x"cc",
          5195 => x"83",
          5196 => x"74",
          5197 => x"0c",
          5198 => x"04",
          5199 => x"61",
          5200 => x"80",
          5201 => x"58",
          5202 => x"0c",
          5203 => x"e1",
          5204 => x"cc",
          5205 => x"56",
          5206 => x"87",
          5207 => x"86",
          5208 => x"87",
          5209 => x"29",
          5210 => x"05",
          5211 => x"53",
          5212 => x"80",
          5213 => x"38",
          5214 => x"76",
          5215 => x"74",
          5216 => x"72",
          5217 => x"38",
          5218 => x"51",
          5219 => x"82",
          5220 => x"81",
          5221 => x"81",
          5222 => x"72",
          5223 => x"80",
          5224 => x"38",
          5225 => x"70",
          5226 => x"53",
          5227 => x"86",
          5228 => x"a6",
          5229 => x"34",
          5230 => x"34",
          5231 => x"14",
          5232 => x"b2",
          5233 => x"cc",
          5234 => x"06",
          5235 => x"54",
          5236 => x"72",
          5237 => x"76",
          5238 => x"38",
          5239 => x"70",
          5240 => x"53",
          5241 => x"85",
          5242 => x"70",
          5243 => x"5b",
          5244 => x"82",
          5245 => x"81",
          5246 => x"76",
          5247 => x"81",
          5248 => x"38",
          5249 => x"56",
          5250 => x"83",
          5251 => x"70",
          5252 => x"80",
          5253 => x"83",
          5254 => x"dc",
          5255 => x"87",
          5256 => x"76",
          5257 => x"05",
          5258 => x"16",
          5259 => x"56",
          5260 => x"d7",
          5261 => x"8d",
          5262 => x"72",
          5263 => x"54",
          5264 => x"57",
          5265 => x"95",
          5266 => x"73",
          5267 => x"3f",
          5268 => x"08",
          5269 => x"57",
          5270 => x"89",
          5271 => x"56",
          5272 => x"d7",
          5273 => x"76",
          5274 => x"f0",
          5275 => x"76",
          5276 => x"e8",
          5277 => x"51",
          5278 => x"82",
          5279 => x"83",
          5280 => x"53",
          5281 => x"2e",
          5282 => x"84",
          5283 => x"ca",
          5284 => x"da",
          5285 => x"cc",
          5286 => x"ff",
          5287 => x"8d",
          5288 => x"14",
          5289 => x"3f",
          5290 => x"08",
          5291 => x"15",
          5292 => x"14",
          5293 => x"34",
          5294 => x"33",
          5295 => x"81",
          5296 => x"54",
          5297 => x"72",
          5298 => x"90",
          5299 => x"ff",
          5300 => x"29",
          5301 => x"33",
          5302 => x"72",
          5303 => x"72",
          5304 => x"38",
          5305 => x"06",
          5306 => x"2e",
          5307 => x"56",
          5308 => x"80",
          5309 => x"da",
          5310 => x"87",
          5311 => x"82",
          5312 => x"88",
          5313 => x"8f",
          5314 => x"56",
          5315 => x"38",
          5316 => x"51",
          5317 => x"82",
          5318 => x"83",
          5319 => x"55",
          5320 => x"80",
          5321 => x"da",
          5322 => x"87",
          5323 => x"80",
          5324 => x"da",
          5325 => x"87",
          5326 => x"ff",
          5327 => x"8d",
          5328 => x"2e",
          5329 => x"88",
          5330 => x"14",
          5331 => x"05",
          5332 => x"75",
          5333 => x"38",
          5334 => x"52",
          5335 => x"51",
          5336 => x"82",
          5337 => x"55",
          5338 => x"08",
          5339 => x"ec",
          5340 => x"cc",
          5341 => x"ff",
          5342 => x"83",
          5343 => x"74",
          5344 => x"26",
          5345 => x"57",
          5346 => x"26",
          5347 => x"57",
          5348 => x"56",
          5349 => x"82",
          5350 => x"15",
          5351 => x"0c",
          5352 => x"0c",
          5353 => x"a4",
          5354 => x"1d",
          5355 => x"54",
          5356 => x"2e",
          5357 => x"af",
          5358 => x"14",
          5359 => x"3f",
          5360 => x"08",
          5361 => x"06",
          5362 => x"72",
          5363 => x"79",
          5364 => x"80",
          5365 => x"d9",
          5366 => x"87",
          5367 => x"15",
          5368 => x"2b",
          5369 => x"8d",
          5370 => x"2e",
          5371 => x"77",
          5372 => x"0c",
          5373 => x"76",
          5374 => x"38",
          5375 => x"70",
          5376 => x"81",
          5377 => x"53",
          5378 => x"89",
          5379 => x"56",
          5380 => x"08",
          5381 => x"38",
          5382 => x"15",
          5383 => x"8c",
          5384 => x"80",
          5385 => x"34",
          5386 => x"09",
          5387 => x"92",
          5388 => x"14",
          5389 => x"3f",
          5390 => x"08",
          5391 => x"06",
          5392 => x"2e",
          5393 => x"80",
          5394 => x"1b",
          5395 => x"db",
          5396 => x"87",
          5397 => x"ea",
          5398 => x"cc",
          5399 => x"34",
          5400 => x"51",
          5401 => x"82",
          5402 => x"83",
          5403 => x"53",
          5404 => x"d5",
          5405 => x"06",
          5406 => x"b4",
          5407 => x"85",
          5408 => x"cc",
          5409 => x"85",
          5410 => x"09",
          5411 => x"38",
          5412 => x"51",
          5413 => x"82",
          5414 => x"86",
          5415 => x"f2",
          5416 => x"06",
          5417 => x"9c",
          5418 => x"d9",
          5419 => x"cc",
          5420 => x"0c",
          5421 => x"51",
          5422 => x"82",
          5423 => x"8c",
          5424 => x"74",
          5425 => x"80",
          5426 => x"53",
          5427 => x"80",
          5428 => x"15",
          5429 => x"94",
          5430 => x"56",
          5431 => x"cc",
          5432 => x"0d",
          5433 => x"0d",
          5434 => x"55",
          5435 => x"b9",
          5436 => x"53",
          5437 => x"b1",
          5438 => x"52",
          5439 => x"a9",
          5440 => x"22",
          5441 => x"57",
          5442 => x"2e",
          5443 => x"99",
          5444 => x"33",
          5445 => x"3f",
          5446 => x"08",
          5447 => x"71",
          5448 => x"74",
          5449 => x"83",
          5450 => x"78",
          5451 => x"52",
          5452 => x"cc",
          5453 => x"0d",
          5454 => x"0d",
          5455 => x"33",
          5456 => x"3d",
          5457 => x"56",
          5458 => x"8b",
          5459 => x"82",
          5460 => x"24",
          5461 => x"87",
          5462 => x"29",
          5463 => x"05",
          5464 => x"55",
          5465 => x"84",
          5466 => x"34",
          5467 => x"80",
          5468 => x"80",
          5469 => x"75",
          5470 => x"75",
          5471 => x"38",
          5472 => x"3d",
          5473 => x"05",
          5474 => x"3f",
          5475 => x"08",
          5476 => x"87",
          5477 => x"3d",
          5478 => x"3d",
          5479 => x"84",
          5480 => x"05",
          5481 => x"89",
          5482 => x"2e",
          5483 => x"77",
          5484 => x"54",
          5485 => x"05",
          5486 => x"84",
          5487 => x"f6",
          5488 => x"87",
          5489 => x"82",
          5490 => x"84",
          5491 => x"5c",
          5492 => x"3d",
          5493 => x"ed",
          5494 => x"87",
          5495 => x"82",
          5496 => x"92",
          5497 => x"d7",
          5498 => x"98",
          5499 => x"73",
          5500 => x"38",
          5501 => x"9c",
          5502 => x"80",
          5503 => x"38",
          5504 => x"95",
          5505 => x"2e",
          5506 => x"aa",
          5507 => x"ea",
          5508 => x"87",
          5509 => x"9e",
          5510 => x"05",
          5511 => x"54",
          5512 => x"38",
          5513 => x"70",
          5514 => x"54",
          5515 => x"8e",
          5516 => x"83",
          5517 => x"88",
          5518 => x"83",
          5519 => x"83",
          5520 => x"06",
          5521 => x"80",
          5522 => x"38",
          5523 => x"51",
          5524 => x"82",
          5525 => x"56",
          5526 => x"0a",
          5527 => x"05",
          5528 => x"3f",
          5529 => x"0b",
          5530 => x"80",
          5531 => x"7a",
          5532 => x"3f",
          5533 => x"9c",
          5534 => x"d2",
          5535 => x"81",
          5536 => x"34",
          5537 => x"80",
          5538 => x"b0",
          5539 => x"54",
          5540 => x"52",
          5541 => x"05",
          5542 => x"3f",
          5543 => x"08",
          5544 => x"cc",
          5545 => x"38",
          5546 => x"82",
          5547 => x"b2",
          5548 => x"84",
          5549 => x"06",
          5550 => x"73",
          5551 => x"38",
          5552 => x"ad",
          5553 => x"2a",
          5554 => x"51",
          5555 => x"2e",
          5556 => x"81",
          5557 => x"80",
          5558 => x"87",
          5559 => x"39",
          5560 => x"51",
          5561 => x"82",
          5562 => x"7b",
          5563 => x"12",
          5564 => x"82",
          5565 => x"81",
          5566 => x"83",
          5567 => x"06",
          5568 => x"80",
          5569 => x"77",
          5570 => x"58",
          5571 => x"08",
          5572 => x"63",
          5573 => x"63",
          5574 => x"57",
          5575 => x"82",
          5576 => x"82",
          5577 => x"88",
          5578 => x"9c",
          5579 => x"d2",
          5580 => x"87",
          5581 => x"87",
          5582 => x"1b",
          5583 => x"0c",
          5584 => x"22",
          5585 => x"77",
          5586 => x"80",
          5587 => x"34",
          5588 => x"1a",
          5589 => x"94",
          5590 => x"85",
          5591 => x"06",
          5592 => x"80",
          5593 => x"38",
          5594 => x"08",
          5595 => x"84",
          5596 => x"cc",
          5597 => x"0c",
          5598 => x"70",
          5599 => x"52",
          5600 => x"39",
          5601 => x"51",
          5602 => x"82",
          5603 => x"57",
          5604 => x"08",
          5605 => x"38",
          5606 => x"87",
          5607 => x"2e",
          5608 => x"83",
          5609 => x"75",
          5610 => x"74",
          5611 => x"07",
          5612 => x"54",
          5613 => x"8a",
          5614 => x"75",
          5615 => x"73",
          5616 => x"98",
          5617 => x"a9",
          5618 => x"ff",
          5619 => x"80",
          5620 => x"76",
          5621 => x"d6",
          5622 => x"87",
          5623 => x"38",
          5624 => x"39",
          5625 => x"82",
          5626 => x"05",
          5627 => x"84",
          5628 => x"0c",
          5629 => x"82",
          5630 => x"97",
          5631 => x"f2",
          5632 => x"63",
          5633 => x"40",
          5634 => x"7e",
          5635 => x"fc",
          5636 => x"51",
          5637 => x"82",
          5638 => x"55",
          5639 => x"08",
          5640 => x"19",
          5641 => x"80",
          5642 => x"74",
          5643 => x"39",
          5644 => x"81",
          5645 => x"56",
          5646 => x"82",
          5647 => x"39",
          5648 => x"1a",
          5649 => x"82",
          5650 => x"0b",
          5651 => x"81",
          5652 => x"39",
          5653 => x"94",
          5654 => x"55",
          5655 => x"83",
          5656 => x"7b",
          5657 => x"89",
          5658 => x"08",
          5659 => x"06",
          5660 => x"81",
          5661 => x"8a",
          5662 => x"05",
          5663 => x"06",
          5664 => x"a8",
          5665 => x"38",
          5666 => x"55",
          5667 => x"19",
          5668 => x"51",
          5669 => x"82",
          5670 => x"55",
          5671 => x"ff",
          5672 => x"ff",
          5673 => x"38",
          5674 => x"0c",
          5675 => x"52",
          5676 => x"cc",
          5677 => x"cc",
          5678 => x"ff",
          5679 => x"87",
          5680 => x"7c",
          5681 => x"57",
          5682 => x"80",
          5683 => x"1a",
          5684 => x"22",
          5685 => x"75",
          5686 => x"38",
          5687 => x"58",
          5688 => x"53",
          5689 => x"1b",
          5690 => x"89",
          5691 => x"cc",
          5692 => x"38",
          5693 => x"33",
          5694 => x"80",
          5695 => x"b0",
          5696 => x"31",
          5697 => x"27",
          5698 => x"80",
          5699 => x"52",
          5700 => x"77",
          5701 => x"7d",
          5702 => x"e1",
          5703 => x"2b",
          5704 => x"76",
          5705 => x"94",
          5706 => x"ff",
          5707 => x"71",
          5708 => x"7b",
          5709 => x"38",
          5710 => x"19",
          5711 => x"51",
          5712 => x"82",
          5713 => x"fe",
          5714 => x"53",
          5715 => x"83",
          5716 => x"b4",
          5717 => x"51",
          5718 => x"7b",
          5719 => x"08",
          5720 => x"76",
          5721 => x"08",
          5722 => x"0c",
          5723 => x"f3",
          5724 => x"75",
          5725 => x"0c",
          5726 => x"04",
          5727 => x"60",
          5728 => x"40",
          5729 => x"80",
          5730 => x"3d",
          5731 => x"77",
          5732 => x"3f",
          5733 => x"08",
          5734 => x"cc",
          5735 => x"91",
          5736 => x"74",
          5737 => x"38",
          5738 => x"b8",
          5739 => x"33",
          5740 => x"70",
          5741 => x"56",
          5742 => x"74",
          5743 => x"a4",
          5744 => x"82",
          5745 => x"34",
          5746 => x"98",
          5747 => x"91",
          5748 => x"56",
          5749 => x"94",
          5750 => x"11",
          5751 => x"76",
          5752 => x"75",
          5753 => x"80",
          5754 => x"38",
          5755 => x"70",
          5756 => x"56",
          5757 => x"fd",
          5758 => x"11",
          5759 => x"77",
          5760 => x"5c",
          5761 => x"38",
          5762 => x"88",
          5763 => x"74",
          5764 => x"52",
          5765 => x"18",
          5766 => x"51",
          5767 => x"82",
          5768 => x"55",
          5769 => x"08",
          5770 => x"ab",
          5771 => x"2e",
          5772 => x"74",
          5773 => x"95",
          5774 => x"19",
          5775 => x"08",
          5776 => x"88",
          5777 => x"55",
          5778 => x"9c",
          5779 => x"09",
          5780 => x"38",
          5781 => x"c2",
          5782 => x"cc",
          5783 => x"38",
          5784 => x"52",
          5785 => x"98",
          5786 => x"cc",
          5787 => x"fe",
          5788 => x"87",
          5789 => x"7c",
          5790 => x"57",
          5791 => x"80",
          5792 => x"1b",
          5793 => x"22",
          5794 => x"75",
          5795 => x"38",
          5796 => x"59",
          5797 => x"53",
          5798 => x"1a",
          5799 => x"bf",
          5800 => x"cc",
          5801 => x"38",
          5802 => x"08",
          5803 => x"56",
          5804 => x"9b",
          5805 => x"53",
          5806 => x"77",
          5807 => x"7d",
          5808 => x"16",
          5809 => x"3f",
          5810 => x"0b",
          5811 => x"78",
          5812 => x"80",
          5813 => x"18",
          5814 => x"08",
          5815 => x"7e",
          5816 => x"3f",
          5817 => x"08",
          5818 => x"7e",
          5819 => x"0c",
          5820 => x"19",
          5821 => x"08",
          5822 => x"84",
          5823 => x"57",
          5824 => x"27",
          5825 => x"56",
          5826 => x"52",
          5827 => x"fa",
          5828 => x"cc",
          5829 => x"38",
          5830 => x"52",
          5831 => x"83",
          5832 => x"b4",
          5833 => x"d5",
          5834 => x"81",
          5835 => x"34",
          5836 => x"7e",
          5837 => x"0c",
          5838 => x"1a",
          5839 => x"94",
          5840 => x"1b",
          5841 => x"5e",
          5842 => x"27",
          5843 => x"55",
          5844 => x"0c",
          5845 => x"90",
          5846 => x"c0",
          5847 => x"90",
          5848 => x"56",
          5849 => x"cc",
          5850 => x"0d",
          5851 => x"0d",
          5852 => x"fc",
          5853 => x"52",
          5854 => x"3f",
          5855 => x"08",
          5856 => x"cc",
          5857 => x"38",
          5858 => x"70",
          5859 => x"81",
          5860 => x"55",
          5861 => x"80",
          5862 => x"16",
          5863 => x"51",
          5864 => x"82",
          5865 => x"57",
          5866 => x"08",
          5867 => x"a4",
          5868 => x"11",
          5869 => x"55",
          5870 => x"16",
          5871 => x"08",
          5872 => x"75",
          5873 => x"e9",
          5874 => x"08",
          5875 => x"51",
          5876 => x"82",
          5877 => x"52",
          5878 => x"c9",
          5879 => x"52",
          5880 => x"c9",
          5881 => x"54",
          5882 => x"15",
          5883 => x"cc",
          5884 => x"87",
          5885 => x"17",
          5886 => x"06",
          5887 => x"90",
          5888 => x"82",
          5889 => x"8a",
          5890 => x"fc",
          5891 => x"70",
          5892 => x"d9",
          5893 => x"cc",
          5894 => x"87",
          5895 => x"38",
          5896 => x"05",
          5897 => x"f1",
          5898 => x"87",
          5899 => x"82",
          5900 => x"87",
          5901 => x"cc",
          5902 => x"72",
          5903 => x"0c",
          5904 => x"04",
          5905 => x"84",
          5906 => x"e5",
          5907 => x"80",
          5908 => x"cc",
          5909 => x"38",
          5910 => x"08",
          5911 => x"34",
          5912 => x"82",
          5913 => x"83",
          5914 => x"ef",
          5915 => x"53",
          5916 => x"05",
          5917 => x"51",
          5918 => x"82",
          5919 => x"55",
          5920 => x"08",
          5921 => x"76",
          5922 => x"93",
          5923 => x"51",
          5924 => x"82",
          5925 => x"55",
          5926 => x"08",
          5927 => x"80",
          5928 => x"70",
          5929 => x"56",
          5930 => x"89",
          5931 => x"94",
          5932 => x"b2",
          5933 => x"05",
          5934 => x"2a",
          5935 => x"51",
          5936 => x"80",
          5937 => x"76",
          5938 => x"52",
          5939 => x"3f",
          5940 => x"08",
          5941 => x"8e",
          5942 => x"cc",
          5943 => x"09",
          5944 => x"38",
          5945 => x"82",
          5946 => x"93",
          5947 => x"e4",
          5948 => x"6f",
          5949 => x"7a",
          5950 => x"9e",
          5951 => x"05",
          5952 => x"51",
          5953 => x"82",
          5954 => x"57",
          5955 => x"08",
          5956 => x"7b",
          5957 => x"94",
          5958 => x"55",
          5959 => x"73",
          5960 => x"ed",
          5961 => x"93",
          5962 => x"55",
          5963 => x"82",
          5964 => x"57",
          5965 => x"08",
          5966 => x"68",
          5967 => x"c9",
          5968 => x"87",
          5969 => x"82",
          5970 => x"82",
          5971 => x"52",
          5972 => x"a4",
          5973 => x"cc",
          5974 => x"52",
          5975 => x"b9",
          5976 => x"cc",
          5977 => x"87",
          5978 => x"a2",
          5979 => x"74",
          5980 => x"3f",
          5981 => x"08",
          5982 => x"cc",
          5983 => x"69",
          5984 => x"d9",
          5985 => x"82",
          5986 => x"2e",
          5987 => x"52",
          5988 => x"d0",
          5989 => x"cc",
          5990 => x"87",
          5991 => x"2e",
          5992 => x"84",
          5993 => x"06",
          5994 => x"57",
          5995 => x"76",
          5996 => x"9e",
          5997 => x"05",
          5998 => x"dc",
          5999 => x"90",
          6000 => x"81",
          6001 => x"56",
          6002 => x"80",
          6003 => x"02",
          6004 => x"81",
          6005 => x"70",
          6006 => x"56",
          6007 => x"81",
          6008 => x"78",
          6009 => x"38",
          6010 => x"99",
          6011 => x"81",
          6012 => x"18",
          6013 => x"18",
          6014 => x"58",
          6015 => x"33",
          6016 => x"ee",
          6017 => x"6f",
          6018 => x"af",
          6019 => x"8d",
          6020 => x"2e",
          6021 => x"8a",
          6022 => x"6f",
          6023 => x"af",
          6024 => x"0b",
          6025 => x"33",
          6026 => x"82",
          6027 => x"70",
          6028 => x"52",
          6029 => x"56",
          6030 => x"8d",
          6031 => x"70",
          6032 => x"51",
          6033 => x"f5",
          6034 => x"54",
          6035 => x"a7",
          6036 => x"74",
          6037 => x"38",
          6038 => x"73",
          6039 => x"81",
          6040 => x"81",
          6041 => x"39",
          6042 => x"81",
          6043 => x"74",
          6044 => x"81",
          6045 => x"91",
          6046 => x"6e",
          6047 => x"59",
          6048 => x"7a",
          6049 => x"5c",
          6050 => x"26",
          6051 => x"7a",
          6052 => x"87",
          6053 => x"3d",
          6054 => x"3d",
          6055 => x"8d",
          6056 => x"54",
          6057 => x"55",
          6058 => x"82",
          6059 => x"53",
          6060 => x"08",
          6061 => x"91",
          6062 => x"72",
          6063 => x"8c",
          6064 => x"73",
          6065 => x"38",
          6066 => x"70",
          6067 => x"81",
          6068 => x"57",
          6069 => x"73",
          6070 => x"08",
          6071 => x"94",
          6072 => x"75",
          6073 => x"97",
          6074 => x"11",
          6075 => x"2b",
          6076 => x"73",
          6077 => x"38",
          6078 => x"16",
          6079 => x"ee",
          6080 => x"cc",
          6081 => x"78",
          6082 => x"55",
          6083 => x"de",
          6084 => x"cc",
          6085 => x"96",
          6086 => x"70",
          6087 => x"94",
          6088 => x"71",
          6089 => x"08",
          6090 => x"53",
          6091 => x"15",
          6092 => x"a6",
          6093 => x"74",
          6094 => x"3f",
          6095 => x"08",
          6096 => x"cc",
          6097 => x"81",
          6098 => x"87",
          6099 => x"2e",
          6100 => x"82",
          6101 => x"88",
          6102 => x"98",
          6103 => x"80",
          6104 => x"38",
          6105 => x"80",
          6106 => x"77",
          6107 => x"08",
          6108 => x"0c",
          6109 => x"70",
          6110 => x"81",
          6111 => x"5a",
          6112 => x"2e",
          6113 => x"52",
          6114 => x"fa",
          6115 => x"cc",
          6116 => x"87",
          6117 => x"38",
          6118 => x"08",
          6119 => x"73",
          6120 => x"c7",
          6121 => x"87",
          6122 => x"73",
          6123 => x"38",
          6124 => x"af",
          6125 => x"73",
          6126 => x"27",
          6127 => x"98",
          6128 => x"a0",
          6129 => x"08",
          6130 => x"0c",
          6131 => x"06",
          6132 => x"2e",
          6133 => x"52",
          6134 => x"a4",
          6135 => x"cc",
          6136 => x"82",
          6137 => x"34",
          6138 => x"c4",
          6139 => x"91",
          6140 => x"53",
          6141 => x"89",
          6142 => x"cc",
          6143 => x"94",
          6144 => x"8c",
          6145 => x"27",
          6146 => x"8c",
          6147 => x"15",
          6148 => x"07",
          6149 => x"16",
          6150 => x"ff",
          6151 => x"80",
          6152 => x"77",
          6153 => x"2e",
          6154 => x"9c",
          6155 => x"53",
          6156 => x"cc",
          6157 => x"0d",
          6158 => x"0d",
          6159 => x"54",
          6160 => x"81",
          6161 => x"53",
          6162 => x"05",
          6163 => x"84",
          6164 => x"e8",
          6165 => x"cc",
          6166 => x"87",
          6167 => x"ea",
          6168 => x"0c",
          6169 => x"51",
          6170 => x"82",
          6171 => x"55",
          6172 => x"08",
          6173 => x"ab",
          6174 => x"98",
          6175 => x"80",
          6176 => x"38",
          6177 => x"70",
          6178 => x"81",
          6179 => x"57",
          6180 => x"ad",
          6181 => x"08",
          6182 => x"d3",
          6183 => x"87",
          6184 => x"17",
          6185 => x"86",
          6186 => x"17",
          6187 => x"75",
          6188 => x"3f",
          6189 => x"08",
          6190 => x"2e",
          6191 => x"85",
          6192 => x"86",
          6193 => x"2e",
          6194 => x"76",
          6195 => x"73",
          6196 => x"0c",
          6197 => x"04",
          6198 => x"76",
          6199 => x"05",
          6200 => x"53",
          6201 => x"82",
          6202 => x"87",
          6203 => x"cc",
          6204 => x"86",
          6205 => x"fb",
          6206 => x"79",
          6207 => x"05",
          6208 => x"56",
          6209 => x"3f",
          6210 => x"08",
          6211 => x"cc",
          6212 => x"38",
          6213 => x"82",
          6214 => x"52",
          6215 => x"f9",
          6216 => x"cc",
          6217 => x"ca",
          6218 => x"cc",
          6219 => x"51",
          6220 => x"82",
          6221 => x"53",
          6222 => x"08",
          6223 => x"81",
          6224 => x"80",
          6225 => x"82",
          6226 => x"a6",
          6227 => x"73",
          6228 => x"3f",
          6229 => x"51",
          6230 => x"82",
          6231 => x"84",
          6232 => x"70",
          6233 => x"2c",
          6234 => x"cc",
          6235 => x"51",
          6236 => x"82",
          6237 => x"87",
          6238 => x"ee",
          6239 => x"57",
          6240 => x"3d",
          6241 => x"3d",
          6242 => x"b0",
          6243 => x"cc",
          6244 => x"87",
          6245 => x"38",
          6246 => x"51",
          6247 => x"82",
          6248 => x"55",
          6249 => x"08",
          6250 => x"80",
          6251 => x"70",
          6252 => x"58",
          6253 => x"85",
          6254 => x"8d",
          6255 => x"2e",
          6256 => x"52",
          6257 => x"bf",
          6258 => x"87",
          6259 => x"3d",
          6260 => x"3d",
          6261 => x"55",
          6262 => x"92",
          6263 => x"52",
          6264 => x"de",
          6265 => x"87",
          6266 => x"82",
          6267 => x"82",
          6268 => x"74",
          6269 => x"98",
          6270 => x"11",
          6271 => x"59",
          6272 => x"75",
          6273 => x"38",
          6274 => x"81",
          6275 => x"5b",
          6276 => x"82",
          6277 => x"39",
          6278 => x"08",
          6279 => x"59",
          6280 => x"09",
          6281 => x"38",
          6282 => x"57",
          6283 => x"3d",
          6284 => x"c1",
          6285 => x"87",
          6286 => x"2e",
          6287 => x"87",
          6288 => x"2e",
          6289 => x"87",
          6290 => x"70",
          6291 => x"08",
          6292 => x"7a",
          6293 => x"7f",
          6294 => x"54",
          6295 => x"77",
          6296 => x"80",
          6297 => x"15",
          6298 => x"cc",
          6299 => x"75",
          6300 => x"52",
          6301 => x"52",
          6302 => x"8e",
          6303 => x"cc",
          6304 => x"87",
          6305 => x"d6",
          6306 => x"33",
          6307 => x"1a",
          6308 => x"54",
          6309 => x"09",
          6310 => x"38",
          6311 => x"ff",
          6312 => x"82",
          6313 => x"83",
          6314 => x"70",
          6315 => x"25",
          6316 => x"59",
          6317 => x"9b",
          6318 => x"51",
          6319 => x"3f",
          6320 => x"08",
          6321 => x"70",
          6322 => x"25",
          6323 => x"59",
          6324 => x"75",
          6325 => x"7a",
          6326 => x"ff",
          6327 => x"7c",
          6328 => x"90",
          6329 => x"11",
          6330 => x"56",
          6331 => x"15",
          6332 => x"87",
          6333 => x"3d",
          6334 => x"3d",
          6335 => x"3d",
          6336 => x"70",
          6337 => x"dd",
          6338 => x"cc",
          6339 => x"87",
          6340 => x"a8",
          6341 => x"33",
          6342 => x"a0",
          6343 => x"33",
          6344 => x"70",
          6345 => x"55",
          6346 => x"73",
          6347 => x"8e",
          6348 => x"08",
          6349 => x"18",
          6350 => x"80",
          6351 => x"38",
          6352 => x"08",
          6353 => x"08",
          6354 => x"c4",
          6355 => x"87",
          6356 => x"88",
          6357 => x"80",
          6358 => x"17",
          6359 => x"51",
          6360 => x"3f",
          6361 => x"08",
          6362 => x"81",
          6363 => x"81",
          6364 => x"cc",
          6365 => x"09",
          6366 => x"38",
          6367 => x"39",
          6368 => x"77",
          6369 => x"cc",
          6370 => x"08",
          6371 => x"98",
          6372 => x"82",
          6373 => x"52",
          6374 => x"be",
          6375 => x"cc",
          6376 => x"17",
          6377 => x"0c",
          6378 => x"80",
          6379 => x"73",
          6380 => x"75",
          6381 => x"38",
          6382 => x"34",
          6383 => x"82",
          6384 => x"89",
          6385 => x"e2",
          6386 => x"53",
          6387 => x"a4",
          6388 => x"3d",
          6389 => x"3f",
          6390 => x"08",
          6391 => x"cc",
          6392 => x"38",
          6393 => x"3d",
          6394 => x"3d",
          6395 => x"d1",
          6396 => x"87",
          6397 => x"82",
          6398 => x"81",
          6399 => x"80",
          6400 => x"70",
          6401 => x"81",
          6402 => x"56",
          6403 => x"81",
          6404 => x"98",
          6405 => x"74",
          6406 => x"38",
          6407 => x"05",
          6408 => x"06",
          6409 => x"55",
          6410 => x"38",
          6411 => x"51",
          6412 => x"82",
          6413 => x"74",
          6414 => x"81",
          6415 => x"56",
          6416 => x"80",
          6417 => x"54",
          6418 => x"08",
          6419 => x"2e",
          6420 => x"73",
          6421 => x"cc",
          6422 => x"52",
          6423 => x"52",
          6424 => x"3f",
          6425 => x"08",
          6426 => x"cc",
          6427 => x"38",
          6428 => x"08",
          6429 => x"cc",
          6430 => x"87",
          6431 => x"82",
          6432 => x"86",
          6433 => x"80",
          6434 => x"87",
          6435 => x"2e",
          6436 => x"87",
          6437 => x"c0",
          6438 => x"ce",
          6439 => x"87",
          6440 => x"87",
          6441 => x"70",
          6442 => x"08",
          6443 => x"51",
          6444 => x"80",
          6445 => x"73",
          6446 => x"38",
          6447 => x"52",
          6448 => x"96",
          6449 => x"cc",
          6450 => x"8c",
          6451 => x"ff",
          6452 => x"82",
          6453 => x"55",
          6454 => x"cc",
          6455 => x"0d",
          6456 => x"0d",
          6457 => x"3d",
          6458 => x"9a",
          6459 => x"cc",
          6460 => x"cc",
          6461 => x"87",
          6462 => x"b0",
          6463 => x"69",
          6464 => x"70",
          6465 => x"98",
          6466 => x"cc",
          6467 => x"87",
          6468 => x"38",
          6469 => x"94",
          6470 => x"cc",
          6471 => x"09",
          6472 => x"88",
          6473 => x"df",
          6474 => x"85",
          6475 => x"51",
          6476 => x"74",
          6477 => x"78",
          6478 => x"8a",
          6479 => x"57",
          6480 => x"82",
          6481 => x"75",
          6482 => x"87",
          6483 => x"38",
          6484 => x"87",
          6485 => x"2e",
          6486 => x"83",
          6487 => x"82",
          6488 => x"ff",
          6489 => x"06",
          6490 => x"54",
          6491 => x"73",
          6492 => x"82",
          6493 => x"52",
          6494 => x"a5",
          6495 => x"cc",
          6496 => x"87",
          6497 => x"9a",
          6498 => x"a0",
          6499 => x"51",
          6500 => x"3f",
          6501 => x"0b",
          6502 => x"78",
          6503 => x"bf",
          6504 => x"88",
          6505 => x"80",
          6506 => x"ff",
          6507 => x"75",
          6508 => x"11",
          6509 => x"f9",
          6510 => x"78",
          6511 => x"80",
          6512 => x"ff",
          6513 => x"78",
          6514 => x"80",
          6515 => x"7f",
          6516 => x"d4",
          6517 => x"c9",
          6518 => x"54",
          6519 => x"15",
          6520 => x"cb",
          6521 => x"87",
          6522 => x"82",
          6523 => x"b2",
          6524 => x"b2",
          6525 => x"96",
          6526 => x"b5",
          6527 => x"53",
          6528 => x"51",
          6529 => x"64",
          6530 => x"8b",
          6531 => x"54",
          6532 => x"15",
          6533 => x"ff",
          6534 => x"82",
          6535 => x"54",
          6536 => x"53",
          6537 => x"51",
          6538 => x"3f",
          6539 => x"cc",
          6540 => x"0d",
          6541 => x"0d",
          6542 => x"05",
          6543 => x"3f",
          6544 => x"3d",
          6545 => x"52",
          6546 => x"d5",
          6547 => x"87",
          6548 => x"82",
          6549 => x"82",
          6550 => x"4d",
          6551 => x"52",
          6552 => x"52",
          6553 => x"3f",
          6554 => x"08",
          6555 => x"cc",
          6556 => x"38",
          6557 => x"05",
          6558 => x"06",
          6559 => x"73",
          6560 => x"a0",
          6561 => x"08",
          6562 => x"ff",
          6563 => x"ff",
          6564 => x"ac",
          6565 => x"92",
          6566 => x"54",
          6567 => x"3f",
          6568 => x"52",
          6569 => x"f8",
          6570 => x"cc",
          6571 => x"87",
          6572 => x"38",
          6573 => x"09",
          6574 => x"38",
          6575 => x"08",
          6576 => x"88",
          6577 => x"39",
          6578 => x"08",
          6579 => x"81",
          6580 => x"38",
          6581 => x"b2",
          6582 => x"cc",
          6583 => x"87",
          6584 => x"c8",
          6585 => x"93",
          6586 => x"ff",
          6587 => x"8d",
          6588 => x"b4",
          6589 => x"af",
          6590 => x"17",
          6591 => x"33",
          6592 => x"70",
          6593 => x"55",
          6594 => x"38",
          6595 => x"54",
          6596 => x"34",
          6597 => x"0b",
          6598 => x"8b",
          6599 => x"84",
          6600 => x"06",
          6601 => x"73",
          6602 => x"e5",
          6603 => x"2e",
          6604 => x"75",
          6605 => x"c6",
          6606 => x"87",
          6607 => x"78",
          6608 => x"bc",
          6609 => x"82",
          6610 => x"80",
          6611 => x"38",
          6612 => x"08",
          6613 => x"ff",
          6614 => x"82",
          6615 => x"79",
          6616 => x"58",
          6617 => x"87",
          6618 => x"c0",
          6619 => x"33",
          6620 => x"2e",
          6621 => x"99",
          6622 => x"75",
          6623 => x"c6",
          6624 => x"54",
          6625 => x"15",
          6626 => x"82",
          6627 => x"9c",
          6628 => x"c8",
          6629 => x"87",
          6630 => x"82",
          6631 => x"8c",
          6632 => x"ff",
          6633 => x"82",
          6634 => x"55",
          6635 => x"cc",
          6636 => x"0d",
          6637 => x"0d",
          6638 => x"05",
          6639 => x"05",
          6640 => x"33",
          6641 => x"53",
          6642 => x"05",
          6643 => x"51",
          6644 => x"82",
          6645 => x"55",
          6646 => x"08",
          6647 => x"78",
          6648 => x"95",
          6649 => x"51",
          6650 => x"82",
          6651 => x"55",
          6652 => x"08",
          6653 => x"80",
          6654 => x"81",
          6655 => x"86",
          6656 => x"38",
          6657 => x"61",
          6658 => x"12",
          6659 => x"7a",
          6660 => x"51",
          6661 => x"74",
          6662 => x"78",
          6663 => x"83",
          6664 => x"51",
          6665 => x"3f",
          6666 => x"08",
          6667 => x"87",
          6668 => x"3d",
          6669 => x"3d",
          6670 => x"82",
          6671 => x"d0",
          6672 => x"3d",
          6673 => x"3f",
          6674 => x"08",
          6675 => x"cc",
          6676 => x"38",
          6677 => x"52",
          6678 => x"05",
          6679 => x"3f",
          6680 => x"08",
          6681 => x"cc",
          6682 => x"02",
          6683 => x"33",
          6684 => x"54",
          6685 => x"a6",
          6686 => x"22",
          6687 => x"71",
          6688 => x"53",
          6689 => x"51",
          6690 => x"3f",
          6691 => x"0b",
          6692 => x"76",
          6693 => x"b9",
          6694 => x"cc",
          6695 => x"82",
          6696 => x"93",
          6697 => x"ea",
          6698 => x"6b",
          6699 => x"53",
          6700 => x"05",
          6701 => x"51",
          6702 => x"82",
          6703 => x"82",
          6704 => x"30",
          6705 => x"cc",
          6706 => x"25",
          6707 => x"79",
          6708 => x"85",
          6709 => x"75",
          6710 => x"73",
          6711 => x"f9",
          6712 => x"80",
          6713 => x"8d",
          6714 => x"54",
          6715 => x"3f",
          6716 => x"08",
          6717 => x"cc",
          6718 => x"38",
          6719 => x"51",
          6720 => x"82",
          6721 => x"57",
          6722 => x"08",
          6723 => x"87",
          6724 => x"87",
          6725 => x"5b",
          6726 => x"18",
          6727 => x"18",
          6728 => x"74",
          6729 => x"81",
          6730 => x"78",
          6731 => x"8b",
          6732 => x"54",
          6733 => x"75",
          6734 => x"38",
          6735 => x"1b",
          6736 => x"55",
          6737 => x"2e",
          6738 => x"39",
          6739 => x"09",
          6740 => x"38",
          6741 => x"80",
          6742 => x"70",
          6743 => x"25",
          6744 => x"80",
          6745 => x"38",
          6746 => x"bc",
          6747 => x"11",
          6748 => x"ff",
          6749 => x"82",
          6750 => x"57",
          6751 => x"08",
          6752 => x"70",
          6753 => x"80",
          6754 => x"83",
          6755 => x"80",
          6756 => x"84",
          6757 => x"a7",
          6758 => x"b4",
          6759 => x"ad",
          6760 => x"87",
          6761 => x"0c",
          6762 => x"cc",
          6763 => x"0d",
          6764 => x"0d",
          6765 => x"3d",
          6766 => x"52",
          6767 => x"ce",
          6768 => x"87",
          6769 => x"87",
          6770 => x"54",
          6771 => x"08",
          6772 => x"8b",
          6773 => x"8b",
          6774 => x"59",
          6775 => x"3f",
          6776 => x"33",
          6777 => x"06",
          6778 => x"57",
          6779 => x"81",
          6780 => x"58",
          6781 => x"06",
          6782 => x"4e",
          6783 => x"ff",
          6784 => x"82",
          6785 => x"80",
          6786 => x"6c",
          6787 => x"53",
          6788 => x"ae",
          6789 => x"87",
          6790 => x"2e",
          6791 => x"88",
          6792 => x"6d",
          6793 => x"55",
          6794 => x"87",
          6795 => x"ff",
          6796 => x"83",
          6797 => x"51",
          6798 => x"26",
          6799 => x"15",
          6800 => x"ff",
          6801 => x"80",
          6802 => x"87",
          6803 => x"94",
          6804 => x"74",
          6805 => x"38",
          6806 => x"82",
          6807 => x"ae",
          6808 => x"87",
          6809 => x"38",
          6810 => x"27",
          6811 => x"89",
          6812 => x"8b",
          6813 => x"27",
          6814 => x"55",
          6815 => x"81",
          6816 => x"8f",
          6817 => x"2a",
          6818 => x"70",
          6819 => x"34",
          6820 => x"74",
          6821 => x"05",
          6822 => x"17",
          6823 => x"70",
          6824 => x"52",
          6825 => x"73",
          6826 => x"c8",
          6827 => x"33",
          6828 => x"73",
          6829 => x"81",
          6830 => x"80",
          6831 => x"02",
          6832 => x"76",
          6833 => x"51",
          6834 => x"2e",
          6835 => x"87",
          6836 => x"57",
          6837 => x"79",
          6838 => x"80",
          6839 => x"70",
          6840 => x"ba",
          6841 => x"87",
          6842 => x"82",
          6843 => x"80",
          6844 => x"52",
          6845 => x"bf",
          6846 => x"87",
          6847 => x"82",
          6848 => x"8d",
          6849 => x"c4",
          6850 => x"e5",
          6851 => x"c6",
          6852 => x"cc",
          6853 => x"09",
          6854 => x"cc",
          6855 => x"76",
          6856 => x"c4",
          6857 => x"74",
          6858 => x"b1",
          6859 => x"cc",
          6860 => x"87",
          6861 => x"38",
          6862 => x"87",
          6863 => x"67",
          6864 => x"dc",
          6865 => x"88",
          6866 => x"34",
          6867 => x"52",
          6868 => x"ab",
          6869 => x"54",
          6870 => x"15",
          6871 => x"ff",
          6872 => x"82",
          6873 => x"54",
          6874 => x"82",
          6875 => x"9c",
          6876 => x"f2",
          6877 => x"62",
          6878 => x"80",
          6879 => x"93",
          6880 => x"55",
          6881 => x"5e",
          6882 => x"3f",
          6883 => x"08",
          6884 => x"cc",
          6885 => x"38",
          6886 => x"58",
          6887 => x"38",
          6888 => x"97",
          6889 => x"08",
          6890 => x"38",
          6891 => x"70",
          6892 => x"81",
          6893 => x"55",
          6894 => x"87",
          6895 => x"39",
          6896 => x"90",
          6897 => x"82",
          6898 => x"8a",
          6899 => x"89",
          6900 => x"7f",
          6901 => x"56",
          6902 => x"3f",
          6903 => x"06",
          6904 => x"72",
          6905 => x"82",
          6906 => x"05",
          6907 => x"7c",
          6908 => x"55",
          6909 => x"27",
          6910 => x"16",
          6911 => x"83",
          6912 => x"76",
          6913 => x"80",
          6914 => x"79",
          6915 => x"9a",
          6916 => x"7f",
          6917 => x"14",
          6918 => x"83",
          6919 => x"82",
          6920 => x"81",
          6921 => x"38",
          6922 => x"08",
          6923 => x"95",
          6924 => x"cc",
          6925 => x"81",
          6926 => x"7b",
          6927 => x"06",
          6928 => x"39",
          6929 => x"56",
          6930 => x"09",
          6931 => x"b9",
          6932 => x"80",
          6933 => x"80",
          6934 => x"78",
          6935 => x"7a",
          6936 => x"38",
          6937 => x"73",
          6938 => x"81",
          6939 => x"ff",
          6940 => x"74",
          6941 => x"ff",
          6942 => x"82",
          6943 => x"58",
          6944 => x"08",
          6945 => x"74",
          6946 => x"16",
          6947 => x"73",
          6948 => x"39",
          6949 => x"7e",
          6950 => x"0c",
          6951 => x"2e",
          6952 => x"88",
          6953 => x"8c",
          6954 => x"1a",
          6955 => x"07",
          6956 => x"1b",
          6957 => x"08",
          6958 => x"16",
          6959 => x"75",
          6960 => x"38",
          6961 => x"90",
          6962 => x"15",
          6963 => x"54",
          6964 => x"34",
          6965 => x"82",
          6966 => x"90",
          6967 => x"e9",
          6968 => x"6d",
          6969 => x"80",
          6970 => x"9d",
          6971 => x"5c",
          6972 => x"3f",
          6973 => x"0b",
          6974 => x"08",
          6975 => x"38",
          6976 => x"08",
          6977 => x"9e",
          6978 => x"08",
          6979 => x"80",
          6980 => x"80",
          6981 => x"87",
          6982 => x"ff",
          6983 => x"52",
          6984 => x"a0",
          6985 => x"87",
          6986 => x"ff",
          6987 => x"06",
          6988 => x"56",
          6989 => x"38",
          6990 => x"70",
          6991 => x"55",
          6992 => x"8b",
          6993 => x"3d",
          6994 => x"83",
          6995 => x"ff",
          6996 => x"82",
          6997 => x"99",
          6998 => x"74",
          6999 => x"38",
          7000 => x"80",
          7001 => x"ff",
          7002 => x"55",
          7003 => x"83",
          7004 => x"78",
          7005 => x"38",
          7006 => x"26",
          7007 => x"81",
          7008 => x"8b",
          7009 => x"79",
          7010 => x"80",
          7011 => x"93",
          7012 => x"39",
          7013 => x"6e",
          7014 => x"89",
          7015 => x"48",
          7016 => x"83",
          7017 => x"61",
          7018 => x"25",
          7019 => x"55",
          7020 => x"8a",
          7021 => x"3d",
          7022 => x"81",
          7023 => x"ff",
          7024 => x"81",
          7025 => x"cc",
          7026 => x"38",
          7027 => x"70",
          7028 => x"87",
          7029 => x"56",
          7030 => x"38",
          7031 => x"55",
          7032 => x"75",
          7033 => x"38",
          7034 => x"70",
          7035 => x"ff",
          7036 => x"83",
          7037 => x"78",
          7038 => x"89",
          7039 => x"81",
          7040 => x"06",
          7041 => x"80",
          7042 => x"77",
          7043 => x"74",
          7044 => x"8d",
          7045 => x"06",
          7046 => x"2e",
          7047 => x"77",
          7048 => x"93",
          7049 => x"74",
          7050 => x"cb",
          7051 => x"7d",
          7052 => x"81",
          7053 => x"38",
          7054 => x"66",
          7055 => x"81",
          7056 => x"b8",
          7057 => x"74",
          7058 => x"38",
          7059 => x"98",
          7060 => x"b8",
          7061 => x"82",
          7062 => x"57",
          7063 => x"80",
          7064 => x"76",
          7065 => x"38",
          7066 => x"51",
          7067 => x"3f",
          7068 => x"08",
          7069 => x"87",
          7070 => x"2a",
          7071 => x"5c",
          7072 => x"87",
          7073 => x"80",
          7074 => x"44",
          7075 => x"0a",
          7076 => x"ec",
          7077 => x"39",
          7078 => x"66",
          7079 => x"81",
          7080 => x"a8",
          7081 => x"74",
          7082 => x"38",
          7083 => x"98",
          7084 => x"a8",
          7085 => x"82",
          7086 => x"57",
          7087 => x"80",
          7088 => x"76",
          7089 => x"38",
          7090 => x"51",
          7091 => x"3f",
          7092 => x"08",
          7093 => x"57",
          7094 => x"08",
          7095 => x"96",
          7096 => x"82",
          7097 => x"10",
          7098 => x"08",
          7099 => x"72",
          7100 => x"59",
          7101 => x"ff",
          7102 => x"5d",
          7103 => x"44",
          7104 => x"11",
          7105 => x"70",
          7106 => x"71",
          7107 => x"06",
          7108 => x"52",
          7109 => x"40",
          7110 => x"09",
          7111 => x"38",
          7112 => x"18",
          7113 => x"39",
          7114 => x"79",
          7115 => x"70",
          7116 => x"58",
          7117 => x"76",
          7118 => x"38",
          7119 => x"7d",
          7120 => x"70",
          7121 => x"55",
          7122 => x"3f",
          7123 => x"08",
          7124 => x"2e",
          7125 => x"9b",
          7126 => x"cc",
          7127 => x"f5",
          7128 => x"38",
          7129 => x"38",
          7130 => x"59",
          7131 => x"38",
          7132 => x"7d",
          7133 => x"81",
          7134 => x"38",
          7135 => x"0b",
          7136 => x"08",
          7137 => x"78",
          7138 => x"1a",
          7139 => x"c0",
          7140 => x"74",
          7141 => x"39",
          7142 => x"55",
          7143 => x"8f",
          7144 => x"fd",
          7145 => x"87",
          7146 => x"f5",
          7147 => x"78",
          7148 => x"79",
          7149 => x"80",
          7150 => x"f1",
          7151 => x"39",
          7152 => x"81",
          7153 => x"06",
          7154 => x"55",
          7155 => x"27",
          7156 => x"81",
          7157 => x"56",
          7158 => x"38",
          7159 => x"80",
          7160 => x"ff",
          7161 => x"8b",
          7162 => x"d0",
          7163 => x"ff",
          7164 => x"84",
          7165 => x"1b",
          7166 => x"b4",
          7167 => x"1c",
          7168 => x"ff",
          7169 => x"8e",
          7170 => x"a1",
          7171 => x"0b",
          7172 => x"7d",
          7173 => x"30",
          7174 => x"84",
          7175 => x"51",
          7176 => x"51",
          7177 => x"3f",
          7178 => x"83",
          7179 => x"90",
          7180 => x"ff",
          7181 => x"93",
          7182 => x"a0",
          7183 => x"39",
          7184 => x"1b",
          7185 => x"86",
          7186 => x"95",
          7187 => x"52",
          7188 => x"ff",
          7189 => x"81",
          7190 => x"1b",
          7191 => x"d0",
          7192 => x"9c",
          7193 => x"a0",
          7194 => x"83",
          7195 => x"06",
          7196 => x"82",
          7197 => x"52",
          7198 => x"51",
          7199 => x"3f",
          7200 => x"1b",
          7201 => x"c6",
          7202 => x"ac",
          7203 => x"a0",
          7204 => x"52",
          7205 => x"ff",
          7206 => x"86",
          7207 => x"51",
          7208 => x"3f",
          7209 => x"80",
          7210 => x"a9",
          7211 => x"1c",
          7212 => x"82",
          7213 => x"80",
          7214 => x"ae",
          7215 => x"b2",
          7216 => x"1b",
          7217 => x"86",
          7218 => x"ff",
          7219 => x"96",
          7220 => x"9f",
          7221 => x"80",
          7222 => x"34",
          7223 => x"1c",
          7224 => x"82",
          7225 => x"ab",
          7226 => x"a0",
          7227 => x"d4",
          7228 => x"fe",
          7229 => x"59",
          7230 => x"3f",
          7231 => x"53",
          7232 => x"51",
          7233 => x"3f",
          7234 => x"87",
          7235 => x"e7",
          7236 => x"2e",
          7237 => x"80",
          7238 => x"54",
          7239 => x"53",
          7240 => x"51",
          7241 => x"3f",
          7242 => x"80",
          7243 => x"ff",
          7244 => x"84",
          7245 => x"d2",
          7246 => x"ff",
          7247 => x"86",
          7248 => x"f2",
          7249 => x"1b",
          7250 => x"82",
          7251 => x"52",
          7252 => x"51",
          7253 => x"3f",
          7254 => x"ec",
          7255 => x"9e",
          7256 => x"d4",
          7257 => x"51",
          7258 => x"3f",
          7259 => x"87",
          7260 => x"52",
          7261 => x"9a",
          7262 => x"54",
          7263 => x"7a",
          7264 => x"ff",
          7265 => x"65",
          7266 => x"7a",
          7267 => x"90",
          7268 => x"80",
          7269 => x"2e",
          7270 => x"9a",
          7271 => x"7a",
          7272 => x"aa",
          7273 => x"84",
          7274 => x"9e",
          7275 => x"0a",
          7276 => x"51",
          7277 => x"ff",
          7278 => x"7d",
          7279 => x"38",
          7280 => x"52",
          7281 => x"9e",
          7282 => x"55",
          7283 => x"62",
          7284 => x"74",
          7285 => x"75",
          7286 => x"7e",
          7287 => x"ff",
          7288 => x"cc",
          7289 => x"38",
          7290 => x"82",
          7291 => x"52",
          7292 => x"9e",
          7293 => x"16",
          7294 => x"56",
          7295 => x"38",
          7296 => x"77",
          7297 => x"8d",
          7298 => x"7d",
          7299 => x"38",
          7300 => x"57",
          7301 => x"83",
          7302 => x"76",
          7303 => x"7a",
          7304 => x"ff",
          7305 => x"82",
          7306 => x"81",
          7307 => x"16",
          7308 => x"56",
          7309 => x"38",
          7310 => x"83",
          7311 => x"86",
          7312 => x"ff",
          7313 => x"38",
          7314 => x"82",
          7315 => x"81",
          7316 => x"06",
          7317 => x"fe",
          7318 => x"53",
          7319 => x"51",
          7320 => x"3f",
          7321 => x"52",
          7322 => x"9c",
          7323 => x"be",
          7324 => x"75",
          7325 => x"81",
          7326 => x"0b",
          7327 => x"77",
          7328 => x"75",
          7329 => x"60",
          7330 => x"80",
          7331 => x"75",
          7332 => x"da",
          7333 => x"85",
          7334 => x"87",
          7335 => x"2a",
          7336 => x"75",
          7337 => x"82",
          7338 => x"87",
          7339 => x"52",
          7340 => x"51",
          7341 => x"3f",
          7342 => x"ca",
          7343 => x"9c",
          7344 => x"54",
          7345 => x"52",
          7346 => x"98",
          7347 => x"56",
          7348 => x"08",
          7349 => x"53",
          7350 => x"51",
          7351 => x"3f",
          7352 => x"87",
          7353 => x"38",
          7354 => x"56",
          7355 => x"56",
          7356 => x"87",
          7357 => x"75",
          7358 => x"0c",
          7359 => x"04",
          7360 => x"7d",
          7361 => x"80",
          7362 => x"05",
          7363 => x"76",
          7364 => x"38",
          7365 => x"11",
          7366 => x"53",
          7367 => x"79",
          7368 => x"3f",
          7369 => x"09",
          7370 => x"38",
          7371 => x"55",
          7372 => x"db",
          7373 => x"70",
          7374 => x"34",
          7375 => x"74",
          7376 => x"81",
          7377 => x"80",
          7378 => x"55",
          7379 => x"76",
          7380 => x"87",
          7381 => x"3d",
          7382 => x"3d",
          7383 => x"84",
          7384 => x"33",
          7385 => x"8a",
          7386 => x"06",
          7387 => x"52",
          7388 => x"3f",
          7389 => x"56",
          7390 => x"be",
          7391 => x"08",
          7392 => x"05",
          7393 => x"75",
          7394 => x"56",
          7395 => x"a1",
          7396 => x"fc",
          7397 => x"53",
          7398 => x"76",
          7399 => x"dc",
          7400 => x"32",
          7401 => x"72",
          7402 => x"70",
          7403 => x"56",
          7404 => x"18",
          7405 => x"88",
          7406 => x"3d",
          7407 => x"3d",
          7408 => x"11",
          7409 => x"80",
          7410 => x"38",
          7411 => x"05",
          7412 => x"8c",
          7413 => x"08",
          7414 => x"3f",
          7415 => x"08",
          7416 => x"16",
          7417 => x"09",
          7418 => x"38",
          7419 => x"55",
          7420 => x"55",
          7421 => x"cc",
          7422 => x"0d",
          7423 => x"0d",
          7424 => x"cc",
          7425 => x"73",
          7426 => x"94",
          7427 => x"0c",
          7428 => x"04",
          7429 => x"02",
          7430 => x"33",
          7431 => x"3d",
          7432 => x"54",
          7433 => x"52",
          7434 => x"ae",
          7435 => x"ff",
          7436 => x"3d",
          7437 => x"00",
          7438 => x"ff",
          7439 => x"ff",
          7440 => x"ff",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"00",
          7471 => x"00",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"00",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"00",
          7480 => x"00",
          7481 => x"00",
          7482 => x"00",
          7483 => x"00",
          7484 => x"00",
          7485 => x"00",
          7486 => x"00",
          7487 => x"00",
          7488 => x"64",
          7489 => x"74",
          7490 => x"64",
          7491 => x"74",
          7492 => x"66",
          7493 => x"74",
          7494 => x"66",
          7495 => x"64",
          7496 => x"66",
          7497 => x"63",
          7498 => x"6d",
          7499 => x"61",
          7500 => x"6d",
          7501 => x"79",
          7502 => x"6d",
          7503 => x"66",
          7504 => x"6d",
          7505 => x"70",
          7506 => x"6d",
          7507 => x"6d",
          7508 => x"6d",
          7509 => x"68",
          7510 => x"68",
          7511 => x"68",
          7512 => x"68",
          7513 => x"63",
          7514 => x"00",
          7515 => x"6a",
          7516 => x"72",
          7517 => x"61",
          7518 => x"72",
          7519 => x"74",
          7520 => x"69",
          7521 => x"00",
          7522 => x"74",
          7523 => x"00",
          7524 => x"74",
          7525 => x"69",
          7526 => x"6d",
          7527 => x"69",
          7528 => x"6b",
          7529 => x"00",
          7530 => x"65",
          7531 => x"44",
          7532 => x"20",
          7533 => x"6f",
          7534 => x"49",
          7535 => x"72",
          7536 => x"20",
          7537 => x"6f",
          7538 => x"00",
          7539 => x"44",
          7540 => x"20",
          7541 => x"20",
          7542 => x"64",
          7543 => x"00",
          7544 => x"4e",
          7545 => x"69",
          7546 => x"66",
          7547 => x"64",
          7548 => x"4e",
          7549 => x"61",
          7550 => x"66",
          7551 => x"64",
          7552 => x"49",
          7553 => x"6c",
          7554 => x"66",
          7555 => x"6e",
          7556 => x"2e",
          7557 => x"41",
          7558 => x"73",
          7559 => x"65",
          7560 => x"64",
          7561 => x"46",
          7562 => x"20",
          7563 => x"65",
          7564 => x"20",
          7565 => x"73",
          7566 => x"0a",
          7567 => x"46",
          7568 => x"20",
          7569 => x"64",
          7570 => x"69",
          7571 => x"6c",
          7572 => x"0a",
          7573 => x"53",
          7574 => x"73",
          7575 => x"69",
          7576 => x"70",
          7577 => x"65",
          7578 => x"64",
          7579 => x"44",
          7580 => x"65",
          7581 => x"6d",
          7582 => x"20",
          7583 => x"69",
          7584 => x"6c",
          7585 => x"0a",
          7586 => x"44",
          7587 => x"20",
          7588 => x"20",
          7589 => x"62",
          7590 => x"2e",
          7591 => x"4e",
          7592 => x"6f",
          7593 => x"74",
          7594 => x"65",
          7595 => x"6c",
          7596 => x"73",
          7597 => x"20",
          7598 => x"6e",
          7599 => x"6e",
          7600 => x"73",
          7601 => x"00",
          7602 => x"46",
          7603 => x"61",
          7604 => x"62",
          7605 => x"65",
          7606 => x"00",
          7607 => x"54",
          7608 => x"6f",
          7609 => x"20",
          7610 => x"72",
          7611 => x"6f",
          7612 => x"61",
          7613 => x"6c",
          7614 => x"2e",
          7615 => x"46",
          7616 => x"20",
          7617 => x"6c",
          7618 => x"65",
          7619 => x"00",
          7620 => x"49",
          7621 => x"66",
          7622 => x"69",
          7623 => x"20",
          7624 => x"6f",
          7625 => x"0a",
          7626 => x"54",
          7627 => x"6d",
          7628 => x"20",
          7629 => x"6e",
          7630 => x"6c",
          7631 => x"0a",
          7632 => x"50",
          7633 => x"6d",
          7634 => x"72",
          7635 => x"6e",
          7636 => x"72",
          7637 => x"2e",
          7638 => x"53",
          7639 => x"65",
          7640 => x"0a",
          7641 => x"55",
          7642 => x"6f",
          7643 => x"65",
          7644 => x"72",
          7645 => x"0a",
          7646 => x"20",
          7647 => x"65",
          7648 => x"73",
          7649 => x"20",
          7650 => x"20",
          7651 => x"65",
          7652 => x"65",
          7653 => x"00",
          7654 => x"72",
          7655 => x"00",
          7656 => x"25",
          7657 => x"00",
          7658 => x"3a",
          7659 => x"25",
          7660 => x"00",
          7661 => x"20",
          7662 => x"20",
          7663 => x"00",
          7664 => x"25",
          7665 => x"00",
          7666 => x"20",
          7667 => x"20",
          7668 => x"7c",
          7669 => x"5a",
          7670 => x"41",
          7671 => x"0a",
          7672 => x"25",
          7673 => x"00",
          7674 => x"30",
          7675 => x"35",
          7676 => x"32",
          7677 => x"76",
          7678 => x"32",
          7679 => x"20",
          7680 => x"2c",
          7681 => x"76",
          7682 => x"32",
          7683 => x"25",
          7684 => x"73",
          7685 => x"0a",
          7686 => x"5a",
          7687 => x"41",
          7688 => x"74",
          7689 => x"75",
          7690 => x"48",
          7691 => x"6c",
          7692 => x"00",
          7693 => x"54",
          7694 => x"72",
          7695 => x"74",
          7696 => x"75",
          7697 => x"00",
          7698 => x"50",
          7699 => x"69",
          7700 => x"72",
          7701 => x"74",
          7702 => x"49",
          7703 => x"4c",
          7704 => x"20",
          7705 => x"65",
          7706 => x"70",
          7707 => x"49",
          7708 => x"4c",
          7709 => x"20",
          7710 => x"65",
          7711 => x"70",
          7712 => x"55",
          7713 => x"30",
          7714 => x"20",
          7715 => x"65",
          7716 => x"70",
          7717 => x"55",
          7718 => x"30",
          7719 => x"20",
          7720 => x"65",
          7721 => x"70",
          7722 => x"55",
          7723 => x"31",
          7724 => x"20",
          7725 => x"65",
          7726 => x"70",
          7727 => x"55",
          7728 => x"31",
          7729 => x"20",
          7730 => x"65",
          7731 => x"70",
          7732 => x"53",
          7733 => x"69",
          7734 => x"75",
          7735 => x"69",
          7736 => x"2e",
          7737 => x"00",
          7738 => x"45",
          7739 => x"6c",
          7740 => x"20",
          7741 => x"65",
          7742 => x"2e",
          7743 => x"61",
          7744 => x"65",
          7745 => x"2e",
          7746 => x"00",
          7747 => x"7a",
          7748 => x"61",
          7749 => x"74",
          7750 => x"30",
          7751 => x"46",
          7752 => x"65",
          7753 => x"6f",
          7754 => x"69",
          7755 => x"6c",
          7756 => x"20",
          7757 => x"63",
          7758 => x"20",
          7759 => x"70",
          7760 => x"73",
          7761 => x"6e",
          7762 => x"6d",
          7763 => x"61",
          7764 => x"2e",
          7765 => x"2a",
          7766 => x"42",
          7767 => x"64",
          7768 => x"20",
          7769 => x"0a",
          7770 => x"49",
          7771 => x"69",
          7772 => x"73",
          7773 => x"0a",
          7774 => x"46",
          7775 => x"65",
          7776 => x"6f",
          7777 => x"69",
          7778 => x"6c",
          7779 => x"2e",
          7780 => x"72",
          7781 => x"64",
          7782 => x"25",
          7783 => x"43",
          7784 => x"72",
          7785 => x"2e",
          7786 => x"00",
          7787 => x"43",
          7788 => x"69",
          7789 => x"2e",
          7790 => x"43",
          7791 => x"61",
          7792 => x"67",
          7793 => x"00",
          7794 => x"25",
          7795 => x"78",
          7796 => x"38",
          7797 => x"3e",
          7798 => x"6c",
          7799 => x"30",
          7800 => x"0a",
          7801 => x"44",
          7802 => x"20",
          7803 => x"6f",
          7804 => x"00",
          7805 => x"0a",
          7806 => x"70",
          7807 => x"65",
          7808 => x"25",
          7809 => x"20",
          7810 => x"58",
          7811 => x"3f",
          7812 => x"00",
          7813 => x"25",
          7814 => x"20",
          7815 => x"58",
          7816 => x"25",
          7817 => x"20",
          7818 => x"58",
          7819 => x"44",
          7820 => x"62",
          7821 => x"67",
          7822 => x"74",
          7823 => x"75",
          7824 => x"0a",
          7825 => x"45",
          7826 => x"6c",
          7827 => x"20",
          7828 => x"65",
          7829 => x"70",
          7830 => x"00",
          7831 => x"44",
          7832 => x"62",
          7833 => x"20",
          7834 => x"74",
          7835 => x"66",
          7836 => x"45",
          7837 => x"6c",
          7838 => x"20",
          7839 => x"74",
          7840 => x"66",
          7841 => x"45",
          7842 => x"75",
          7843 => x"67",
          7844 => x"64",
          7845 => x"20",
          7846 => x"78",
          7847 => x"2e",
          7848 => x"43",
          7849 => x"69",
          7850 => x"63",
          7851 => x"20",
          7852 => x"30",
          7853 => x"2e",
          7854 => x"00",
          7855 => x"43",
          7856 => x"20",
          7857 => x"75",
          7858 => x"64",
          7859 => x"64",
          7860 => x"25",
          7861 => x"0a",
          7862 => x"52",
          7863 => x"61",
          7864 => x"6e",
          7865 => x"70",
          7866 => x"63",
          7867 => x"6f",
          7868 => x"2e",
          7869 => x"43",
          7870 => x"20",
          7871 => x"6f",
          7872 => x"6e",
          7873 => x"2e",
          7874 => x"5a",
          7875 => x"62",
          7876 => x"25",
          7877 => x"25",
          7878 => x"73",
          7879 => x"00",
          7880 => x"25",
          7881 => x"25",
          7882 => x"73",
          7883 => x"25",
          7884 => x"25",
          7885 => x"42",
          7886 => x"63",
          7887 => x"61",
          7888 => x"0a",
          7889 => x"52",
          7890 => x"69",
          7891 => x"2e",
          7892 => x"45",
          7893 => x"6c",
          7894 => x"20",
          7895 => x"65",
          7896 => x"70",
          7897 => x"2e",
          7898 => x"25",
          7899 => x"64",
          7900 => x"20",
          7901 => x"25",
          7902 => x"64",
          7903 => x"25",
          7904 => x"53",
          7905 => x"43",
          7906 => x"69",
          7907 => x"61",
          7908 => x"6e",
          7909 => x"20",
          7910 => x"6f",
          7911 => x"6f",
          7912 => x"6f",
          7913 => x"67",
          7914 => x"3a",
          7915 => x"76",
          7916 => x"73",
          7917 => x"70",
          7918 => x"65",
          7919 => x"64",
          7920 => x"20",
          7921 => x"57",
          7922 => x"44",
          7923 => x"20",
          7924 => x"30",
          7925 => x"25",
          7926 => x"29",
          7927 => x"20",
          7928 => x"53",
          7929 => x"4d",
          7930 => x"20",
          7931 => x"30",
          7932 => x"25",
          7933 => x"29",
          7934 => x"20",
          7935 => x"49",
          7936 => x"20",
          7937 => x"4d",
          7938 => x"30",
          7939 => x"25",
          7940 => x"29",
          7941 => x"20",
          7942 => x"42",
          7943 => x"20",
          7944 => x"20",
          7945 => x"30",
          7946 => x"25",
          7947 => x"29",
          7948 => x"20",
          7949 => x"52",
          7950 => x"20",
          7951 => x"20",
          7952 => x"30",
          7953 => x"25",
          7954 => x"29",
          7955 => x"20",
          7956 => x"53",
          7957 => x"41",
          7958 => x"20",
          7959 => x"65",
          7960 => x"65",
          7961 => x"25",
          7962 => x"29",
          7963 => x"20",
          7964 => x"54",
          7965 => x"52",
          7966 => x"20",
          7967 => x"69",
          7968 => x"73",
          7969 => x"25",
          7970 => x"29",
          7971 => x"20",
          7972 => x"49",
          7973 => x"20",
          7974 => x"4c",
          7975 => x"68",
          7976 => x"65",
          7977 => x"25",
          7978 => x"29",
          7979 => x"20",
          7980 => x"57",
          7981 => x"42",
          7982 => x"20",
          7983 => x"0a",
          7984 => x"20",
          7985 => x"57",
          7986 => x"32",
          7987 => x"20",
          7988 => x"49",
          7989 => x"4c",
          7990 => x"20",
          7991 => x"50",
          7992 => x"00",
          7993 => x"20",
          7994 => x"53",
          7995 => x"00",
          7996 => x"41",
          7997 => x"65",
          7998 => x"73",
          7999 => x"20",
          8000 => x"43",
          8001 => x"52",
          8002 => x"74",
          8003 => x"63",
          8004 => x"20",
          8005 => x"72",
          8006 => x"20",
          8007 => x"30",
          8008 => x"00",
          8009 => x"20",
          8010 => x"43",
          8011 => x"4d",
          8012 => x"72",
          8013 => x"74",
          8014 => x"20",
          8015 => x"72",
          8016 => x"20",
          8017 => x"30",
          8018 => x"00",
          8019 => x"20",
          8020 => x"53",
          8021 => x"6b",
          8022 => x"61",
          8023 => x"41",
          8024 => x"65",
          8025 => x"20",
          8026 => x"20",
          8027 => x"30",
          8028 => x"00",
          8029 => x"4d",
          8030 => x"3a",
          8031 => x"20",
          8032 => x"5a",
          8033 => x"49",
          8034 => x"20",
          8035 => x"20",
          8036 => x"20",
          8037 => x"20",
          8038 => x"20",
          8039 => x"30",
          8040 => x"00",
          8041 => x"20",
          8042 => x"53",
          8043 => x"65",
          8044 => x"6c",
          8045 => x"20",
          8046 => x"71",
          8047 => x"20",
          8048 => x"20",
          8049 => x"64",
          8050 => x"34",
          8051 => x"7a",
          8052 => x"20",
          8053 => x"53",
          8054 => x"4d",
          8055 => x"6f",
          8056 => x"46",
          8057 => x"20",
          8058 => x"20",
          8059 => x"20",
          8060 => x"64",
          8061 => x"34",
          8062 => x"7a",
          8063 => x"20",
          8064 => x"57",
          8065 => x"62",
          8066 => x"20",
          8067 => x"41",
          8068 => x"6c",
          8069 => x"20",
          8070 => x"71",
          8071 => x"64",
          8072 => x"34",
          8073 => x"7a",
          8074 => x"53",
          8075 => x"6c",
          8076 => x"4d",
          8077 => x"75",
          8078 => x"46",
          8079 => x"00",
          8080 => x"45",
          8081 => x"45",
          8082 => x"69",
          8083 => x"55",
          8084 => x"6f",
          8085 => x"00",
          8086 => x"01",
          8087 => x"00",
          8088 => x"00",
          8089 => x"01",
          8090 => x"00",
          8091 => x"00",
          8092 => x"01",
          8093 => x"00",
          8094 => x"00",
          8095 => x"01",
          8096 => x"00",
          8097 => x"00",
          8098 => x"01",
          8099 => x"00",
          8100 => x"00",
          8101 => x"01",
          8102 => x"00",
          8103 => x"00",
          8104 => x"01",
          8105 => x"00",
          8106 => x"00",
          8107 => x"01",
          8108 => x"00",
          8109 => x"00",
          8110 => x"01",
          8111 => x"00",
          8112 => x"00",
          8113 => x"01",
          8114 => x"00",
          8115 => x"00",
          8116 => x"01",
          8117 => x"00",
          8118 => x"00",
          8119 => x"04",
          8120 => x"00",
          8121 => x"00",
          8122 => x"04",
          8123 => x"00",
          8124 => x"00",
          8125 => x"04",
          8126 => x"00",
          8127 => x"00",
          8128 => x"03",
          8129 => x"00",
          8130 => x"00",
          8131 => x"04",
          8132 => x"00",
          8133 => x"00",
          8134 => x"04",
          8135 => x"00",
          8136 => x"00",
          8137 => x"04",
          8138 => x"00",
          8139 => x"00",
          8140 => x"03",
          8141 => x"00",
          8142 => x"00",
          8143 => x"03",
          8144 => x"00",
          8145 => x"00",
          8146 => x"03",
          8147 => x"00",
          8148 => x"00",
          8149 => x"03",
          8150 => x"00",
          8151 => x"1b",
          8152 => x"1b",
          8153 => x"1b",
          8154 => x"1b",
          8155 => x"1b",
          8156 => x"1b",
          8157 => x"1b",
          8158 => x"1b",
          8159 => x"1b",
          8160 => x"1b",
          8161 => x"1b",
          8162 => x"10",
          8163 => x"0e",
          8164 => x"0d",
          8165 => x"0b",
          8166 => x"08",
          8167 => x"06",
          8168 => x"05",
          8169 => x"04",
          8170 => x"03",
          8171 => x"02",
          8172 => x"01",
          8173 => x"68",
          8174 => x"6f",
          8175 => x"68",
          8176 => x"00",
          8177 => x"21",
          8178 => x"25",
          8179 => x"20",
          8180 => x"0a",
          8181 => x"46",
          8182 => x"65",
          8183 => x"6f",
          8184 => x"73",
          8185 => x"74",
          8186 => x"68",
          8187 => x"6f",
          8188 => x"66",
          8189 => x"20",
          8190 => x"45",
          8191 => x"0a",
          8192 => x"43",
          8193 => x"6f",
          8194 => x"70",
          8195 => x"63",
          8196 => x"74",
          8197 => x"69",
          8198 => x"72",
          8199 => x"69",
          8200 => x"20",
          8201 => x"61",
          8202 => x"6e",
          8203 => x"00",
          8204 => x"53",
          8205 => x"22",
          8206 => x"3a",
          8207 => x"3e",
          8208 => x"7c",
          8209 => x"46",
          8210 => x"46",
          8211 => x"32",
          8212 => x"eb",
          8213 => x"53",
          8214 => x"35",
          8215 => x"4e",
          8216 => x"41",
          8217 => x"20",
          8218 => x"41",
          8219 => x"20",
          8220 => x"4e",
          8221 => x"41",
          8222 => x"20",
          8223 => x"41",
          8224 => x"20",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"80",
          8230 => x"8e",
          8231 => x"45",
          8232 => x"49",
          8233 => x"90",
          8234 => x"99",
          8235 => x"59",
          8236 => x"9c",
          8237 => x"41",
          8238 => x"a5",
          8239 => x"a8",
          8240 => x"ac",
          8241 => x"b0",
          8242 => x"b4",
          8243 => x"b8",
          8244 => x"bc",
          8245 => x"c0",
          8246 => x"c4",
          8247 => x"c8",
          8248 => x"cc",
          8249 => x"d0",
          8250 => x"d4",
          8251 => x"d8",
          8252 => x"dc",
          8253 => x"e0",
          8254 => x"e4",
          8255 => x"e8",
          8256 => x"ec",
          8257 => x"f0",
          8258 => x"f4",
          8259 => x"f8",
          8260 => x"fc",
          8261 => x"2b",
          8262 => x"3d",
          8263 => x"5c",
          8264 => x"3c",
          8265 => x"7f",
          8266 => x"00",
          8267 => x"00",
          8268 => x"01",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"01",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"01",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"01",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"01",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"01",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"01",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"01",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"01",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"01",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"01",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"01",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"01",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"01",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"01",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"01",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"01",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"01",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"01",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"01",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"01",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"01",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"01",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"01",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"01",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"01",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"01",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"01",
          8389 => x"01",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"05",
          8395 => x"05",
          8396 => x"05",
          8397 => x"00",
          8398 => x"01",
          8399 => x"01",
          8400 => x"01",
          8401 => x"01",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"01",
          8428 => x"00",
          8429 => x"01",
          8430 => x"00",
          8431 => x"02",
          8432 => x"00",
          8433 => x"00",
          8434 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
