-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87fa",
          2049 => x"f80d0b0b",
          2050 => x"0b93e904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"cd040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b93b0",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b83bf",
          2210 => x"84738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93b50400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0bac",
          2219 => x"cc2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0bab",
          2227 => x"ab2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"96040b0b",
          2317 => x"0b8ca604",
          2318 => x"0b0b0b8c",
          2319 => x"b6040b0b",
          2320 => x"0b8cc604",
          2321 => x"0b0b0b8c",
          2322 => x"d6040b0b",
          2323 => x"0b8ce604",
          2324 => x"0b0b0b8c",
          2325 => x"f6040b0b",
          2326 => x"0b8d8604",
          2327 => x"0b0b0b8d",
          2328 => x"96040b0b",
          2329 => x"0b8da604",
          2330 => x"0b0b0b8d",
          2331 => x"b6040b0b",
          2332 => x"0b8dc604",
          2333 => x"0b0b0b8d",
          2334 => x"d7040b0b",
          2335 => x"0b8de804",
          2336 => x"0b0b0b8d",
          2337 => x"f9040b0b",
          2338 => x"0b8e8a04",
          2339 => x"0b0b0b8e",
          2340 => x"9b040b0b",
          2341 => x"0b8eac04",
          2342 => x"0b0b0b8e",
          2343 => x"bd040b0b",
          2344 => x"0b8ece04",
          2345 => x"0b0b0b8e",
          2346 => x"df040b0b",
          2347 => x"0b8ef004",
          2348 => x"0b0b0b8f",
          2349 => x"81040b0b",
          2350 => x"0b8f9204",
          2351 => x"0b0b0b8f",
          2352 => x"a3040b0b",
          2353 => x"0b8fb404",
          2354 => x"0b0b0b8f",
          2355 => x"c5040b0b",
          2356 => x"0b8fd604",
          2357 => x"0b0b0b8f",
          2358 => x"e7040b0b",
          2359 => x"0b8ff804",
          2360 => x"0b0b0b90",
          2361 => x"89040b0b",
          2362 => x"0b909a04",
          2363 => x"0b0b0b90",
          2364 => x"ab040b0b",
          2365 => x"0b90bc04",
          2366 => x"0b0b0b90",
          2367 => x"cd040b0b",
          2368 => x"0b90de04",
          2369 => x"0b0b0b90",
          2370 => x"ef040b0b",
          2371 => x"0b918004",
          2372 => x"0b0b0b91",
          2373 => x"91040b0b",
          2374 => x"0b91a204",
          2375 => x"0b0b0b91",
          2376 => x"b3040b0b",
          2377 => x"0b91c404",
          2378 => x"0b0b0b91",
          2379 => x"d5040b0b",
          2380 => x"0b91e604",
          2381 => x"0b0b0b91",
          2382 => x"f7040b0b",
          2383 => x"0b928804",
          2384 => x"0b0b0b92",
          2385 => x"99040b0b",
          2386 => x"0b92aa04",
          2387 => x"0b0b0b92",
          2388 => x"bb040b0b",
          2389 => x"0b92cb04",
          2390 => x"0b0b0b92",
          2391 => x"dc040b0b",
          2392 => x"0b92ed04",
          2393 => x"0b0b0b92",
          2394 => x"fe04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0484bb90",
          2434 => x"0c80d697",
          2435 => x"2d84bb90",
          2436 => x"0880c080",
          2437 => x"900484bb",
          2438 => x"900ca2ee",
          2439 => x"2d84bb90",
          2440 => x"0880c080",
          2441 => x"900484bb",
          2442 => x"900ca0f3",
          2443 => x"2d84bb90",
          2444 => x"0880c080",
          2445 => x"900484bb",
          2446 => x"900ca0e0",
          2447 => x"2d84bb90",
          2448 => x"0880c080",
          2449 => x"900484bb",
          2450 => x"900c94a3",
          2451 => x"2d84bb90",
          2452 => x"0880c080",
          2453 => x"900484bb",
          2454 => x"900ca1f6",
          2455 => x"2d84bb90",
          2456 => x"0880c080",
          2457 => x"900484bb",
          2458 => x"900caf86",
          2459 => x"2d84bb90",
          2460 => x"0880c080",
          2461 => x"900484bb",
          2462 => x"900cad82",
          2463 => x"2d84bb90",
          2464 => x"0880c080",
          2465 => x"900484bb",
          2466 => x"900c9488",
          2467 => x"2d84bb90",
          2468 => x"0880c080",
          2469 => x"900484bb",
          2470 => x"900c95a8",
          2471 => x"2d84bb90",
          2472 => x"0880c080",
          2473 => x"900484bb",
          2474 => x"900c95d1",
          2475 => x"2d84bb90",
          2476 => x"0880c080",
          2477 => x"900484bb",
          2478 => x"900cb18a",
          2479 => x"2d84bb90",
          2480 => x"0880c080",
          2481 => x"900484bb",
          2482 => x"900c80d4",
          2483 => x"fc2d84bb",
          2484 => x"900880c0",
          2485 => x"80900484",
          2486 => x"bb900c80",
          2487 => x"d5e12d84",
          2488 => x"bb900880",
          2489 => x"c0809004",
          2490 => x"84bb900c",
          2491 => x"80d2b82d",
          2492 => x"84bb9008",
          2493 => x"80c08090",
          2494 => x"0484bb90",
          2495 => x"0c80d3eb",
          2496 => x"2d84bb90",
          2497 => x"0880c080",
          2498 => x"900484bb",
          2499 => x"900c82ca",
          2500 => x"f62d84bb",
          2501 => x"900880c0",
          2502 => x"80900484",
          2503 => x"bb900c82",
          2504 => x"e3892d84",
          2505 => x"bb900880",
          2506 => x"c0809004",
          2507 => x"84bb900c",
          2508 => x"82d4c52d",
          2509 => x"84bb9008",
          2510 => x"80c08090",
          2511 => x"0484bb90",
          2512 => x"0c82d9a5",
          2513 => x"2d84bb90",
          2514 => x"0880c080",
          2515 => x"900484bb",
          2516 => x"900c82ed",
          2517 => x"a62d84bb",
          2518 => x"900880c0",
          2519 => x"80900484",
          2520 => x"bb900c82",
          2521 => x"fafc2d84",
          2522 => x"bb900880",
          2523 => x"c0809004",
          2524 => x"84bb900c",
          2525 => x"82deb82d",
          2526 => x"84bb9008",
          2527 => x"80c08090",
          2528 => x"0484bb90",
          2529 => x"0c82f295",
          2530 => x"2d84bb90",
          2531 => x"0880c080",
          2532 => x"900484bb",
          2533 => x"900c82f3",
          2534 => x"e22d84bb",
          2535 => x"900880c0",
          2536 => x"80900484",
          2537 => x"bb900c82",
          2538 => x"f4b72d84",
          2539 => x"bb900880",
          2540 => x"c0809004",
          2541 => x"84bb900c",
          2542 => x"8385b12d",
          2543 => x"84bb9008",
          2544 => x"80c08090",
          2545 => x"0484bb90",
          2546 => x"0c82fff6",
          2547 => x"2d84bb90",
          2548 => x"0880c080",
          2549 => x"900484bb",
          2550 => x"900c838c",
          2551 => x"952d84bb",
          2552 => x"900880c0",
          2553 => x"80900484",
          2554 => x"bb900c82",
          2555 => x"f6942d84",
          2556 => x"bb900880",
          2557 => x"c0809004",
          2558 => x"84bb900c",
          2559 => x"83958c2d",
          2560 => x"84bb9008",
          2561 => x"80c08090",
          2562 => x"0484bb90",
          2563 => x"0c839697",
          2564 => x"2d84bb90",
          2565 => x"0880c080",
          2566 => x"900484bb",
          2567 => x"900c82e5",
          2568 => x"d92d84bb",
          2569 => x"900880c0",
          2570 => x"80900484",
          2571 => x"bb900c82",
          2572 => x"e3f02d84",
          2573 => x"bb900880",
          2574 => x"c0809004",
          2575 => x"84bb900c",
          2576 => x"82e7972d",
          2577 => x"84bb9008",
          2578 => x"80c08090",
          2579 => x"0484bb90",
          2580 => x"0c82f6fe",
          2581 => x"2d84bb90",
          2582 => x"0880c080",
          2583 => x"900484bb",
          2584 => x"900c8397",
          2585 => x"a92d84bb",
          2586 => x"900880c0",
          2587 => x"80900484",
          2588 => x"bb900c83",
          2589 => x"9b862d84",
          2590 => x"bb900880",
          2591 => x"c0809004",
          2592 => x"84bb900c",
          2593 => x"83a1f82d",
          2594 => x"84bb9008",
          2595 => x"80c08090",
          2596 => x"0484bb90",
          2597 => x"0c82c8c7",
          2598 => x"2d84bb90",
          2599 => x"0880c080",
          2600 => x"900484bb",
          2601 => x"900c83a5",
          2602 => x"a12d84bb",
          2603 => x"900880c0",
          2604 => x"80900484",
          2605 => x"bb900c83",
          2606 => x"baa22d84",
          2607 => x"bb900880",
          2608 => x"c0809004",
          2609 => x"84bb900c",
          2610 => x"83b8d42d",
          2611 => x"84bb9008",
          2612 => x"80c08090",
          2613 => x"0484bb90",
          2614 => x"0c81f5ab",
          2615 => x"2d84bb90",
          2616 => x"0880c080",
          2617 => x"900484bb",
          2618 => x"900c81f6",
          2619 => x"aa2d84bb",
          2620 => x"900880c0",
          2621 => x"80900484",
          2622 => x"bb900c81",
          2623 => x"f7a92d84",
          2624 => x"bb900880",
          2625 => x"c0809004",
          2626 => x"84bb900c",
          2627 => x"80d0ba2d",
          2628 => x"84bb9008",
          2629 => x"80c08090",
          2630 => x"0484bb90",
          2631 => x"0c80d28a",
          2632 => x"2d84bb90",
          2633 => x"0880c080",
          2634 => x"900484bb",
          2635 => x"900c80d7",
          2636 => x"b52d84bb",
          2637 => x"900880c0",
          2638 => x"80900484",
          2639 => x"bb900cb1",
          2640 => x"9a2d84bb",
          2641 => x"900880c0",
          2642 => x"80900484",
          2643 => x"bb900c81",
          2644 => x"dcc92d84",
          2645 => x"bb900880",
          2646 => x"c0809004",
          2647 => x"84bb900c",
          2648 => x"81de842d",
          2649 => x"84bb9008",
          2650 => x"80c08090",
          2651 => x"0484bb90",
          2652 => x"0c81f385",
          2653 => x"2d84bb90",
          2654 => x"0880c080",
          2655 => x"900484bb",
          2656 => x"900c81d6",
          2657 => x"d92d84bb",
          2658 => x"900880c0",
          2659 => x"8090043c",
          2660 => x"04101010",
          2661 => x"10101010",
          2662 => x"10101010",
          2663 => x"10101010",
          2664 => x"10101010",
          2665 => x"10101010",
          2666 => x"10101010",
          2667 => x"10101010",
          2668 => x"53510400",
          2669 => x"007381ff",
          2670 => x"06738306",
          2671 => x"09810583",
          2672 => x"05101010",
          2673 => x"2b0772fc",
          2674 => x"060c5151",
          2675 => x"04727280",
          2676 => x"728106ff",
          2677 => x"05097206",
          2678 => x"05711052",
          2679 => x"720a100a",
          2680 => x"5372ed38",
          2681 => x"51515351",
          2682 => x"0484bb84",
          2683 => x"7084e6f0",
          2684 => x"278e3880",
          2685 => x"71708405",
          2686 => x"530c0b0b",
          2687 => x"0b93ec04",
          2688 => x"8c815180",
          2689 => x"ceca0400",
          2690 => x"fc3d0d87",
          2691 => x"3d707084",
          2692 => x"05520856",
          2693 => x"53745284",
          2694 => x"e6e80851",
          2695 => x"81c53f86",
          2696 => x"3d0d04fa",
          2697 => x"3d0d787a",
          2698 => x"7c851133",
          2699 => x"81328106",
          2700 => x"80732507",
          2701 => x"56585557",
          2702 => x"80527272",
          2703 => x"2e098106",
          2704 => x"80d338ff",
          2705 => x"1477748a",
          2706 => x"32703070",
          2707 => x"72079f2a",
          2708 => x"51555556",
          2709 => x"54807425",
          2710 => x"b7387180",
          2711 => x"2eb23875",
          2712 => x"518efa3f",
          2713 => x"84bb8408",
          2714 => x"5384bb84",
          2715 => x"08ff2eae",
          2716 => x"3884bb84",
          2717 => x"08757081",
          2718 => x"055734ff",
          2719 => x"14738a32",
          2720 => x"70307072",
          2721 => x"079f2a51",
          2722 => x"54545473",
          2723 => x"8024cb38",
          2724 => x"80753476",
          2725 => x"527184bb",
          2726 => x"840c883d",
          2727 => x"0d04800b",
          2728 => x"84bb840c",
          2729 => x"883d0d04",
          2730 => x"f53d0d7d",
          2731 => x"54860284",
          2732 => x"05990534",
          2733 => x"7356fe0a",
          2734 => x"588e3d88",
          2735 => x"05537e52",
          2736 => x"8d3de405",
          2737 => x"519d3f73",
          2738 => x"19548074",
          2739 => x"348d3d0d",
          2740 => x"04fd3d0d",
          2741 => x"863d8805",
          2742 => x"53765275",
          2743 => x"51853f85",
          2744 => x"3d0d04f1",
          2745 => x"3d0d6163",
          2746 => x"65425d5d",
          2747 => x"80708c1f",
          2748 => x"0c851e33",
          2749 => x"70812a81",
          2750 => x"32810655",
          2751 => x"555bff54",
          2752 => x"727b2e09",
          2753 => x"810680d2",
          2754 => x"387b3357",
          2755 => x"767b2e80",
          2756 => x"c538811c",
          2757 => x"7b810654",
          2758 => x"5c72802e",
          2759 => x"818138d0",
          2760 => x"175f7e89",
          2761 => x"2681a338",
          2762 => x"76b03270",
          2763 => x"30708025",
          2764 => x"51545578",
          2765 => x"ae387280",
          2766 => x"2ea9387a",
          2767 => x"832a7081",
          2768 => x"32810640",
          2769 => x"547e802e",
          2770 => x"9e387a82",
          2771 => x"80075b7b",
          2772 => x"335776ff",
          2773 => x"bd388c1d",
          2774 => x"08547384",
          2775 => x"bb840c91",
          2776 => x"3d0d047a",
          2777 => x"832a5478",
          2778 => x"10101079",
          2779 => x"10057098",
          2780 => x"2b70982c",
          2781 => x"19708180",
          2782 => x"0a298b0a",
          2783 => x"0570982c",
          2784 => x"525a5b56",
          2785 => x"5f807924",
          2786 => x"81863873",
          2787 => x"81065372",
          2788 => x"ffbd3878",
          2789 => x"7c335858",
          2790 => x"76fef738",
          2791 => x"ffb83976",
          2792 => x"a52e0981",
          2793 => x"06933881",
          2794 => x"73745a5a",
          2795 => x"5b8a7c33",
          2796 => x"585a76fe",
          2797 => x"dd38ff9e",
          2798 => x"397c5276",
          2799 => x"518baf3f",
          2800 => x"7b335776",
          2801 => x"fecc38ff",
          2802 => x"8d397a83",
          2803 => x"2a708106",
          2804 => x"5455788a",
          2805 => x"38817074",
          2806 => x"0640547e",
          2807 => x"9538e017",
          2808 => x"537280d8",
          2809 => x"26973872",
          2810 => x"101083cb",
          2811 => x"94055473",
          2812 => x"080473e0",
          2813 => x"18545980",
          2814 => x"d87327eb",
          2815 => x"387c5276",
          2816 => x"518aeb3f",
          2817 => x"807c3358",
          2818 => x"5b76fe86",
          2819 => x"38fec739",
          2820 => x"80ff59fe",
          2821 => x"f639885a",
          2822 => x"7f608405",
          2823 => x"71087d83",
          2824 => x"ffcf065e",
          2825 => x"58415484",
          2826 => x"bb945e79",
          2827 => x"52755193",
          2828 => x"9a3f84bb",
          2829 => x"840881ff",
          2830 => x"0684bb84",
          2831 => x"0818df05",
          2832 => x"56537289",
          2833 => x"26883884",
          2834 => x"bb8408b0",
          2835 => x"0555747e",
          2836 => x"70810540",
          2837 => x"34795275",
          2838 => x"5190ca3f",
          2839 => x"84bb8408",
          2840 => x"5684bb84",
          2841 => x"08c5387d",
          2842 => x"84bb9431",
          2843 => x"982b7bb2",
          2844 => x"0640567e",
          2845 => x"802e8f38",
          2846 => x"77848080",
          2847 => x"29fc8080",
          2848 => x"0570902c",
          2849 => x"59557a86",
          2850 => x"2a708106",
          2851 => x"555f7380",
          2852 => x"2e9e3877",
          2853 => x"84808029",
          2854 => x"f8808005",
          2855 => x"5379902e",
          2856 => x"8b387784",
          2857 => x"808029fc",
          2858 => x"80800553",
          2859 => x"72902c58",
          2860 => x"7a832a70",
          2861 => x"81065455",
          2862 => x"72802e9e",
          2863 => x"3875982c",
          2864 => x"7081ff06",
          2865 => x"54547873",
          2866 => x"2486cc38",
          2867 => x"7a83fff7",
          2868 => x"0670832a",
          2869 => x"71862a41",
          2870 => x"565b7481",
          2871 => x"06547380",
          2872 => x"2e85f038",
          2873 => x"77793190",
          2874 => x"2b70902c",
          2875 => x"7c838006",
          2876 => x"56595373",
          2877 => x"802e8596",
          2878 => x"387a812a",
          2879 => x"81065473",
          2880 => x"85eb387a",
          2881 => x"842a8106",
          2882 => x"54738698",
          2883 => x"387a852a",
          2884 => x"81065473",
          2885 => x"8697387e",
          2886 => x"81065473",
          2887 => x"858f387a",
          2888 => x"882a8106",
          2889 => x"5f7e802e",
          2890 => x"b2387778",
          2891 => x"84808029",
          2892 => x"fc808005",
          2893 => x"70902c5a",
          2894 => x"40548074",
          2895 => x"259d387c",
          2896 => x"52b05188",
          2897 => x"a93f7778",
          2898 => x"84808029",
          2899 => x"fc808005",
          2900 => x"70902c5a",
          2901 => x"40547380",
          2902 => x"24e53874",
          2903 => x"81065372",
          2904 => x"802eb238",
          2905 => x"78798180",
          2906 => x"0a2981ff",
          2907 => x"0a057098",
          2908 => x"2c5b5555",
          2909 => x"8075259d",
          2910 => x"387c52b0",
          2911 => x"5187ef3f",
          2912 => x"78798180",
          2913 => x"0a2981ff",
          2914 => x"0a057098",
          2915 => x"2c5b5555",
          2916 => x"748024e5",
          2917 => x"387a872a",
          2918 => x"7081065c",
          2919 => x"557a802e",
          2920 => x"81b93876",
          2921 => x"80e32e84",
          2922 => x"d8387680",
          2923 => x"f32e81ca",
          2924 => x"387680d3",
          2925 => x"2e81e238",
          2926 => x"7d84bb94",
          2927 => x"2e96387c",
          2928 => x"52ff1e70",
          2929 => x"33525e87",
          2930 => x"a53f7d84",
          2931 => x"bb942e09",
          2932 => x"8106ec38",
          2933 => x"7481065b",
          2934 => x"7a802efc",
          2935 => x"a7387778",
          2936 => x"84808029",
          2937 => x"fc808005",
          2938 => x"70902c5a",
          2939 => x"40558075",
          2940 => x"25fc9138",
          2941 => x"7c52a051",
          2942 => x"86f43fe2",
          2943 => x"397a9007",
          2944 => x"5b7aa007",
          2945 => x"7c33585b",
          2946 => x"76fa8738",
          2947 => x"fac8397a",
          2948 => x"80c0075b",
          2949 => x"80f85790",
          2950 => x"60618405",
          2951 => x"71087e83",
          2952 => x"ffcf065f",
          2953 => x"5942555a",
          2954 => x"fbfd397f",
          2955 => x"60840577",
          2956 => x"fe800a06",
          2957 => x"83133370",
          2958 => x"982b7207",
          2959 => x"7c848080",
          2960 => x"29fc8080",
          2961 => x"0570902c",
          2962 => x"5e525a56",
          2963 => x"57415f7a",
          2964 => x"872a7081",
          2965 => x"065c557a",
          2966 => x"fec93877",
          2967 => x"78848080",
          2968 => x"29fc8080",
          2969 => x"0570902c",
          2970 => x"5a545f80",
          2971 => x"7f25feb3",
          2972 => x"387c52a0",
          2973 => x"5185f73f",
          2974 => x"e239ff1a",
          2975 => x"7083ffff",
          2976 => x"065b5779",
          2977 => x"83ffff2e",
          2978 => x"feca387c",
          2979 => x"52757081",
          2980 => x"05573351",
          2981 => x"85d83fe2",
          2982 => x"39ff1a70",
          2983 => x"83ffff06",
          2984 => x"5b547983",
          2985 => x"ffff2efe",
          2986 => x"ab387c52",
          2987 => x"75708105",
          2988 => x"57335185",
          2989 => x"b93fe239",
          2990 => x"75fc0a06",
          2991 => x"81fc0a07",
          2992 => x"78848080",
          2993 => x"29fc8080",
          2994 => x"0570902c",
          2995 => x"5a585680",
          2996 => x"e37b872a",
          2997 => x"7081065d",
          2998 => x"56577afd",
          2999 => x"c638fefb",
          3000 => x"397f6084",
          3001 => x"05710870",
          3002 => x"53404156",
          3003 => x"807e2482",
          3004 => x"df387a83",
          3005 => x"ffbf065b",
          3006 => x"84bb945e",
          3007 => x"faad397a",
          3008 => x"84077c33",
          3009 => x"585b76f8",
          3010 => x"8938f8ca",
          3011 => x"397a8807",
          3012 => x"5b807c33",
          3013 => x"585976f7",
          3014 => x"f938f8ba",
          3015 => x"397f6084",
          3016 => x"05710877",
          3017 => x"81065658",
          3018 => x"415f7282",
          3019 => x"8a387551",
          3020 => x"87f63f84",
          3021 => x"bb840883",
          3022 => x"ffff0678",
          3023 => x"7131902b",
          3024 => x"545a7290",
          3025 => x"2c58fe87",
          3026 => x"397a80c0",
          3027 => x"077c3358",
          3028 => x"5b76f7be",
          3029 => x"38f7ff39",
          3030 => x"7f608405",
          3031 => x"71087781",
          3032 => x"065d5841",
          3033 => x"547981cf",
          3034 => x"38755187",
          3035 => x"bb3f84bb",
          3036 => x"840883ff",
          3037 => x"ff067871",
          3038 => x"31902b54",
          3039 => x"5ac4397a",
          3040 => x"8180077c",
          3041 => x"33585b76",
          3042 => x"f78838f7",
          3043 => x"c9397778",
          3044 => x"84808029",
          3045 => x"fc808005",
          3046 => x"70902c5a",
          3047 => x"54548074",
          3048 => x"25fad638",
          3049 => x"7c52a051",
          3050 => x"83c43fe2",
          3051 => x"397c52b0",
          3052 => x"5183bb3f",
          3053 => x"79902e09",
          3054 => x"8106fae3",
          3055 => x"387c5276",
          3056 => x"5183ab3f",
          3057 => x"7a882a81",
          3058 => x"065f7e80",
          3059 => x"2efb8c38",
          3060 => x"fad83975",
          3061 => x"982c7871",
          3062 => x"31902b70",
          3063 => x"902c7d83",
          3064 => x"8006575a",
          3065 => x"515373fa",
          3066 => x"9038ffa2",
          3067 => x"397c52ad",
          3068 => x"5182fb3f",
          3069 => x"7e810654",
          3070 => x"73802efa",
          3071 => x"a238ffad",
          3072 => x"397c5275",
          3073 => x"982a5182",
          3074 => x"e53f7481",
          3075 => x"065b7a80",
          3076 => x"2ef7f138",
          3077 => x"fbc83978",
          3078 => x"7431982b",
          3079 => x"70982c5a",
          3080 => x"53f9b739",
          3081 => x"7c52ab51",
          3082 => x"82c43fc8",
          3083 => x"397c52a0",
          3084 => x"5182bb3f",
          3085 => x"ffbe3978",
          3086 => x"52755188",
          3087 => x"8b3f84bb",
          3088 => x"840883ff",
          3089 => x"ff067871",
          3090 => x"31902b54",
          3091 => x"5afdf339",
          3092 => x"7a82077e",
          3093 => x"307183ff",
          3094 => x"bf065257",
          3095 => x"5bfd9939",
          3096 => x"fe3d0d84",
          3097 => x"e6e40853",
          3098 => x"75527451",
          3099 => x"f3b53f84",
          3100 => x"3d0d04fa",
          3101 => x"3d0d7855",
          3102 => x"800b84e6",
          3103 => x"e8088511",
          3104 => x"3370812a",
          3105 => x"81327081",
          3106 => x"06515658",
          3107 => x"5557ff56",
          3108 => x"72772e09",
          3109 => x"810680d5",
          3110 => x"38747081",
          3111 => x"05563353",
          3112 => x"72772eb0",
          3113 => x"3884e6e8",
          3114 => x"08527251",
          3115 => x"90140853",
          3116 => x"722d84bb",
          3117 => x"8408802e",
          3118 => x"8338ff57",
          3119 => x"74708105",
          3120 => x"56335372",
          3121 => x"802e8838",
          3122 => x"84e6e808",
          3123 => x"54d73984",
          3124 => x"e6e80854",
          3125 => x"84e6e808",
          3126 => x"528a5190",
          3127 => x"14085574",
          3128 => x"2d84bb84",
          3129 => x"08802e83",
          3130 => x"38ff5776",
          3131 => x"567584bb",
          3132 => x"840c883d",
          3133 => x"0d04fa3d",
          3134 => x"0d787a56",
          3135 => x"54800b85",
          3136 => x"16337081",
          3137 => x"2a813270",
          3138 => x"81065155",
          3139 => x"5757ff56",
          3140 => x"72772e09",
          3141 => x"81069238",
          3142 => x"73708105",
          3143 => x"55335372",
          3144 => x"772e0981",
          3145 => x"06983876",
          3146 => x"567584bb",
          3147 => x"840c883d",
          3148 => x"0d047370",
          3149 => x"81055533",
          3150 => x"5372802e",
          3151 => x"ea387452",
          3152 => x"72519015",
          3153 => x"0853722d",
          3154 => x"84bb8408",
          3155 => x"802ee338",
          3156 => x"ff747081",
          3157 => x"05563354",
          3158 => x"5772e338",
          3159 => x"ca39ff3d",
          3160 => x"0d84e6e8",
          3161 => x"08527351",
          3162 => x"853f833d",
          3163 => x"0d04fa3d",
          3164 => x"0d787a85",
          3165 => x"11337081",
          3166 => x"2a813281",
          3167 => x"06565656",
          3168 => x"57ff5672",
          3169 => x"ae387382",
          3170 => x"2a810654",
          3171 => x"73802eac",
          3172 => x"388c1508",
          3173 => x"53728816",
          3174 => x"08259138",
          3175 => x"74085676",
          3176 => x"76347408",
          3177 => x"8105750c",
          3178 => x"8c150853",
          3179 => x"81138c16",
          3180 => x"0c765675",
          3181 => x"84bb840c",
          3182 => x"883d0d04",
          3183 => x"74527681",
          3184 => x"ff065190",
          3185 => x"15085473",
          3186 => x"2dff5684",
          3187 => x"bb8408e3",
          3188 => x"388c1508",
          3189 => x"81058c16",
          3190 => x"0c7656d7",
          3191 => x"39fb3d0d",
          3192 => x"77851133",
          3193 => x"7081ff06",
          3194 => x"70813281",
          3195 => x"06555556",
          3196 => x"56ff5471",
          3197 => x"b3387286",
          3198 => x"2a810652",
          3199 => x"71b33872",
          3200 => x"822a8106",
          3201 => x"5271802e",
          3202 => x"80c33875",
          3203 => x"08703353",
          3204 => x"5371802e",
          3205 => x"80f03881",
          3206 => x"13760c8c",
          3207 => x"16088105",
          3208 => x"8c170c71",
          3209 => x"81ff0654",
          3210 => x"7384bb84",
          3211 => x"0c873d0d",
          3212 => x"0474ffbf",
          3213 => x"06537285",
          3214 => x"17348c16",
          3215 => x"0881058c",
          3216 => x"170c8416",
          3217 => x"3384bb84",
          3218 => x"0c873d0d",
          3219 => x"04755194",
          3220 => x"16085574",
          3221 => x"2d84bb84",
          3222 => x"085284bb",
          3223 => x"84088025",
          3224 => x"ffb93885",
          3225 => x"16337090",
          3226 => x"07545284",
          3227 => x"bb8408ff",
          3228 => x"2e853871",
          3229 => x"a0075372",
          3230 => x"851734ff",
          3231 => x"547384bb",
          3232 => x"840c873d",
          3233 => x"0d0474a0",
          3234 => x"07537285",
          3235 => x"1734ff54",
          3236 => x"ec39fd3d",
          3237 => x"0d757771",
          3238 => x"54545471",
          3239 => x"70810553",
          3240 => x"335170f7",
          3241 => x"38ff1252",
          3242 => x"72708105",
          3243 => x"54335170",
          3244 => x"72708105",
          3245 => x"543470f0",
          3246 => x"387384bb",
          3247 => x"840c853d",
          3248 => x"0d04fc3d",
          3249 => x"0d767971",
          3250 => x"7a555552",
          3251 => x"5470802e",
          3252 => x"9d387372",
          3253 => x"27a13870",
          3254 => x"802e9338",
          3255 => x"71708105",
          3256 => x"53337370",
          3257 => x"81055534",
          3258 => x"ff115170",
          3259 => x"ef387384",
          3260 => x"bb840c86",
          3261 => x"3d0d0470",
          3262 => x"12557375",
          3263 => x"27d93870",
          3264 => x"14755353",
          3265 => x"ff13ff13",
          3266 => x"53537133",
          3267 => x"7334ff11",
          3268 => x"5170802e",
          3269 => x"d938ff13",
          3270 => x"ff135353",
          3271 => x"71337334",
          3272 => x"ff115170",
          3273 => x"df38c739",
          3274 => x"fe3d0d74",
          3275 => x"70535371",
          3276 => x"70810553",
          3277 => x"335170f7",
          3278 => x"38ff1270",
          3279 => x"743184bb",
          3280 => x"840c5184",
          3281 => x"3d0d04fd",
          3282 => x"3d0d7577",
          3283 => x"71545454",
          3284 => x"72708105",
          3285 => x"54335170",
          3286 => x"72708105",
          3287 => x"543470f0",
          3288 => x"387384bb",
          3289 => x"840c853d",
          3290 => x"0d04fd3d",
          3291 => x"0d757871",
          3292 => x"79555552",
          3293 => x"5470802e",
          3294 => x"93387170",
          3295 => x"81055333",
          3296 => x"73708105",
          3297 => x"5534ff11",
          3298 => x"5170ef38",
          3299 => x"7384bb84",
          3300 => x"0c853d0d",
          3301 => x"04fc3d0d",
          3302 => x"76787a55",
          3303 => x"56547280",
          3304 => x"2ea13873",
          3305 => x"33757081",
          3306 => x"05573352",
          3307 => x"5271712e",
          3308 => x"0981069a",
          3309 => x"38811454",
          3310 => x"71802eb7",
          3311 => x"38ff1353",
          3312 => x"72e13880",
          3313 => x"517084bb",
          3314 => x"840c863d",
          3315 => x"0d047280",
          3316 => x"2ef13873",
          3317 => x"3353ff51",
          3318 => x"72802ee9",
          3319 => x"38ff1533",
          3320 => x"52815171",
          3321 => x"802ede38",
          3322 => x"72723184",
          3323 => x"bb840c86",
          3324 => x"3d0d0471",
          3325 => x"84bb840c",
          3326 => x"863d0d04",
          3327 => x"fb3d0d77",
          3328 => x"79537052",
          3329 => x"5680c13f",
          3330 => x"84bb8408",
          3331 => x"84bb8408",
          3332 => x"81055255",
          3333 => x"81b4b23f",
          3334 => x"84bb8408",
          3335 => x"5484bb84",
          3336 => x"08802e9b",
          3337 => x"3884bb84",
          3338 => x"08155480",
          3339 => x"74347453",
          3340 => x"755284bb",
          3341 => x"840851fe",
          3342 => x"b13f84bb",
          3343 => x"84085473",
          3344 => x"84bb840c",
          3345 => x"873d0d04",
          3346 => x"fd3d0d75",
          3347 => x"77717154",
          3348 => x"55535471",
          3349 => x"802e9f38",
          3350 => x"72708105",
          3351 => x"54335170",
          3352 => x"802e8c38",
          3353 => x"ff125271",
          3354 => x"ff2e0981",
          3355 => x"06ea38ff",
          3356 => x"13707531",
          3357 => x"52527084",
          3358 => x"bb840c85",
          3359 => x"3d0d04fd",
          3360 => x"3d0d7577",
          3361 => x"79725553",
          3362 => x"54547080",
          3363 => x"2e8e3872",
          3364 => x"72708105",
          3365 => x"5434ff11",
          3366 => x"5170f438",
          3367 => x"7384bb84",
          3368 => x"0c853d0d",
          3369 => x"04fa3d0d",
          3370 => x"787a5854",
          3371 => x"a0527680",
          3372 => x"2e8b3876",
          3373 => x"5180f53f",
          3374 => x"84bb8408",
          3375 => x"52e01253",
          3376 => x"73802e8d",
          3377 => x"38735180",
          3378 => x"e33f7184",
          3379 => x"bb840831",
          3380 => x"53805272",
          3381 => x"9f2680cb",
          3382 => x"38735272",
          3383 => x"9f2e80c3",
          3384 => x"38811374",
          3385 => x"712aa072",
          3386 => x"3176712b",
          3387 => x"57545455",
          3388 => x"80567476",
          3389 => x"2ea83872",
          3390 => x"10749f2a",
          3391 => x"07741077",
          3392 => x"07787231",
          3393 => x"ff119f2c",
          3394 => x"7081067b",
          3395 => x"72067571",
          3396 => x"31ff1c5c",
          3397 => x"56525255",
          3398 => x"58555374",
          3399 => x"da387310",
          3400 => x"76075271",
          3401 => x"84bb840c",
          3402 => x"883d0d04",
          3403 => x"fc3d0d76",
          3404 => x"70fc8080",
          3405 => x"06703070",
          3406 => x"72078025",
          3407 => x"70842b90",
          3408 => x"71317571",
          3409 => x"2a7083fe",
          3410 => x"80067030",
          3411 => x"70802583",
          3412 => x"2b887131",
          3413 => x"74712a70",
          3414 => x"81f00670",
          3415 => x"30708025",
          3416 => x"822b8471",
          3417 => x"3174712a",
          3418 => x"5553751b",
          3419 => x"05738c06",
          3420 => x"70307080",
          3421 => x"25108271",
          3422 => x"3177712a",
          3423 => x"70812a81",
          3424 => x"32708106",
          3425 => x"70308274",
          3426 => x"31067519",
          3427 => x"0584bb84",
          3428 => x"0c515254",
          3429 => x"55515456",
          3430 => x"5a535555",
          3431 => x"55515656",
          3432 => x"56565158",
          3433 => x"56545286",
          3434 => x"3d0d04fd",
          3435 => x"3d0d7577",
          3436 => x"70547153",
          3437 => x"54548194",
          3438 => x"3f84bb84",
          3439 => x"08732974",
          3440 => x"713184bb",
          3441 => x"840c5385",
          3442 => x"3d0d04fa",
          3443 => x"3d0d787a",
          3444 => x"5854a053",
          3445 => x"76802e8b",
          3446 => x"387651fe",
          3447 => x"cf3f84bb",
          3448 => x"840853e0",
          3449 => x"13527380",
          3450 => x"2e8d3873",
          3451 => x"51febd3f",
          3452 => x"7284bb84",
          3453 => x"08315273",
          3454 => x"53719f26",
          3455 => x"80c53880",
          3456 => x"53719f2e",
          3457 => x"be388112",
          3458 => x"74712aa0",
          3459 => x"72317671",
          3460 => x"2b575454",
          3461 => x"55805674",
          3462 => x"762ea838",
          3463 => x"7210749f",
          3464 => x"2a077410",
          3465 => x"77077872",
          3466 => x"31ff119f",
          3467 => x"2c708106",
          3468 => x"7b720675",
          3469 => x"7131ff1c",
          3470 => x"5c565252",
          3471 => x"55585553",
          3472 => x"74da3872",
          3473 => x"84bb840c",
          3474 => x"883d0d04",
          3475 => x"fa3d0d78",
          3476 => x"9f2c7a9f",
          3477 => x"2c7a9f2c",
          3478 => x"7b327c9f",
          3479 => x"2c7d3273",
          3480 => x"73327174",
          3481 => x"31577275",
          3482 => x"31565956",
          3483 => x"595556fc",
          3484 => x"b43f84bb",
          3485 => x"84087532",
          3486 => x"753184bb",
          3487 => x"840c883d",
          3488 => x"0d04f73d",
          3489 => x"0d7b7d5b",
          3490 => x"5780707b",
          3491 => x"0c770870",
          3492 => x"33565659",
          3493 => x"73a02e09",
          3494 => x"81068f38",
          3495 => x"81157078",
          3496 => x"0c703355",
          3497 => x"5573a02e",
          3498 => x"f33873ad",
          3499 => x"2e80f538",
          3500 => x"73b02e81",
          3501 => x"8338d014",
          3502 => x"58805677",
          3503 => x"892680db",
          3504 => x"388a5880",
          3505 => x"56a07427",
          3506 => x"80c43880",
          3507 => x"e0742789",
          3508 => x"38e01470",
          3509 => x"81ff0655",
          3510 => x"53d01470",
          3511 => x"81ff0651",
          3512 => x"53907327",
          3513 => x"8f38f913",
          3514 => x"7081ff06",
          3515 => x"54548973",
          3516 => x"27818938",
          3517 => x"72782781",
          3518 => x"83387776",
          3519 => x"29138116",
          3520 => x"70790c70",
          3521 => x"33565656",
          3522 => x"73a026ff",
          3523 => x"be387880",
          3524 => x"2e843875",
          3525 => x"3056757a",
          3526 => x"0c815675",
          3527 => x"84bb840c",
          3528 => x"8b3d0d04",
          3529 => x"81701670",
          3530 => x"790c7033",
          3531 => x"56565973",
          3532 => x"b02e0981",
          3533 => x"06feff38",
          3534 => x"81157078",
          3535 => x"0c703355",
          3536 => x"557380e2",
          3537 => x"2ea63890",
          3538 => x"587380f8",
          3539 => x"2ea03881",
          3540 => x"56a07427",
          3541 => x"c638d014",
          3542 => x"53805688",
          3543 => x"58897327",
          3544 => x"fee13875",
          3545 => x"84bb840c",
          3546 => x"8b3d0d04",
          3547 => x"82588115",
          3548 => x"70780c70",
          3549 => x"33555580",
          3550 => x"56feca39",
          3551 => x"800b84bb",
          3552 => x"840c8b3d",
          3553 => x"0d04f73d",
          3554 => x"0d7b7d5b",
          3555 => x"5780707b",
          3556 => x"0c770870",
          3557 => x"33565659",
          3558 => x"73a02e09",
          3559 => x"81068f38",
          3560 => x"81157078",
          3561 => x"0c703355",
          3562 => x"5573a02e",
          3563 => x"f33873ad",
          3564 => x"2e80f538",
          3565 => x"73b02e81",
          3566 => x"8338d014",
          3567 => x"58805677",
          3568 => x"892680db",
          3569 => x"388a5880",
          3570 => x"56a07427",
          3571 => x"80c43880",
          3572 => x"e0742789",
          3573 => x"38e01470",
          3574 => x"81ff0655",
          3575 => x"53d01470",
          3576 => x"81ff0651",
          3577 => x"53907327",
          3578 => x"8f38f913",
          3579 => x"7081ff06",
          3580 => x"54548973",
          3581 => x"27818938",
          3582 => x"72782781",
          3583 => x"83387776",
          3584 => x"29138116",
          3585 => x"70790c70",
          3586 => x"33565656",
          3587 => x"73a026ff",
          3588 => x"be387880",
          3589 => x"2e843875",
          3590 => x"3056757a",
          3591 => x"0c815675",
          3592 => x"84bb840c",
          3593 => x"8b3d0d04",
          3594 => x"81701670",
          3595 => x"790c7033",
          3596 => x"56565973",
          3597 => x"b02e0981",
          3598 => x"06feff38",
          3599 => x"81157078",
          3600 => x"0c703355",
          3601 => x"557380e2",
          3602 => x"2ea63890",
          3603 => x"587380f8",
          3604 => x"2ea03881",
          3605 => x"56a07427",
          3606 => x"c638d014",
          3607 => x"53805688",
          3608 => x"58897327",
          3609 => x"fee13875",
          3610 => x"84bb840c",
          3611 => x"8b3d0d04",
          3612 => x"82588115",
          3613 => x"70780c70",
          3614 => x"33555580",
          3615 => x"56feca39",
          3616 => x"800b84bb",
          3617 => x"840c8b3d",
          3618 => x"0d0480d8",
          3619 => x"aa3f84bb",
          3620 => x"840881ff",
          3621 => x"0684bb84",
          3622 => x"0c04ff3d",
          3623 => x"0d735271",
          3624 => x"93268c38",
          3625 => x"71101083",
          3626 => x"bf940552",
          3627 => x"71080483",
          3628 => x"cfac51ef",
          3629 => x"be3f833d",
          3630 => x"0d0483cf",
          3631 => x"bc51efb3",
          3632 => x"3f833d0d",
          3633 => x"0483cfd4",
          3634 => x"51efa83f",
          3635 => x"833d0d04",
          3636 => x"83cfec51",
          3637 => x"ef9d3f83",
          3638 => x"3d0d0483",
          3639 => x"d08451ef",
          3640 => x"923f833d",
          3641 => x"0d0483d0",
          3642 => x"9451ef87",
          3643 => x"3f833d0d",
          3644 => x"0483d0b4",
          3645 => x"51eefc3f",
          3646 => x"833d0d04",
          3647 => x"83d0c451",
          3648 => x"eef13f83",
          3649 => x"3d0d0483",
          3650 => x"d0ec51ee",
          3651 => x"e63f833d",
          3652 => x"0d0483d1",
          3653 => x"8051eedb",
          3654 => x"3f833d0d",
          3655 => x"0483d19c",
          3656 => x"51eed03f",
          3657 => x"833d0d04",
          3658 => x"83d1b451",
          3659 => x"eec53f83",
          3660 => x"3d0d0483",
          3661 => x"d1cc51ee",
          3662 => x"ba3f833d",
          3663 => x"0d0483d1",
          3664 => x"e451eeaf",
          3665 => x"3f833d0d",
          3666 => x"0483d1f4",
          3667 => x"51eea43f",
          3668 => x"833d0d04",
          3669 => x"83d28851",
          3670 => x"ee993f83",
          3671 => x"3d0d0483",
          3672 => x"d29851ee",
          3673 => x"8e3f833d",
          3674 => x"0d0483d2",
          3675 => x"a851ee83",
          3676 => x"3f833d0d",
          3677 => x"0483d2b8",
          3678 => x"51edf83f",
          3679 => x"833d0d04",
          3680 => x"83d2c851",
          3681 => x"eded3f83",
          3682 => x"3d0d0483",
          3683 => x"d2d451ed",
          3684 => x"e23f833d",
          3685 => x"0d04feec",
          3686 => x"3d0d8197",
          3687 => x"3d080284",
          3688 => x"0584e305",
          3689 => x"335b5880",
          3690 => x"0b81993d",
          3691 => x"08793070",
          3692 => x"7b077325",
          3693 => x"51575759",
          3694 => x"78577587",
          3695 => x"ff268338",
          3696 => x"81577477",
          3697 => x"077081ff",
          3698 => x"06515593",
          3699 => x"577480e2",
          3700 => x"38815377",
          3701 => x"528c3d70",
          3702 => x"52588297",
          3703 => x"993f84bb",
          3704 => x"84085784",
          3705 => x"bb840880",
          3706 => x"2e80d138",
          3707 => x"775182af",
          3708 => x"983f7630",
          3709 => x"70780780",
          3710 => x"257b3070",
          3711 => x"9f2a7206",
          3712 => x"53575758",
          3713 => x"77802eaa",
          3714 => x"3887c098",
          3715 => x"88085574",
          3716 => x"87e72680",
          3717 => x"e3387452",
          3718 => x"7887e829",
          3719 => x"51f5863f",
          3720 => x"84bb8408",
          3721 => x"5483d384",
          3722 => x"53785283",
          3723 => x"d2e051df",
          3724 => x"d73f7684",
          3725 => x"bb840c81",
          3726 => x"963d0d04",
          3727 => x"84bb8408",
          3728 => x"87c09888",
          3729 => x"0c84bb84",
          3730 => x"08598196",
          3731 => x"3dfbd405",
          3732 => x"54848053",
          3733 => x"75527751",
          3734 => x"829fea3f",
          3735 => x"84bb8408",
          3736 => x"5784bb84",
          3737 => x"08ff8538",
          3738 => x"7a557480",
          3739 => x"2efefd38",
          3740 => x"74197517",
          3741 => x"5759d339",
          3742 => x"87e85274",
          3743 => x"51f4a63f",
          3744 => x"84bb8408",
          3745 => x"527851f4",
          3746 => x"9c3f84bb",
          3747 => x"84085483",
          3748 => x"d3845378",
          3749 => x"5283d2e0",
          3750 => x"51deed3f",
          3751 => x"ff9439f8",
          3752 => x"3d0d7c02",
          3753 => x"8405b705",
          3754 => x"335859ff",
          3755 => x"5880537b",
          3756 => x"527a51fd",
          3757 => x"e13f84bb",
          3758 => x"84088b38",
          3759 => x"76802e91",
          3760 => x"3876812e",
          3761 => x"8a387784",
          3762 => x"bb840c8a",
          3763 => x"3d0d0478",
          3764 => x"0484e6e4",
          3765 => x"56615560",
          3766 => x"5484bb84",
          3767 => x"537f527e",
          3768 => x"51782d84",
          3769 => x"bb840884",
          3770 => x"bb840c8a",
          3771 => x"3d0d04f3",
          3772 => x"3d0d7f61",
          3773 => x"63028c05",
          3774 => x"80cf0533",
          3775 => x"73731568",
          3776 => x"415f5c5c",
          3777 => x"5f5d5e78",
          3778 => x"802e8382",
          3779 => x"387a5283",
          3780 => x"d38c51dd",
          3781 => x"f33f83d3",
          3782 => x"9451ddec",
          3783 => x"3f805473",
          3784 => x"7927b238",
          3785 => x"7c902e81",
          3786 => x"ed387ca0",
          3787 => x"2e82a838",
          3788 => x"73185372",
          3789 => x"7a2781a7",
          3790 => x"38723352",
          3791 => x"83d39851",
          3792 => x"ddc63f81",
          3793 => x"1484e6e8",
          3794 => x"085354a0",
          3795 => x"51ec9f3f",
          3796 => x"787426dc",
          3797 => x"3883d3a0",
          3798 => x"51ddad3f",
          3799 => x"80567579",
          3800 => x"2780c038",
          3801 => x"75187033",
          3802 => x"55538055",
          3803 => x"727a2783",
          3804 => x"38815580",
          3805 => x"539f7427",
          3806 => x"83388153",
          3807 => x"74730670",
          3808 => x"81ff0656",
          3809 => x"5774802e",
          3810 => x"883880fe",
          3811 => x"742781ee",
          3812 => x"3884e6e8",
          3813 => x"0852a051",
          3814 => x"ebd43f81",
          3815 => x"16567876",
          3816 => x"26c23883",
          3817 => x"d3a451e9",
          3818 => x"ca3f7818",
          3819 => x"791c5c58",
          3820 => x"80519dc8",
          3821 => x"3f84bb84",
          3822 => x"08982b70",
          3823 => x"982c5854",
          3824 => x"76a02e81",
          3825 => x"ee38769b",
          3826 => x"2e82c338",
          3827 => x"7b1e5776",
          3828 => x"7826feb9",
          3829 => x"38ff0b84",
          3830 => x"bb840c8f",
          3831 => x"3d0d0483",
          3832 => x"d3a851dc",
          3833 => x"a33f8114",
          3834 => x"84e6e808",
          3835 => x"5354a051",
          3836 => x"eafc3f78",
          3837 => x"7426feb8",
          3838 => x"38feda39",
          3839 => x"83d3b851",
          3840 => x"dc863f82",
          3841 => x"1484e6e8",
          3842 => x"085354a0",
          3843 => x"51eadf3f",
          3844 => x"737927fe",
          3845 => x"c0387318",
          3846 => x"53727a27",
          3847 => x"df387222",
          3848 => x"5283d3ac",
          3849 => x"51dbe13f",
          3850 => x"821484e6",
          3851 => x"e8085354",
          3852 => x"a051eaba",
          3853 => x"3f787426",
          3854 => x"dd38fe99",
          3855 => x"3983d3b4",
          3856 => x"51dbc53f",
          3857 => x"841484e6",
          3858 => x"e8085354",
          3859 => x"a051ea9e",
          3860 => x"3f737927",
          3861 => x"fdff3873",
          3862 => x"1853727a",
          3863 => x"27df3872",
          3864 => x"085283d3",
          3865 => x"8c51dba0",
          3866 => x"3f841484",
          3867 => x"e6e80853",
          3868 => x"54a051e9",
          3869 => x"f93f7874",
          3870 => x"26dd38fd",
          3871 => x"d83984e6",
          3872 => x"e8085273",
          3873 => x"51e9e73f",
          3874 => x"811656fe",
          3875 => x"913980d0",
          3876 => x"a63f84bb",
          3877 => x"840881ff",
          3878 => x"06538859",
          3879 => x"72a82efc",
          3880 => x"ec38a059",
          3881 => x"7280d02e",
          3882 => x"098106fc",
          3883 => x"e0389059",
          3884 => x"fcdb3980",
          3885 => x"519bc53f",
          3886 => x"84bb8408",
          3887 => x"982b7098",
          3888 => x"2c70a032",
          3889 => x"7030729b",
          3890 => x"32703070",
          3891 => x"72077375",
          3892 => x"07065155",
          3893 => x"58595758",
          3894 => x"53728025",
          3895 => x"fde83880",
          3896 => x"519b993f",
          3897 => x"84bb8408",
          3898 => x"982b7098",
          3899 => x"2c70a032",
          3900 => x"7030729b",
          3901 => x"32703070",
          3902 => x"72077375",
          3903 => x"07065155",
          3904 => x"58595758",
          3905 => x"53807324",
          3906 => x"ffa938fd",
          3907 => x"b939800b",
          3908 => x"84bb840c",
          3909 => x"8f3d0d04",
          3910 => x"fe3d0d87",
          3911 => x"c0968008",
          3912 => x"53aadd3f",
          3913 => x"81519d8d",
          3914 => x"3f83d4d0",
          3915 => x"519d9e3f",
          3916 => x"80519d81",
          3917 => x"3f72812a",
          3918 => x"70810651",
          3919 => x"527182b7",
          3920 => x"3872822a",
          3921 => x"70810651",
          3922 => x"52718289",
          3923 => x"3872832a",
          3924 => x"70810651",
          3925 => x"527181db",
          3926 => x"3872842a",
          3927 => x"70810651",
          3928 => x"527181ad",
          3929 => x"3872852a",
          3930 => x"70810651",
          3931 => x"527180ff",
          3932 => x"3872862a",
          3933 => x"70810651",
          3934 => x"527180d2",
          3935 => x"3872872a",
          3936 => x"70810651",
          3937 => x"5271a938",
          3938 => x"72882a81",
          3939 => x"06537288",
          3940 => x"38a9f53f",
          3941 => x"843d0d04",
          3942 => x"81519c99",
          3943 => x"3f83d4e8",
          3944 => x"519caa3f",
          3945 => x"80519c8d",
          3946 => x"3fa9dd3f",
          3947 => x"843d0d04",
          3948 => x"81519c81",
          3949 => x"3f83d4fc",
          3950 => x"519c923f",
          3951 => x"80519bf5",
          3952 => x"3f72882a",
          3953 => x"81065372",
          3954 => x"802ec638",
          3955 => x"cb398151",
          3956 => x"9be33f83",
          3957 => x"d590519b",
          3958 => x"f43f8051",
          3959 => x"9bd73f72",
          3960 => x"872a7081",
          3961 => x"06515271",
          3962 => x"802eff9c",
          3963 => x"38c23981",
          3964 => x"519bc23f",
          3965 => x"83d5a451",
          3966 => x"9bd33f80",
          3967 => x"519bb63f",
          3968 => x"72862a70",
          3969 => x"81065152",
          3970 => x"71802efe",
          3971 => x"f038ffbe",
          3972 => x"3981519b",
          3973 => x"a03f83d5",
          3974 => x"b8519bb1",
          3975 => x"3f80519b",
          3976 => x"943f7285",
          3977 => x"2a708106",
          3978 => x"51527180",
          3979 => x"2efec238",
          3980 => x"ffbd3981",
          3981 => x"519afe3f",
          3982 => x"83d5cc51",
          3983 => x"9b8f3f80",
          3984 => x"519af23f",
          3985 => x"72842a70",
          3986 => x"81065152",
          3987 => x"71802efe",
          3988 => x"9438ffbd",
          3989 => x"3981519a",
          3990 => x"dc3f83d5",
          3991 => x"e0519aed",
          3992 => x"3f80519a",
          3993 => x"d03f7283",
          3994 => x"2a708106",
          3995 => x"51527180",
          3996 => x"2efde638",
          3997 => x"ffbd3981",
          3998 => x"519aba3f",
          3999 => x"83d5f051",
          4000 => x"9acb3f80",
          4001 => x"519aae3f",
          4002 => x"72822a70",
          4003 => x"81065152",
          4004 => x"71802efd",
          4005 => x"b838ffbd",
          4006 => x"39ca3d0d",
          4007 => x"80704141",
          4008 => x"ff6184de",
          4009 => x"900c4281",
          4010 => x"52605181",
          4011 => x"b7c93f84",
          4012 => x"bb840881",
          4013 => x"ff069b3d",
          4014 => x"40597861",
          4015 => x"2e84b538",
          4016 => x"83d6c451",
          4017 => x"e3ad3f98",
          4018 => x"3d4383d6",
          4019 => x"fc51d6b8",
          4020 => x"3f7e4880",
          4021 => x"f8538052",
          4022 => x"7e51eba3",
          4023 => x"3f0b0b83",
          4024 => x"eff83370",
          4025 => x"81ff065b",
          4026 => x"5979802e",
          4027 => x"82f13879",
          4028 => x"812e8388",
          4029 => x"387881ff",
          4030 => x"065e7d82",
          4031 => x"2e83c138",
          4032 => x"67705a5a",
          4033 => x"79802e83",
          4034 => x"e0387933",
          4035 => x"5c7ba02e",
          4036 => x"0981068c",
          4037 => x"38811a70",
          4038 => x"335d5a7b",
          4039 => x"a02ef638",
          4040 => x"805c7b9b",
          4041 => x"26be387b",
          4042 => x"902983ef",
          4043 => x"fc057008",
          4044 => x"525be7f4",
          4045 => x"3f84bb84",
          4046 => x"0884bb84",
          4047 => x"08547a53",
          4048 => x"7b08525d",
          4049 => x"e8cf3f84",
          4050 => x"bb84088b",
          4051 => x"38841b33",
          4052 => x"5e7d812e",
          4053 => x"83843881",
          4054 => x"1c7081ff",
          4055 => x"065d5b9b",
          4056 => x"7c27c438",
          4057 => x"9a3d335c",
          4058 => x"7b802efe",
          4059 => x"dd3880f8",
          4060 => x"527e51e9",
          4061 => x"873f84bb",
          4062 => x"84085e84",
          4063 => x"bb840880",
          4064 => x"2e8dce38",
          4065 => x"84bb8408",
          4066 => x"48b83dff",
          4067 => x"80055191",
          4068 => x"a93f84bb",
          4069 => x"84086062",
          4070 => x"065c5c7a",
          4071 => x"802e8184",
          4072 => x"3884bb84",
          4073 => x"0851e780",
          4074 => x"3f84bb84",
          4075 => x"088f2680",
          4076 => x"f338810b",
          4077 => x"a53d5e5b",
          4078 => x"7a822e8d",
          4079 => x"8a387a82",
          4080 => x"248ce738",
          4081 => x"7a812e82",
          4082 => x"e8387b54",
          4083 => x"805383d7",
          4084 => x"80527c51",
          4085 => x"d5d23f83",
          4086 => x"f3c05884",
          4087 => x"bbb4577d",
          4088 => x"56675580",
          4089 => x"5490800a",
          4090 => x"5390800a",
          4091 => x"527c51f5",
          4092 => x"ae3f84bb",
          4093 => x"840884bb",
          4094 => x"84080970",
          4095 => x"30707207",
          4096 => x"8025515b",
          4097 => x"5b42805a",
          4098 => x"7a832683",
          4099 => x"38815a78",
          4100 => x"7a065978",
          4101 => x"802e8d38",
          4102 => x"811b7081",
          4103 => x"ff065c5a",
          4104 => x"7aff9538",
          4105 => x"7f813261",
          4106 => x"8132075d",
          4107 => x"7c81f238",
          4108 => x"61ff2e81",
          4109 => x"ec387d51",
          4110 => x"81969e3f",
          4111 => x"83d6fc51",
          4112 => x"d3c63f7e",
          4113 => x"4880f853",
          4114 => x"80527e51",
          4115 => x"e8b13f0b",
          4116 => x"0b83eff8",
          4117 => x"337081ff",
          4118 => x"065b5979",
          4119 => x"fd913881",
          4120 => x"5383d6a8",
          4121 => x"5284de94",
          4122 => x"51828a8a",
          4123 => x"3f84bb84",
          4124 => x"0880c538",
          4125 => x"810b0b0b",
          4126 => x"83eff834",
          4127 => x"84de9453",
          4128 => x"80f8527e",
          4129 => x"5182f7cc",
          4130 => x"3f84bb84",
          4131 => x"08802ea0",
          4132 => x"3884bb84",
          4133 => x"0851dfdb",
          4134 => x"3f0b0b83",
          4135 => x"eff83370",
          4136 => x"81ff065f",
          4137 => x"597d822e",
          4138 => x"098106fc",
          4139 => x"d3389139",
          4140 => x"84de9451",
          4141 => x"82a1d23f",
          4142 => x"820b0b0b",
          4143 => x"83eff834",
          4144 => x"805583d6",
          4145 => x"b8548053",
          4146 => x"80f8527e",
          4147 => x"51a7d73f",
          4148 => x"67705a5a",
          4149 => x"79fcb338",
          4150 => x"90397c1a",
          4151 => x"630c851b",
          4152 => x"33597881",
          4153 => x"8926fcfc",
          4154 => x"38781010",
          4155 => x"83bfe405",
          4156 => x"5a790804",
          4157 => x"835383d7",
          4158 => x"88527e51",
          4159 => x"e4ec3f60",
          4160 => x"537e5284",
          4161 => x"c8b05182",
          4162 => x"86bd3f84",
          4163 => x"bb840861",
          4164 => x"2e098106",
          4165 => x"fbaa3881",
          4166 => x"709a3d45",
          4167 => x"4141fbaa",
          4168 => x"3983d78c",
          4169 => x"51decc3f",
          4170 => x"7d518194",
          4171 => x"ac3ffe8c",
          4172 => x"3983d79c",
          4173 => x"567b5583",
          4174 => x"d7a05480",
          4175 => x"5383d7a4",
          4176 => x"527c51d2",
          4177 => x"e33ffd8f",
          4178 => x"39818de4",
          4179 => x"3ffafb39",
          4180 => x"9af93ffa",
          4181 => x"f5398152",
          4182 => x"835180c0",
          4183 => x"dc3ffaea",
          4184 => x"39818f8e",
          4185 => x"3ffae339",
          4186 => x"83d7b451",
          4187 => x"de853f80",
          4188 => x"59780483",
          4189 => x"d7c851dd",
          4190 => x"fa3fd0ed",
          4191 => x"3ffacb39",
          4192 => x"b83dff84",
          4193 => x"1153ff80",
          4194 => x"0551ebfa",
          4195 => x"3f84bb84",
          4196 => x"08802efa",
          4197 => x"b5386852",
          4198 => x"83d7e451",
          4199 => x"d0ea3f68",
          4200 => x"5a792d84",
          4201 => x"bb840880",
          4202 => x"2efa9f38",
          4203 => x"84bb8408",
          4204 => x"5283d880",
          4205 => x"51d0d13f",
          4206 => x"fa9039b8",
          4207 => x"3dff8411",
          4208 => x"53ff8005",
          4209 => x"51ebbf3f",
          4210 => x"84bb8408",
          4211 => x"802ef9fa",
          4212 => x"38685283",
          4213 => x"d89c51d0",
          4214 => x"af3f6859",
          4215 => x"7804b83d",
          4216 => x"fef41153",
          4217 => x"ff800551",
          4218 => x"e9983f84",
          4219 => x"bb840880",
          4220 => x"2ef9d738",
          4221 => x"b83dfef0",
          4222 => x"1153ff80",
          4223 => x"0551e982",
          4224 => x"3f84bb84",
          4225 => x"0886d038",
          4226 => x"64597808",
          4227 => x"53785283",
          4228 => x"d8b851cf",
          4229 => x"f33f84e6",
          4230 => x"e4085380",
          4231 => x"f8527e51",
          4232 => x"d0813f7e",
          4233 => x"487e3359",
          4234 => x"78ae2ef9",
          4235 => x"9d38789f",
          4236 => x"2687d338",
          4237 => x"64840570",
          4238 => x"4659cf39",
          4239 => x"b83dfef4",
          4240 => x"1153ff80",
          4241 => x"0551e8ba",
          4242 => x"3f84bb84",
          4243 => x"08802ef8",
          4244 => x"f938b83d",
          4245 => x"fef01153",
          4246 => x"ff800551",
          4247 => x"e8a43f84",
          4248 => x"bb840886",
          4249 => x"b0386459",
          4250 => x"78225378",
          4251 => x"5283d8c8",
          4252 => x"51cf953f",
          4253 => x"84e6e408",
          4254 => x"5380f852",
          4255 => x"7e51cfa3",
          4256 => x"3f7e487e",
          4257 => x"335978ae",
          4258 => x"2ef8bf38",
          4259 => x"789f2687",
          4260 => x"ca386482",
          4261 => x"05704659",
          4262 => x"cf39b83d",
          4263 => x"ff841153",
          4264 => x"ff800551",
          4265 => x"e9e03f84",
          4266 => x"bb840880",
          4267 => x"2ef89b38",
          4268 => x"b83dfefc",
          4269 => x"1153ff80",
          4270 => x"0551e9ca",
          4271 => x"3f84bb84",
          4272 => x"08802ef8",
          4273 => x"8538b83d",
          4274 => x"fef81153",
          4275 => x"ff800551",
          4276 => x"e9b43f84",
          4277 => x"bb840880",
          4278 => x"2ef7ef38",
          4279 => x"83d8d451",
          4280 => x"cea63f68",
          4281 => x"675d5978",
          4282 => x"7c27838d",
          4283 => x"38657033",
          4284 => x"7a335f5c",
          4285 => x"5a7a7d2e",
          4286 => x"95387a55",
          4287 => x"79547833",
          4288 => x"53785283",
          4289 => x"d8e451cd",
          4290 => x"ff3f6666",
          4291 => x"5b5c8119",
          4292 => x"811b4759",
          4293 => x"d239b83d",
          4294 => x"ff841153",
          4295 => x"ff800551",
          4296 => x"e8e43f84",
          4297 => x"bb840880",
          4298 => x"2ef79f38",
          4299 => x"b83dfefc",
          4300 => x"1153ff80",
          4301 => x"0551e8ce",
          4302 => x"3f84bb84",
          4303 => x"08802ef7",
          4304 => x"8938b83d",
          4305 => x"fef81153",
          4306 => x"ff800551",
          4307 => x"e8b83f84",
          4308 => x"bb840880",
          4309 => x"2ef6f338",
          4310 => x"83d98051",
          4311 => x"cdaa3f68",
          4312 => x"5a796727",
          4313 => x"82933865",
          4314 => x"5c797081",
          4315 => x"055b337c",
          4316 => x"34658105",
          4317 => x"46eb39b8",
          4318 => x"3dff8411",
          4319 => x"53ff8005",
          4320 => x"51e8833f",
          4321 => x"84bb8408",
          4322 => x"802ef6be",
          4323 => x"38b83dfe",
          4324 => x"fc1153ff",
          4325 => x"800551e7",
          4326 => x"ed3f84bb",
          4327 => x"8408b138",
          4328 => x"68703354",
          4329 => x"5283d98c",
          4330 => x"51ccdd3f",
          4331 => x"84e6e408",
          4332 => x"5380f852",
          4333 => x"7e51cceb",
          4334 => x"3f7e487e",
          4335 => x"335978ae",
          4336 => x"2ef68738",
          4337 => x"789f2684",
          4338 => x"97386881",
          4339 => x"0549d139",
          4340 => x"68590280",
          4341 => x"db053379",
          4342 => x"34688105",
          4343 => x"49b83dfe",
          4344 => x"fc1153ff",
          4345 => x"800551e7",
          4346 => x"9d3f84bb",
          4347 => x"8408802e",
          4348 => x"f5d83868",
          4349 => x"590280db",
          4350 => x"05337934",
          4351 => x"68810549",
          4352 => x"b83dfefc",
          4353 => x"1153ff80",
          4354 => x"0551e6fa",
          4355 => x"3f84bb84",
          4356 => x"08ffbd38",
          4357 => x"f5b439b8",
          4358 => x"3dff8411",
          4359 => x"53ff8005",
          4360 => x"51e6e33f",
          4361 => x"84bb8408",
          4362 => x"802ef59e",
          4363 => x"38b83dfe",
          4364 => x"fc1153ff",
          4365 => x"800551e6",
          4366 => x"cd3f84bb",
          4367 => x"8408802e",
          4368 => x"f58838b8",
          4369 => x"3dfef811",
          4370 => x"53ff8005",
          4371 => x"51e6b73f",
          4372 => x"84bb8408",
          4373 => x"863884bb",
          4374 => x"84084683",
          4375 => x"d99851cb",
          4376 => x"a73f6867",
          4377 => x"5b59787a",
          4378 => x"278f3865",
          4379 => x"5b7a7970",
          4380 => x"84055b0c",
          4381 => x"797926f5",
          4382 => x"388a51d9",
          4383 => x"e13ff4ca",
          4384 => x"39b83dff",
          4385 => x"80055187",
          4386 => x"b13f84bb",
          4387 => x"8408b93d",
          4388 => x"ff800552",
          4389 => x"5988f33f",
          4390 => x"815384bb",
          4391 => x"84085278",
          4392 => x"51e9f33f",
          4393 => x"84bb8408",
          4394 => x"802ef49e",
          4395 => x"3884bb84",
          4396 => x"0851e7e6",
          4397 => x"3ff49339",
          4398 => x"b83dff84",
          4399 => x"1153ff80",
          4400 => x"0551e5c2",
          4401 => x"3f84bb84",
          4402 => x"08913883",
          4403 => x"f488335a",
          4404 => x"79802e83",
          4405 => x"c03883f3",
          4406 => x"c00849b8",
          4407 => x"3dfefc11",
          4408 => x"53ff8005",
          4409 => x"51e59f3f",
          4410 => x"84bb8408",
          4411 => x"913883f4",
          4412 => x"88335a79",
          4413 => x"802e838a",
          4414 => x"3883f3c4",
          4415 => x"0847b83d",
          4416 => x"fef81153",
          4417 => x"ff800551",
          4418 => x"e4fc3f84",
          4419 => x"bb840880",
          4420 => x"2ea53880",
          4421 => x"665c5c7a",
          4422 => x"882e8338",
          4423 => x"815c7a90",
          4424 => x"32703070",
          4425 => x"72079f2a",
          4426 => x"7e065c5f",
          4427 => x"5d79802e",
          4428 => x"88387aa0",
          4429 => x"2e833888",
          4430 => x"4683d9a8",
          4431 => x"51d6b43f",
          4432 => x"80556854",
          4433 => x"65536652",
          4434 => x"6851eba3",
          4435 => x"3f83d9b4",
          4436 => x"51d6a03f",
          4437 => x"f2f43964",
          4438 => x"64710c59",
          4439 => x"64840545",
          4440 => x"b83dfef0",
          4441 => x"1153ff80",
          4442 => x"0551e296",
          4443 => x"3f84bb84",
          4444 => x"08802ef2",
          4445 => x"d5386464",
          4446 => x"710c5964",
          4447 => x"840545b8",
          4448 => x"3dfef011",
          4449 => x"53ff8005",
          4450 => x"51e1f73f",
          4451 => x"84bb8408",
          4452 => x"c638f2b6",
          4453 => x"39645e02",
          4454 => x"80ce0522",
          4455 => x"7e708205",
          4456 => x"40237d45",
          4457 => x"b83dfef0",
          4458 => x"1153ff80",
          4459 => x"0551e1d2",
          4460 => x"3f84bb84",
          4461 => x"08802ef2",
          4462 => x"9138645e",
          4463 => x"0280ce05",
          4464 => x"227e7082",
          4465 => x"0540237d",
          4466 => x"45b83dfe",
          4467 => x"f01153ff",
          4468 => x"800551e1",
          4469 => x"ad3f84bb",
          4470 => x"8408ffb9",
          4471 => x"38f1eb39",
          4472 => x"b83dfefc",
          4473 => x"1153ff80",
          4474 => x"0551e39a",
          4475 => x"3f84bb84",
          4476 => x"08802e81",
          4477 => x"dc38685c",
          4478 => x"0280db05",
          4479 => x"337c3468",
          4480 => x"810549fb",
          4481 => x"9b39b83d",
          4482 => x"fef01153",
          4483 => x"ff800551",
          4484 => x"e0f03f84",
          4485 => x"bb840880",
          4486 => x"2e819838",
          4487 => x"6464710c",
          4488 => x"5d648405",
          4489 => x"704659f7",
          4490 => x"e1397a83",
          4491 => x"2e098106",
          4492 => x"f398387b",
          4493 => x"5583d7a0",
          4494 => x"54805383",
          4495 => x"d9c0527c",
          4496 => x"51c8e53f",
          4497 => x"f391397b",
          4498 => x"527c51d9",
          4499 => x"fa3ff387",
          4500 => x"3983d9cc",
          4501 => x"51d49c3f",
          4502 => x"f0f039b8",
          4503 => x"3dfef011",
          4504 => x"53ff8005",
          4505 => x"51e09b3f",
          4506 => x"84bb8408",
          4507 => x"802eb838",
          4508 => x"64590280",
          4509 => x"ce052279",
          4510 => x"7082055b",
          4511 => x"237845f7",
          4512 => x"e73983f4",
          4513 => x"89335c7b",
          4514 => x"802e80cf",
          4515 => x"3883f3cc",
          4516 => x"0847fcea",
          4517 => x"3983f489",
          4518 => x"335c7b80",
          4519 => x"2ea13883",
          4520 => x"f3c80849",
          4521 => x"fcb53983",
          4522 => x"d9f851d3",
          4523 => x"c63f6459",
          4524 => x"f7b63983",
          4525 => x"d9f851d3",
          4526 => x"ba3f6459",
          4527 => x"f6cc3983",
          4528 => x"f48a3359",
          4529 => x"78802ea5",
          4530 => x"3883f3d0",
          4531 => x"0849fc8b",
          4532 => x"3983d9f8",
          4533 => x"51d39c3f",
          4534 => x"f9c63983",
          4535 => x"f48a3359",
          4536 => x"78802e9b",
          4537 => x"3883f3d4",
          4538 => x"0847fc92",
          4539 => x"3983f48b",
          4540 => x"335e7d80",
          4541 => x"2e9b3883",
          4542 => x"f3d80849",
          4543 => x"fbdd3983",
          4544 => x"f48b335e",
          4545 => x"7d802e9b",
          4546 => x"3883f3dc",
          4547 => x"0847fbee",
          4548 => x"3983f486",
          4549 => x"335d7c80",
          4550 => x"2e9b3883",
          4551 => x"f3e00849",
          4552 => x"fbb93983",
          4553 => x"f486335d",
          4554 => x"7c802e94",
          4555 => x"3883f3e4",
          4556 => x"0847fbca",
          4557 => x"3983f3f0",
          4558 => x"08fc8005",
          4559 => x"49fb9c39",
          4560 => x"83f3f008",
          4561 => x"880547fb",
          4562 => x"b539f33d",
          4563 => x"0d800b84",
          4564 => x"bbb43487",
          4565 => x"c0948c70",
          4566 => x"08565787",
          4567 => x"84805274",
          4568 => x"51dac23f",
          4569 => x"84bb8408",
          4570 => x"902b7708",
          4571 => x"57558784",
          4572 => x"80527551",
          4573 => x"daaf3f74",
          4574 => x"84bb8408",
          4575 => x"07770c87",
          4576 => x"c0949c70",
          4577 => x"08565787",
          4578 => x"84805274",
          4579 => x"51da963f",
          4580 => x"84bb8408",
          4581 => x"902b7708",
          4582 => x"57558784",
          4583 => x"80527551",
          4584 => x"da833f74",
          4585 => x"84bb8408",
          4586 => x"07770c8c",
          4587 => x"80830b87",
          4588 => x"c094840c",
          4589 => x"8c80830b",
          4590 => x"87c09494",
          4591 => x"0c81beba",
          4592 => x"5c81c9b9",
          4593 => x"5d830284",
          4594 => x"05a10534",
          4595 => x"805e84e6",
          4596 => x"e40b893d",
          4597 => x"7088130c",
          4598 => x"70720c84",
          4599 => x"e6e80c56",
          4600 => x"b8bd3f89",
          4601 => x"9e3f9598",
          4602 => x"3fba9851",
          4603 => x"958d3f83",
          4604 => x"d3c05283",
          4605 => x"d3c451c4",
          4606 => x"8f3f83f3",
          4607 => x"f4702252",
          4608 => x"5594983f",
          4609 => x"83d3cc54",
          4610 => x"83d3d853",
          4611 => x"81153352",
          4612 => x"83d3e051",
          4613 => x"c3f23f8d",
          4614 => x"b23f83d3",
          4615 => x"fc51d0d3",
          4616 => x"3f805283",
          4617 => x"d48051c3",
          4618 => x"df3f9080",
          4619 => x"0a5283d4",
          4620 => x"a851c3d4",
          4621 => x"3fece23f",
          4622 => x"8004fb3d",
          4623 => x"0d777008",
          4624 => x"56568075",
          4625 => x"52537473",
          4626 => x"2e818338",
          4627 => x"74337081",
          4628 => x"ff065252",
          4629 => x"70a02e09",
          4630 => x"81069138",
          4631 => x"81157033",
          4632 => x"7081ff06",
          4633 => x"53535570",
          4634 => x"a02ef138",
          4635 => x"7181ff06",
          4636 => x"5473a22e",
          4637 => x"81823874",
          4638 => x"5272812e",
          4639 => x"80e73880",
          4640 => x"72337081",
          4641 => x"ff065354",
          4642 => x"5470a02e",
          4643 => x"83388154",
          4644 => x"70802e8b",
          4645 => x"3873802e",
          4646 => x"86388112",
          4647 => x"52e13980",
          4648 => x"7381ff06",
          4649 => x"525470a0",
          4650 => x"2e098106",
          4651 => x"83388154",
          4652 => x"70a23270",
          4653 => x"30708025",
          4654 => x"76075252",
          4655 => x"5372802e",
          4656 => x"88388072",
          4657 => x"70810554",
          4658 => x"3471760c",
          4659 => x"74517084",
          4660 => x"bb840c87",
          4661 => x"3d0d0470",
          4662 => x"802ec438",
          4663 => x"73802eff",
          4664 => x"be388112",
          4665 => x"52807233",
          4666 => x"7081ff06",
          4667 => x"53545470",
          4668 => x"a22ee438",
          4669 => x"8154e039",
          4670 => x"81155581",
          4671 => x"75535372",
          4672 => x"812e0981",
          4673 => x"06fef838",
          4674 => x"dc39fc3d",
          4675 => x"0d765372",
          4676 => x"088b3880",
          4677 => x"0b84bb84",
          4678 => x"0c863d0d",
          4679 => x"04863dfc",
          4680 => x"05527251",
          4681 => x"dadc3f84",
          4682 => x"bb840880",
          4683 => x"2ee53874",
          4684 => x"84bb840c",
          4685 => x"863d0d04",
          4686 => x"fc3d0d76",
          4687 => x"821133ff",
          4688 => x"05525381",
          4689 => x"52708b26",
          4690 => x"81983883",
          4691 => x"1333ff05",
          4692 => x"54825273",
          4693 => x"9e26818a",
          4694 => x"38841333",
          4695 => x"51835270",
          4696 => x"972680fe",
          4697 => x"38851333",
          4698 => x"54845273",
          4699 => x"bb2680f2",
          4700 => x"38861333",
          4701 => x"55855274",
          4702 => x"bb2680e6",
          4703 => x"38881322",
          4704 => x"55865274",
          4705 => x"87e72680",
          4706 => x"d9388a13",
          4707 => x"22548752",
          4708 => x"7387e726",
          4709 => x"80cc3881",
          4710 => x"0b87c098",
          4711 => x"9c0c7222",
          4712 => x"87c098bc",
          4713 => x"0c821333",
          4714 => x"87c098b8",
          4715 => x"0c831333",
          4716 => x"87c098b4",
          4717 => x"0c841333",
          4718 => x"87c098b0",
          4719 => x"0c851333",
          4720 => x"87c098ac",
          4721 => x"0c861333",
          4722 => x"87c098a8",
          4723 => x"0c7487c0",
          4724 => x"98a40c73",
          4725 => x"87c098a0",
          4726 => x"0c800b87",
          4727 => x"c0989c0c",
          4728 => x"80527184",
          4729 => x"bb840c86",
          4730 => x"3d0d04f3",
          4731 => x"3d0d7f5b",
          4732 => x"87c0989c",
          4733 => x"5d817d0c",
          4734 => x"87c098bc",
          4735 => x"085e7d7b",
          4736 => x"2387c098",
          4737 => x"b8085c7b",
          4738 => x"821c3487",
          4739 => x"c098b408",
          4740 => x"5a79831c",
          4741 => x"3487c098",
          4742 => x"b0085c7b",
          4743 => x"841c3487",
          4744 => x"c098ac08",
          4745 => x"5a79851c",
          4746 => x"3487c098",
          4747 => x"a8085c7b",
          4748 => x"861c3487",
          4749 => x"c098a408",
          4750 => x"5c7b881c",
          4751 => x"2387c098",
          4752 => x"a0085a79",
          4753 => x"8a1c2380",
          4754 => x"7d0c7983",
          4755 => x"ffff0659",
          4756 => x"7b83ffff",
          4757 => x"0658861b",
          4758 => x"3357851b",
          4759 => x"3356841b",
          4760 => x"3355831b",
          4761 => x"3354821b",
          4762 => x"33537d83",
          4763 => x"ffff0652",
          4764 => x"83d9fc51",
          4765 => x"ffbf913f",
          4766 => x"8f3d0d04",
          4767 => x"fe3d0d02",
          4768 => x"93053353",
          4769 => x"72812ea8",
          4770 => x"38725180",
          4771 => x"e9de3f84",
          4772 => x"bb840898",
          4773 => x"2b70982c",
          4774 => x"515271ff",
          4775 => x"2e098106",
          4776 => x"86387283",
          4777 => x"2ee33871",
          4778 => x"84bb840c",
          4779 => x"843d0d04",
          4780 => x"725180e9",
          4781 => x"b73f84bb",
          4782 => x"8408982b",
          4783 => x"70982c51",
          4784 => x"5271ff2e",
          4785 => x"098106df",
          4786 => x"38725180",
          4787 => x"e99e3f84",
          4788 => x"bb840898",
          4789 => x"2b70982c",
          4790 => x"515271ff",
          4791 => x"2ed238c7",
          4792 => x"39fd3d0d",
          4793 => x"80705452",
          4794 => x"71882b54",
          4795 => x"815180e8",
          4796 => x"fb3f84bb",
          4797 => x"8408982b",
          4798 => x"70982c51",
          4799 => x"5271ff2e",
          4800 => x"eb387372",
          4801 => x"07811454",
          4802 => x"52837325",
          4803 => x"db387184",
          4804 => x"bb840c85",
          4805 => x"3d0d04fc",
          4806 => x"3d0d029b",
          4807 => x"053383f3",
          4808 => x"bc337081",
          4809 => x"ff065355",
          4810 => x"5570802e",
          4811 => x"80f43887",
          4812 => x"c0949408",
          4813 => x"70962a70",
          4814 => x"81065354",
          4815 => x"5270802e",
          4816 => x"8c387191",
          4817 => x"2a708106",
          4818 => x"515170e3",
          4819 => x"38728132",
          4820 => x"81065372",
          4821 => x"802e8a38",
          4822 => x"71932a81",
          4823 => x"065271cf",
          4824 => x"387381ff",
          4825 => x"065187c0",
          4826 => x"94805270",
          4827 => x"802e8638",
          4828 => x"87c09490",
          4829 => x"5274720c",
          4830 => x"7484bb84",
          4831 => x"0c863d0d",
          4832 => x"0471912a",
          4833 => x"70810651",
          4834 => x"51709738",
          4835 => x"72813281",
          4836 => x"06537280",
          4837 => x"2ecb3871",
          4838 => x"932a8106",
          4839 => x"5271802e",
          4840 => x"c03887c0",
          4841 => x"94840870",
          4842 => x"962a7081",
          4843 => x"06535452",
          4844 => x"70cf38d8",
          4845 => x"39ff3d0d",
          4846 => x"028f0533",
          4847 => x"7030709f",
          4848 => x"2a515252",
          4849 => x"7083f3bc",
          4850 => x"34833d0d",
          4851 => x"04fa3d0d",
          4852 => x"78558075",
          4853 => x"33705652",
          4854 => x"5770772e",
          4855 => x"80e73881",
          4856 => x"1583f3bc",
          4857 => x"337081ff",
          4858 => x"06545755",
          4859 => x"71802e80",
          4860 => x"ff3887c0",
          4861 => x"94940870",
          4862 => x"962a7081",
          4863 => x"06535452",
          4864 => x"70802e8c",
          4865 => x"3871912a",
          4866 => x"70810651",
          4867 => x"5170e338",
          4868 => x"72813281",
          4869 => x"06537280",
          4870 => x"2e8a3871",
          4871 => x"932a8106",
          4872 => x"5271cf38",
          4873 => x"7581ff06",
          4874 => x"5187c094",
          4875 => x"80527080",
          4876 => x"2e863887",
          4877 => x"c0949052",
          4878 => x"73720c81",
          4879 => x"17753355",
          4880 => x"5773ff9b",
          4881 => x"387684bb",
          4882 => x"840c883d",
          4883 => x"0d047191",
          4884 => x"2a708106",
          4885 => x"51517098",
          4886 => x"38728132",
          4887 => x"81065372",
          4888 => x"802ec138",
          4889 => x"71932a81",
          4890 => x"06527180",
          4891 => x"2effb538",
          4892 => x"87c09484",
          4893 => x"0870962a",
          4894 => x"70810653",
          4895 => x"545270ce",
          4896 => x"38d739ff",
          4897 => x"3d0d87c0",
          4898 => x"9e800870",
          4899 => x"9c2a8a06",
          4900 => x"52527080",
          4901 => x"2e84ab38",
          4902 => x"87c09ea4",
          4903 => x"0883f3c0",
          4904 => x"0c87c09e",
          4905 => x"a80883f3",
          4906 => x"c40c87c0",
          4907 => x"9e940883",
          4908 => x"f3c80c87",
          4909 => x"c09e9808",
          4910 => x"83f3cc0c",
          4911 => x"87c09e9c",
          4912 => x"0883f3d0",
          4913 => x"0c87c09e",
          4914 => x"a00883f3",
          4915 => x"d40c87c0",
          4916 => x"9eac0883",
          4917 => x"f3d80c87",
          4918 => x"c09eb008",
          4919 => x"83f3dc0c",
          4920 => x"87c09eb4",
          4921 => x"0883f3e0",
          4922 => x"0c87c09e",
          4923 => x"b80883f3",
          4924 => x"e40c87c0",
          4925 => x"9ebc0883",
          4926 => x"f3e80c87",
          4927 => x"c09ec008",
          4928 => x"83f3ec0c",
          4929 => x"87c09ec4",
          4930 => x"0883f3f0",
          4931 => x"0c87c09e",
          4932 => x"80085271",
          4933 => x"83f3f423",
          4934 => x"87c09e84",
          4935 => x"0883f3f8",
          4936 => x"0c87c09e",
          4937 => x"880883f3",
          4938 => x"fc0c87c0",
          4939 => x"9e8c0883",
          4940 => x"f4800c81",
          4941 => x"0b83f484",
          4942 => x"34800b87",
          4943 => x"c09e9008",
          4944 => x"7084800a",
          4945 => x"06515252",
          4946 => x"7082fb38",
          4947 => x"7183f485",
          4948 => x"34800b87",
          4949 => x"c09e9008",
          4950 => x"7088800a",
          4951 => x"06515252",
          4952 => x"70802e83",
          4953 => x"38815271",
          4954 => x"83f48634",
          4955 => x"800b87c0",
          4956 => x"9e900870",
          4957 => x"90800a06",
          4958 => x"51525270",
          4959 => x"802e8338",
          4960 => x"81527183",
          4961 => x"f4873480",
          4962 => x"0b87c09e",
          4963 => x"90087088",
          4964 => x"80800651",
          4965 => x"52527080",
          4966 => x"2e833881",
          4967 => x"527183f4",
          4968 => x"8834800b",
          4969 => x"87c09e90",
          4970 => x"0870a080",
          4971 => x"80065152",
          4972 => x"5270802e",
          4973 => x"83388152",
          4974 => x"7183f489",
          4975 => x"34800b87",
          4976 => x"c09e9008",
          4977 => x"70908080",
          4978 => x"06515252",
          4979 => x"70802e83",
          4980 => x"38815271",
          4981 => x"83f48a34",
          4982 => x"800b87c0",
          4983 => x"9e900870",
          4984 => x"84808006",
          4985 => x"51525270",
          4986 => x"802e8338",
          4987 => x"81527183",
          4988 => x"f48b3480",
          4989 => x"0b87c09e",
          4990 => x"90087082",
          4991 => x"80800651",
          4992 => x"52527080",
          4993 => x"2e833881",
          4994 => x"527183f4",
          4995 => x"8c34800b",
          4996 => x"87c09e90",
          4997 => x"08708180",
          4998 => x"80065152",
          4999 => x"5270802e",
          5000 => x"83388152",
          5001 => x"7183f48d",
          5002 => x"34800b87",
          5003 => x"c09e9008",
          5004 => x"7080c080",
          5005 => x"06515252",
          5006 => x"70802e83",
          5007 => x"38815271",
          5008 => x"83f48e34",
          5009 => x"800b87c0",
          5010 => x"9e900870",
          5011 => x"a0800651",
          5012 => x"52527080",
          5013 => x"2e833881",
          5014 => x"527183f4",
          5015 => x"8f3487c0",
          5016 => x"9e900898",
          5017 => x"8006708a",
          5018 => x"2a535171",
          5019 => x"83f49034",
          5020 => x"800b87c0",
          5021 => x"9e900870",
          5022 => x"84800651",
          5023 => x"52527080",
          5024 => x"2e833881",
          5025 => x"527183f4",
          5026 => x"913487c0",
          5027 => x"9e900883",
          5028 => x"f0067084",
          5029 => x"2a535171",
          5030 => x"83f49234",
          5031 => x"800b87c0",
          5032 => x"9e900870",
          5033 => x"88065152",
          5034 => x"5270802e",
          5035 => x"83388152",
          5036 => x"7183f493",
          5037 => x"3487c09e",
          5038 => x"90088706",
          5039 => x"517083f4",
          5040 => x"9434833d",
          5041 => x"0d048152",
          5042 => x"fd8239fb",
          5043 => x"3d0d83da",
          5044 => x"9451ffb6",
          5045 => x"b33f83f4",
          5046 => x"84335473",
          5047 => x"86a03883",
          5048 => x"daa851c3",
          5049 => x"8e3f83f4",
          5050 => x"86335574",
          5051 => x"85f03883",
          5052 => x"f48b3354",
          5053 => x"7385c738",
          5054 => x"83f48833",
          5055 => x"5675859e",
          5056 => x"3883f489",
          5057 => x"33557484",
          5058 => x"f53883f4",
          5059 => x"8a335473",
          5060 => x"84cc3883",
          5061 => x"f48f3356",
          5062 => x"7584a938",
          5063 => x"83f49333",
          5064 => x"54738486",
          5065 => x"3883f491",
          5066 => x"33557483",
          5067 => x"e33883f4",
          5068 => x"85335675",
          5069 => x"83c53883",
          5070 => x"f4873354",
          5071 => x"7383a738",
          5072 => x"83f48c33",
          5073 => x"55748389",
          5074 => x"3883f48d",
          5075 => x"33567582",
          5076 => x"ea3883f4",
          5077 => x"8e335473",
          5078 => x"81e13883",
          5079 => x"dac051c2",
          5080 => x"923f83f3",
          5081 => x"e8085283",
          5082 => x"dacc51ff",
          5083 => x"b59a3f83",
          5084 => x"f3ec0852",
          5085 => x"83daf451",
          5086 => x"ffb58d3f",
          5087 => x"83f3f008",
          5088 => x"5283db9c",
          5089 => x"51ffb580",
          5090 => x"3f83dbc4",
          5091 => x"51c1e43f",
          5092 => x"83f3f422",
          5093 => x"5283dbcc",
          5094 => x"51ffb4ec",
          5095 => x"3f83f3f8",
          5096 => x"0856bd84",
          5097 => x"c0527551",
          5098 => x"c9fb3f84",
          5099 => x"bb8408bd",
          5100 => x"84c02976",
          5101 => x"71315454",
          5102 => x"84bb8408",
          5103 => x"5283dbf4",
          5104 => x"51ffb4c4",
          5105 => x"3f83f48b",
          5106 => x"335574b9",
          5107 => x"3883f486",
          5108 => x"33557485",
          5109 => x"38873d0d",
          5110 => x"0483f480",
          5111 => x"0856bd84",
          5112 => x"c0527551",
          5113 => x"c9bf3f84",
          5114 => x"bb8408bd",
          5115 => x"84c02976",
          5116 => x"71315454",
          5117 => x"84bb8408",
          5118 => x"5283dca0",
          5119 => x"51ffb488",
          5120 => x"3f873d0d",
          5121 => x"0483f3fc",
          5122 => x"0856bd84",
          5123 => x"c0527551",
          5124 => x"c9933f84",
          5125 => x"bb8408bd",
          5126 => x"84c02976",
          5127 => x"71315454",
          5128 => x"84bb8408",
          5129 => x"5283dccc",
          5130 => x"51ffb3dc",
          5131 => x"3f83f486",
          5132 => x"33557480",
          5133 => x"2eff9e38",
          5134 => x"ff9f3983",
          5135 => x"dcf851c0",
          5136 => x"b23f83da",
          5137 => x"c051c0ab",
          5138 => x"3f83f3e8",
          5139 => x"085283da",
          5140 => x"cc51ffb3",
          5141 => x"b33f83f3",
          5142 => x"ec085283",
          5143 => x"daf451ff",
          5144 => x"b3a63f83",
          5145 => x"f3f00852",
          5146 => x"83db9c51",
          5147 => x"ffb3993f",
          5148 => x"83dbc451",
          5149 => x"ffbffc3f",
          5150 => x"83f3f422",
          5151 => x"5283dbcc",
          5152 => x"51ffb384",
          5153 => x"3f83f3f8",
          5154 => x"0856bd84",
          5155 => x"c0527551",
          5156 => x"c8933f84",
          5157 => x"bb8408bd",
          5158 => x"84c02976",
          5159 => x"71315454",
          5160 => x"84bb8408",
          5161 => x"5283dbf4",
          5162 => x"51ffb2dc",
          5163 => x"3f83f48b",
          5164 => x"33557480",
          5165 => x"2efe9638",
          5166 => x"fecb3983",
          5167 => x"dd8051ff",
          5168 => x"bfb13f83",
          5169 => x"f48e3354",
          5170 => x"73802efd",
          5171 => x"8e38feeb",
          5172 => x"3983dd88",
          5173 => x"51ffbf9b",
          5174 => x"3f83f48d",
          5175 => x"33567580",
          5176 => x"2efcef38",
          5177 => x"d63983dd",
          5178 => x"9451ffbf",
          5179 => x"863f83f4",
          5180 => x"8c335574",
          5181 => x"802efcd1",
          5182 => x"38d73983",
          5183 => x"dda051ff",
          5184 => x"bef13f83",
          5185 => x"f4873354",
          5186 => x"73802efc",
          5187 => x"b338d739",
          5188 => x"83f49233",
          5189 => x"5283ddb4",
          5190 => x"51ffb1ec",
          5191 => x"3f83f485",
          5192 => x"33567580",
          5193 => x"2efc9038",
          5194 => x"d23983f4",
          5195 => x"94335283",
          5196 => x"ddd451ff",
          5197 => x"b1d23f83",
          5198 => x"f4913355",
          5199 => x"74802efb",
          5200 => x"ed38cd39",
          5201 => x"83f49033",
          5202 => x"5283ddf4",
          5203 => x"51ffb1b8",
          5204 => x"3f83f493",
          5205 => x"33547380",
          5206 => x"2efbca38",
          5207 => x"cd3983f3",
          5208 => x"d00883f3",
          5209 => x"d4081154",
          5210 => x"5283de94",
          5211 => x"51ffb198",
          5212 => x"3f83f48f",
          5213 => x"33567580",
          5214 => x"2efba138",
          5215 => x"c73983f3",
          5216 => x"c80883f3",
          5217 => x"cc081154",
          5218 => x"5283deb0",
          5219 => x"51ffb0f8",
          5220 => x"3f83f48a",
          5221 => x"33547380",
          5222 => x"2efaf838",
          5223 => x"c13983f3",
          5224 => x"c00883f3",
          5225 => x"c4081154",
          5226 => x"5283decc",
          5227 => x"51ffb0d8",
          5228 => x"3f83f489",
          5229 => x"33557480",
          5230 => x"2efacf38",
          5231 => x"c13983f3",
          5232 => x"d80883f3",
          5233 => x"dc081154",
          5234 => x"5283dee8",
          5235 => x"51ffb0b8",
          5236 => x"3f83f488",
          5237 => x"33567580",
          5238 => x"2efaa638",
          5239 => x"c13983f3",
          5240 => x"e00883f3",
          5241 => x"e4081154",
          5242 => x"5283df84",
          5243 => x"51ffb098",
          5244 => x"3f83f48b",
          5245 => x"33547380",
          5246 => x"2ef9fd38",
          5247 => x"c13983df",
          5248 => x"a051ffb0",
          5249 => x"833f83da",
          5250 => x"a851ffbc",
          5251 => x"e63f83f4",
          5252 => x"86335574",
          5253 => x"802ef9d7",
          5254 => x"38c439ff",
          5255 => x"3d0d028e",
          5256 => x"05335271",
          5257 => x"85268c38",
          5258 => x"71101083",
          5259 => x"c48c0552",
          5260 => x"71080483",
          5261 => x"dfb451ff",
          5262 => x"afce3f83",
          5263 => x"3d0d0483",
          5264 => x"dfbc51ff",
          5265 => x"afc23f83",
          5266 => x"3d0d0483",
          5267 => x"dfc451ff",
          5268 => x"afb63f83",
          5269 => x"3d0d0483",
          5270 => x"dfcc51ff",
          5271 => x"afaa3f83",
          5272 => x"3d0d0483",
          5273 => x"dfd451ff",
          5274 => x"af9e3f83",
          5275 => x"3d0d0483",
          5276 => x"dfdc51ff",
          5277 => x"af923f83",
          5278 => x"3d0d0471",
          5279 => x"88800c04",
          5280 => x"800b87c0",
          5281 => x"96840c04",
          5282 => x"83f49808",
          5283 => x"87c09684",
          5284 => x"0c04d93d",
          5285 => x"0daa3d08",
          5286 => x"ad3d085a",
          5287 => x"5a817057",
          5288 => x"58805283",
          5289 => x"f4ec0851",
          5290 => x"8287fb3f",
          5291 => x"84bb8408",
          5292 => x"80ed388b",
          5293 => x"3d57ff0b",
          5294 => x"83f4ec08",
          5295 => x"545580f8",
          5296 => x"52765182",
          5297 => x"d38e3f84",
          5298 => x"bb840880",
          5299 => x"2ea43876",
          5300 => x"51c0d53f",
          5301 => x"84bb8408",
          5302 => x"81175755",
          5303 => x"800b84bb",
          5304 => x"8408258e",
          5305 => x"3884bb84",
          5306 => x"08ff0570",
          5307 => x"18555580",
          5308 => x"74347409",
          5309 => x"70307072",
          5310 => x"079f2a51",
          5311 => x"55557876",
          5312 => x"2e853873",
          5313 => x"ffb03883",
          5314 => x"f4ec088c",
          5315 => x"11085351",
          5316 => x"8287933f",
          5317 => x"84bb8408",
          5318 => x"8f387876",
          5319 => x"2e9a3877",
          5320 => x"84bb840c",
          5321 => x"a93d0d04",
          5322 => x"83e3b851",
          5323 => x"ffadd93f",
          5324 => x"78762e09",
          5325 => x"8106e838",
          5326 => x"76527951",
          5327 => x"c0893f79",
          5328 => x"51ffbfe4",
          5329 => x"3fab3d08",
          5330 => x"5684bb84",
          5331 => x"08763476",
          5332 => x"5283e3e4",
          5333 => x"51ffadb0",
          5334 => x"3f800b84",
          5335 => x"bb840ca9",
          5336 => x"3d0d04d8",
          5337 => x"3d0dab3d",
          5338 => x"08ad3d08",
          5339 => x"71725d72",
          5340 => x"3357575a",
          5341 => x"5773a02e",
          5342 => x"81923880",
          5343 => x"0b8d3d59",
          5344 => x"56751010",
          5345 => x"1083f4f8",
          5346 => x"05700852",
          5347 => x"54ffbf98",
          5348 => x"3f84bb84",
          5349 => x"08537952",
          5350 => x"730851ff",
          5351 => x"bff73f84",
          5352 => x"bb840890",
          5353 => x"38841433",
          5354 => x"5473812e",
          5355 => x"81883873",
          5356 => x"822e9938",
          5357 => x"81167081",
          5358 => x"ff065754",
          5359 => x"827627c1",
          5360 => x"38805473",
          5361 => x"84bb840c",
          5362 => x"aa3d0d04",
          5363 => x"811a5aaa",
          5364 => x"3dff8411",
          5365 => x"53ff8005",
          5366 => x"51c7ab3f",
          5367 => x"84bb8408",
          5368 => x"802ed138",
          5369 => x"ff1b5378",
          5370 => x"527651fd",
          5371 => x"a53f84bb",
          5372 => x"840881ff",
          5373 => x"06547380",
          5374 => x"2ec93881",
          5375 => x"167081ff",
          5376 => x"06575482",
          5377 => x"7627fef9",
          5378 => x"38ffb639",
          5379 => x"78337705",
          5380 => x"56767627",
          5381 => x"fee53881",
          5382 => x"15705b70",
          5383 => x"33555573",
          5384 => x"a02e0981",
          5385 => x"06fed438",
          5386 => x"757526eb",
          5387 => x"38800b8d",
          5388 => x"3d5956fe",
          5389 => x"cc397384",
          5390 => x"bb840853",
          5391 => x"83f4ec08",
          5392 => x"52568284",
          5393 => x"e13f84bb",
          5394 => x"840880d0",
          5395 => x"3883f4ec",
          5396 => x"085380f8",
          5397 => x"52775182",
          5398 => x"cffa3f84",
          5399 => x"bb840880",
          5400 => x"2eba3877",
          5401 => x"51ffbdc0",
          5402 => x"3f84bb84",
          5403 => x"0855800b",
          5404 => x"84bb8408",
          5405 => x"259d3884",
          5406 => x"bb8408ff",
          5407 => x"05701958",
          5408 => x"55807734",
          5409 => x"77537552",
          5410 => x"811683e3",
          5411 => x"ac5256ff",
          5412 => x"aaf63f74",
          5413 => x"ff2e0981",
          5414 => x"06ffb238",
          5415 => x"810b84bb",
          5416 => x"840caa3d",
          5417 => x"0d04cd3d",
          5418 => x"0db63d08",
          5419 => x"b83d08ba",
          5420 => x"3d08bc3d",
          5421 => x"08be3d08",
          5422 => x"425b5842",
          5423 => x"5c800bb5",
          5424 => x"3d3483f4",
          5425 => x"f4335d75",
          5426 => x"83f4f034",
          5427 => x"83f4ec08",
          5428 => x"55749e38",
          5429 => x"747681ff",
          5430 => x"06565774",
          5431 => x"802e82ed",
          5432 => x"3877802e",
          5433 => x"91883881",
          5434 => x"7078065a",
          5435 => x"5678908b",
          5436 => x"3877802e",
          5437 => x"90f83894",
          5438 => x"3db53d40",
          5439 => x"408051ea",
          5440 => x"fb3f84bb",
          5441 => x"8408982b",
          5442 => x"70982c5b",
          5443 => x"5779ff2e",
          5444 => x"81d73879",
          5445 => x"81ff0684",
          5446 => x"e2c03370",
          5447 => x"982b7098",
          5448 => x"2c84e2bc",
          5449 => x"3370982b",
          5450 => x"70972c71",
          5451 => x"982c0570",
          5452 => x"101083df",
          5453 => x"e0057008",
          5454 => x"15703351",
          5455 => x"53495d5a",
          5456 => x"525b585c",
          5457 => x"59815774",
          5458 => x"792e80cd",
          5459 => x"38787527",
          5460 => x"81a83875",
          5461 => x"81800a29",
          5462 => x"81ff0a05",
          5463 => x"70982c57",
          5464 => x"42807624",
          5465 => x"81ec3875",
          5466 => x"10167082",
          5467 => x"2b565780",
          5468 => x"0b83dfe4",
          5469 => x"16334357",
          5470 => x"77622591",
          5471 => x"3883dfe0",
          5472 => x"15081870",
          5473 => x"33564278",
          5474 => x"752e81b6",
          5475 => x"3876802e",
          5476 => x"c2387584",
          5477 => x"e2bc3481",
          5478 => x"5776802e",
          5479 => x"81ba3881",
          5480 => x"1b70982b",
          5481 => x"70982c84",
          5482 => x"e2bc3370",
          5483 => x"982b7097",
          5484 => x"2c71982c",
          5485 => x"0570822b",
          5486 => x"83dfe411",
          5487 => x"335f535e",
          5488 => x"5e585d57",
          5489 => x"577a782e",
          5490 => x"81b13876",
          5491 => x"84e2c034",
          5492 => x"8051e9a8",
          5493 => x"3f84bb84",
          5494 => x"08982b70",
          5495 => x"982c5b57",
          5496 => x"79ff2e09",
          5497 => x"8106feab",
          5498 => x"387d802e",
          5499 => x"fe8f387d",
          5500 => x"2dfe8a39",
          5501 => x"815776ff",
          5502 => x"99387581",
          5503 => x"800a2981",
          5504 => x"800a0570",
          5505 => x"982c7081",
          5506 => x"ff065957",
          5507 => x"42769526",
          5508 => x"80c03875",
          5509 => x"10167082",
          5510 => x"2b515580",
          5511 => x"0b83dfe4",
          5512 => x"16334357",
          5513 => x"776225ce",
          5514 => x"3883dfe0",
          5515 => x"15081870",
          5516 => x"33435578",
          5517 => x"622effbc",
          5518 => x"3876802e",
          5519 => x"ffbc38fe",
          5520 => x"d1398157",
          5521 => x"76802efe",
          5522 => x"8a38fec6",
          5523 => x"398157fd",
          5524 => x"90398057",
          5525 => x"76fec838",
          5526 => x"7684e2c0",
          5527 => x"347684e2",
          5528 => x"bc34797f",
          5529 => x"3476600c",
          5530 => x"63557495",
          5531 => x"26fd8e38",
          5532 => x"74101083",
          5533 => x"c4a40557",
          5534 => x"76080483",
          5535 => x"dfe81508",
          5536 => x"600c800b",
          5537 => x"84e2c034",
          5538 => x"800b84e2",
          5539 => x"bc34d939",
          5540 => x"84e2c833",
          5541 => x"5675802e",
          5542 => x"fce33884",
          5543 => x"e6e80852",
          5544 => x"8851ffb5",
          5545 => x"c93f84e2",
          5546 => x"c833ff05",
          5547 => x"5b7a84e2",
          5548 => x"c834fcc9",
          5549 => x"3984e2c8",
          5550 => x"337081ff",
          5551 => x"0684e2c4",
          5552 => x"335a5755",
          5553 => x"757827fc",
          5554 => x"b43884e6",
          5555 => x"e8085281",
          5556 => x"15426184",
          5557 => x"e2c8347b",
          5558 => x"16703352",
          5559 => x"55ffb58e",
          5560 => x"3ffc9a39",
          5561 => x"7c932e90",
          5562 => x"bd387c92",
          5563 => x"2690387c",
          5564 => x"101083f4",
          5565 => x"a0057008",
          5566 => x"5758758f",
          5567 => x"a538800b",
          5568 => x"84e2c434",
          5569 => x"807c3484",
          5570 => x"e2c43384",
          5571 => x"e2c83356",
          5572 => x"5674802e",
          5573 => x"b63884e6",
          5574 => x"e8085288",
          5575 => x"51ffb4ce",
          5576 => x"3f84e6e8",
          5577 => x"0852a051",
          5578 => x"ffb4c33f",
          5579 => x"84e6e808",
          5580 => x"528851ff",
          5581 => x"b4b83f84",
          5582 => x"e2c833ff",
          5583 => x"05597884",
          5584 => x"e2c83478",
          5585 => x"81ff0655",
          5586 => x"74cc387b",
          5587 => x"51ffa5b8",
          5588 => x"3f7584e2",
          5589 => x"c834fba5",
          5590 => x"397c8a38",
          5591 => x"83f4e808",
          5592 => x"56758cf1",
          5593 => x"38ff1d70",
          5594 => x"81ff0658",
          5595 => x"58769226",
          5596 => x"90387c10",
          5597 => x"1083f498",
          5598 => x"05700857",
          5599 => x"55758dbc",
          5600 => x"387c9326",
          5601 => x"faf7387c",
          5602 => x"101083f4",
          5603 => x"9c057008",
          5604 => x"57597580",
          5605 => x"2efae638",
          5606 => x"7551ffb7",
          5607 => x"8b3f84bb",
          5608 => x"840884e2",
          5609 => x"c43484bb",
          5610 => x"840881ff",
          5611 => x"06810553",
          5612 => x"75527b51",
          5613 => x"ffb7b33f",
          5614 => x"84e2c433",
          5615 => x"84e2c833",
          5616 => x"56567480",
          5617 => x"2eff8438",
          5618 => x"84e6e808",
          5619 => x"528851ff",
          5620 => x"b39c3f84",
          5621 => x"e6e80852",
          5622 => x"a051ffb3",
          5623 => x"913f84e6",
          5624 => x"e8085288",
          5625 => x"51ffb386",
          5626 => x"3f84e2c8",
          5627 => x"33ff0555",
          5628 => x"7484e2c8",
          5629 => x"347481ff",
          5630 => x"0655c739",
          5631 => x"84e2c833",
          5632 => x"7081ff06",
          5633 => x"84e2c433",
          5634 => x"5c575575",
          5635 => x"7a27f9ed",
          5636 => x"3884e6e8",
          5637 => x"08528115",
          5638 => x"577684e2",
          5639 => x"c8347b16",
          5640 => x"70335255",
          5641 => x"ffb2c73f",
          5642 => x"84e2c833",
          5643 => x"7081ff06",
          5644 => x"84e2c433",
          5645 => x"5a575575",
          5646 => x"7827f9c1",
          5647 => x"3884e6e8",
          5648 => x"08528115",
          5649 => x"577684e2",
          5650 => x"c8347b16",
          5651 => x"70335255",
          5652 => x"ffb29b3f",
          5653 => x"84e2c833",
          5654 => x"7081ff06",
          5655 => x"84e2c433",
          5656 => x"5a575577",
          5657 => x"7626ffa9",
          5658 => x"38f99239",
          5659 => x"84e2c833",
          5660 => x"84e2c433",
          5661 => x"56567476",
          5662 => x"2ef98238",
          5663 => x"ff155b7a",
          5664 => x"84e2c434",
          5665 => x"75982b70",
          5666 => x"982c7c81",
          5667 => x"ff064457",
          5668 => x"59617624",
          5669 => x"80ef3884",
          5670 => x"e6e80852",
          5671 => x"a051ffb1",
          5672 => x"cd3f84e2",
          5673 => x"c8337098",
          5674 => x"2b70982c",
          5675 => x"84e2c433",
          5676 => x"5a574356",
          5677 => x"747724f8",
          5678 => x"c43884e6",
          5679 => x"e8085288",
          5680 => x"51ffb1aa",
          5681 => x"3f748180",
          5682 => x"0a298180",
          5683 => x"0a057098",
          5684 => x"2c84e2c4",
          5685 => x"335d5659",
          5686 => x"747b24f8",
          5687 => x"a03884e6",
          5688 => x"e8085288",
          5689 => x"51ffb186",
          5690 => x"3f748180",
          5691 => x"0a298180",
          5692 => x"0a057098",
          5693 => x"2c84e2c4",
          5694 => x"335d5659",
          5695 => x"7a7525ff",
          5696 => x"b938f7f9",
          5697 => x"397b1658",
          5698 => x"81183378",
          5699 => x"3484e6e8",
          5700 => x"08527733",
          5701 => x"51ffb0d6",
          5702 => x"3f758180",
          5703 => x"0a298180",
          5704 => x"0a057098",
          5705 => x"2c84e2c4",
          5706 => x"335c5755",
          5707 => x"757a25fe",
          5708 => x"e6387b16",
          5709 => x"58811833",
          5710 => x"783484e6",
          5711 => x"e8085277",
          5712 => x"3351ffb0",
          5713 => x"a93f7581",
          5714 => x"800a2981",
          5715 => x"800a0570",
          5716 => x"982c84e2",
          5717 => x"c4335c57",
          5718 => x"55797624",
          5719 => x"ffa738fe",
          5720 => x"b63984e2",
          5721 => x"c8335574",
          5722 => x"802ef791",
          5723 => x"3884e6e8",
          5724 => x"08528851",
          5725 => x"ffaff73f",
          5726 => x"84e2c833",
          5727 => x"ff055776",
          5728 => x"84e2c834",
          5729 => x"7681ff06",
          5730 => x"55dd3984",
          5731 => x"e2c4337c",
          5732 => x"05418061",
          5733 => x"3484e6e8",
          5734 => x"08528a51",
          5735 => x"ffafcf3f",
          5736 => x"84e2c452",
          5737 => x"7b51f3bb",
          5738 => x"3f84bb84",
          5739 => x"0881ff06",
          5740 => x"58778ada",
          5741 => x"3884e2c4",
          5742 => x"33577680",
          5743 => x"2e80f038",
          5744 => x"83f4f433",
          5745 => x"70101083",
          5746 => x"f49c0570",
          5747 => x"08574156",
          5748 => x"748bc238",
          5749 => x"75822b87",
          5750 => x"fc0683f4",
          5751 => x"9c058118",
          5752 => x"70535759",
          5753 => x"80e8e23f",
          5754 => x"84bb8408",
          5755 => x"790c83f4",
          5756 => x"f4337010",
          5757 => x"1083f49c",
          5758 => x"05700854",
          5759 => x"4383e394",
          5760 => x"525bffa0",
          5761 => x"833f83f4",
          5762 => x"f4337010",
          5763 => x"1083f49c",
          5764 => x"05700857",
          5765 => x"5e5e748b",
          5766 => x"cf3883f4",
          5767 => x"ec085675",
          5768 => x"802e8c38",
          5769 => x"83f4f033",
          5770 => x"5877802e",
          5771 => x"8bde3880",
          5772 => x"0b84e2c8",
          5773 => x"34800b84",
          5774 => x"e2c4347b",
          5775 => x"84bb840c",
          5776 => x"b53d0d04",
          5777 => x"84e2c833",
          5778 => x"5574802e",
          5779 => x"b63884e6",
          5780 => x"e8085288",
          5781 => x"51ffae96",
          5782 => x"3f84e6e8",
          5783 => x"0852a051",
          5784 => x"ffae8b3f",
          5785 => x"84e6e808",
          5786 => x"528851ff",
          5787 => x"ae803f84",
          5788 => x"e2c833ff",
          5789 => x"05426184",
          5790 => x"e2c83461",
          5791 => x"81ff0655",
          5792 => x"74cc3883",
          5793 => x"d38051ff",
          5794 => x"9efe3f80",
          5795 => x"0b84e2c8",
          5796 => x"34800b84",
          5797 => x"e2c434f4",
          5798 => x"e43984e2",
          5799 => x"c8337081",
          5800 => x"ff065c56",
          5801 => x"7a802ef4",
          5802 => x"d43884e2",
          5803 => x"c433ff05",
          5804 => x"5a7984e2",
          5805 => x"c434ff16",
          5806 => x"587784e2",
          5807 => x"c83484e6",
          5808 => x"e8085288",
          5809 => x"51ffada6",
          5810 => x"3f84e2c8",
          5811 => x"3370982b",
          5812 => x"70982c84",
          5813 => x"e2c4335a",
          5814 => x"525a5676",
          5815 => x"762480ef",
          5816 => x"3884e6e8",
          5817 => x"0852a051",
          5818 => x"ffad833f",
          5819 => x"84e2c833",
          5820 => x"70982b70",
          5821 => x"982c84e2",
          5822 => x"c4335c57",
          5823 => x"59567479",
          5824 => x"24f3fa38",
          5825 => x"84e6e808",
          5826 => x"528851ff",
          5827 => x"ace03f74",
          5828 => x"81800a29",
          5829 => x"81800a05",
          5830 => x"70982c84",
          5831 => x"e2c4335c",
          5832 => x"5155747a",
          5833 => x"24f3d638",
          5834 => x"84e6e808",
          5835 => x"528851ff",
          5836 => x"acbc3f74",
          5837 => x"81800a29",
          5838 => x"81800a05",
          5839 => x"70982c84",
          5840 => x"e2c4335c",
          5841 => x"51557975",
          5842 => x"25ffb938",
          5843 => x"f3af397b",
          5844 => x"16578117",
          5845 => x"33773484",
          5846 => x"e6e80852",
          5847 => x"763351ff",
          5848 => x"ac8c3f75",
          5849 => x"81800a29",
          5850 => x"81800a05",
          5851 => x"70982c84",
          5852 => x"e2c43344",
          5853 => x"575b7562",
          5854 => x"25fee638",
          5855 => x"7b165781",
          5856 => x"17337734",
          5857 => x"84e6e808",
          5858 => x"52763351",
          5859 => x"ffabdf3f",
          5860 => x"7581800a",
          5861 => x"2981800a",
          5862 => x"0570982c",
          5863 => x"84e2c433",
          5864 => x"44575b61",
          5865 => x"7624ffa7",
          5866 => x"38feb639",
          5867 => x"837c3480",
          5868 => x"0b811d34",
          5869 => x"84e2c833",
          5870 => x"5574802e",
          5871 => x"b63884e6",
          5872 => x"e8085288",
          5873 => x"51ffaba6",
          5874 => x"3f84e6e8",
          5875 => x"0852a051",
          5876 => x"ffab9b3f",
          5877 => x"84e6e808",
          5878 => x"528851ff",
          5879 => x"ab903f84",
          5880 => x"e2c833ff",
          5881 => x"055d7c84",
          5882 => x"e2c8347c",
          5883 => x"81ff0655",
          5884 => x"74cc3883",
          5885 => x"d38051ff",
          5886 => x"9c8e3f80",
          5887 => x"0b84e2c8",
          5888 => x"34800b84",
          5889 => x"e2c4347b",
          5890 => x"84bb840c",
          5891 => x"b53d0d04",
          5892 => x"84e2c833",
          5893 => x"7081ff06",
          5894 => x"58587661",
          5895 => x"2ef1de38",
          5896 => x"84e2c433",
          5897 => x"55767527",
          5898 => x"ae387498",
          5899 => x"2b70982c",
          5900 => x"57427676",
          5901 => x"24a1387b",
          5902 => x"165b7a33",
          5903 => x"811c3475",
          5904 => x"81800a29",
          5905 => x"81ff0a05",
          5906 => x"70982c84",
          5907 => x"e2c83352",
          5908 => x"57587578",
          5909 => x"25e13881",
          5910 => x"18557484",
          5911 => x"e2c83477",
          5912 => x"81ff067c",
          5913 => x"0559b43d",
          5914 => x"33793484",
          5915 => x"e2c43357",
          5916 => x"7661258b",
          5917 => x"38811756",
          5918 => x"7584e2c4",
          5919 => x"34755784",
          5920 => x"e2c83370",
          5921 => x"81800a29",
          5922 => x"81ff0a05",
          5923 => x"70982c79",
          5924 => x"81ff0645",
          5925 => x"585c5861",
          5926 => x"76248190",
          5927 => x"3877982b",
          5928 => x"70982c78",
          5929 => x"81ff065b",
          5930 => x"575a7579",
          5931 => x"25f0ce38",
          5932 => x"84e6e808",
          5933 => x"528851ff",
          5934 => x"a9b43f75",
          5935 => x"81800a29",
          5936 => x"81800a05",
          5937 => x"70982c84",
          5938 => x"e2c43357",
          5939 => x"57427575",
          5940 => x"25f0aa38",
          5941 => x"84e6e808",
          5942 => x"528851ff",
          5943 => x"a9903f75",
          5944 => x"81800a29",
          5945 => x"81800a05",
          5946 => x"70982c84",
          5947 => x"e2c43357",
          5948 => x"57427476",
          5949 => x"24ffb938",
          5950 => x"f0833984",
          5951 => x"a85180e2",
          5952 => x"c83f84bb",
          5953 => x"840883f4",
          5954 => x"ec0c84bb",
          5955 => x"84085283",
          5956 => x"e2c051ff",
          5957 => x"99f23f83",
          5958 => x"f4ec0855",
          5959 => x"7486a638",
          5960 => x"7583f4f0",
          5961 => x"3477efcf",
          5962 => x"3880c339",
          5963 => x"84e6e808",
          5964 => x"527b1670",
          5965 => x"335258ff",
          5966 => x"a8b43f75",
          5967 => x"81800a29",
          5968 => x"81800a05",
          5969 => x"70982c84",
          5970 => x"e2c43352",
          5971 => x"57577676",
          5972 => x"24da3884",
          5973 => x"e2c83370",
          5974 => x"982b7098",
          5975 => x"2c7981ff",
          5976 => x"065c585b",
          5977 => x"58757925",
          5978 => x"ef9338fe",
          5979 => x"c33983f4",
          5980 => x"ec08802e",
          5981 => x"ef813883",
          5982 => x"f49c5793",
          5983 => x"56760855",
          5984 => x"74bb38ff",
          5985 => x"16841858",
          5986 => x"56758025",
          5987 => x"f038800b",
          5988 => x"83f4f434",
          5989 => x"83f4ec08",
          5990 => x"5574802e",
          5991 => x"eed93874",
          5992 => x"5181e7e5",
          5993 => x"3f83f4ec",
          5994 => x"085180db",
          5995 => x"ac3f800b",
          5996 => x"83f4ec0c",
          5997 => x"943db53d",
          5998 => x"4040eec1",
          5999 => x"39745180",
          6000 => x"db973f80",
          6001 => x"770cff16",
          6002 => x"84185856",
          6003 => x"758025ff",
          6004 => x"ac38ffba",
          6005 => x"397551ff",
          6006 => x"aace3f84",
          6007 => x"bb840884",
          6008 => x"e2c43484",
          6009 => x"bb840881",
          6010 => x"ff068105",
          6011 => x"5375527b",
          6012 => x"51ffaaf6",
          6013 => x"3f930b84",
          6014 => x"e2c43384",
          6015 => x"e2c83357",
          6016 => x"575d7480",
          6017 => x"2ef2c438",
          6018 => x"84e6e808",
          6019 => x"528851ff",
          6020 => x"a6dc3f84",
          6021 => x"e6e80852",
          6022 => x"a051ffa6",
          6023 => x"d13f84e6",
          6024 => x"e8085288",
          6025 => x"51ffa6c6",
          6026 => x"3f84e2c8",
          6027 => x"33ff0559",
          6028 => x"7884e2c8",
          6029 => x"347881ff",
          6030 => x"0655c739",
          6031 => x"7551ffa9",
          6032 => x"e73f84bb",
          6033 => x"840884e2",
          6034 => x"c43484bb",
          6035 => x"840881ff",
          6036 => x"06810553",
          6037 => x"75527b51",
          6038 => x"ffaa8f3f",
          6039 => x"7684e2c4",
          6040 => x"3384e2c8",
          6041 => x"3357575d",
          6042 => x"74802ef1",
          6043 => x"de3884e6",
          6044 => x"e8085288",
          6045 => x"51ffa5f6",
          6046 => x"3f84e6e8",
          6047 => x"0852a051",
          6048 => x"ffa5eb3f",
          6049 => x"84e6e808",
          6050 => x"528851ff",
          6051 => x"a5e03f84",
          6052 => x"e2c833ff",
          6053 => x"05577684",
          6054 => x"e2c83476",
          6055 => x"81ff0655",
          6056 => x"c7397551",
          6057 => x"ffa9813f",
          6058 => x"84bb8408",
          6059 => x"84e2c434",
          6060 => x"84bb8408",
          6061 => x"81ff0681",
          6062 => x"05537552",
          6063 => x"7b51ffa9",
          6064 => x"a93f811d",
          6065 => x"7081ff06",
          6066 => x"84e2c433",
          6067 => x"84e2c833",
          6068 => x"58525e56",
          6069 => x"74802ef0",
          6070 => x"f23884e6",
          6071 => x"e8085288",
          6072 => x"51ffa58a",
          6073 => x"3f84e6e8",
          6074 => x"0852a051",
          6075 => x"ffa4ff3f",
          6076 => x"84e6e808",
          6077 => x"528851ff",
          6078 => x"a4f43f84",
          6079 => x"e2c833ff",
          6080 => x"055b7a84",
          6081 => x"e2c8347a",
          6082 => x"81ff0655",
          6083 => x"c739807c",
          6084 => x"34800b84",
          6085 => x"e2c83480",
          6086 => x"0b84e2c4",
          6087 => x"347b84bb",
          6088 => x"840cb53d",
          6089 => x"0d0483f4",
          6090 => x"9c085675",
          6091 => x"802eefce",
          6092 => x"387551ff",
          6093 => x"a7f23f84",
          6094 => x"bb840884",
          6095 => x"e2c43484",
          6096 => x"bb840881",
          6097 => x"ff068105",
          6098 => x"5375527b",
          6099 => x"51ffa89a",
          6100 => x"3f84e2c4",
          6101 => x"3384e2c8",
          6102 => x"33565674",
          6103 => x"802eefeb",
          6104 => x"3884e6e8",
          6105 => x"08528851",
          6106 => x"ffa4833f",
          6107 => x"84e6e808",
          6108 => x"52a051ff",
          6109 => x"a3f83f84",
          6110 => x"e6e80852",
          6111 => x"8851ffa3",
          6112 => x"ed3f84e2",
          6113 => x"c833ff05",
          6114 => x"597884e2",
          6115 => x"c8347881",
          6116 => x"ff0655c7",
          6117 => x"39745180",
          6118 => x"d7bf3f83",
          6119 => x"f4f43370",
          6120 => x"822b87fc",
          6121 => x"0683f49c",
          6122 => x"05811970",
          6123 => x"54525a56",
          6124 => x"80dd963f",
          6125 => x"84bb8408",
          6126 => x"790c83f4",
          6127 => x"f4337010",
          6128 => x"1083f49c",
          6129 => x"05700854",
          6130 => x"4383e394",
          6131 => x"525bff94",
          6132 => x"b73f83f4",
          6133 => x"f4337010",
          6134 => x"1083f49c",
          6135 => x"05700857",
          6136 => x"5e5e7480",
          6137 => x"2ef4b338",
          6138 => x"75537b52",
          6139 => x"7451ffa6",
          6140 => x"f93f83f4",
          6141 => x"f4338105",
          6142 => x"7081ff06",
          6143 => x"56569375",
          6144 => x"27839f38",
          6145 => x"7783f4f4",
          6146 => x"34f48f39",
          6147 => x"b53dfef8",
          6148 => x"05547653",
          6149 => x"7b527551",
          6150 => x"81d98a3f",
          6151 => x"83f4ec08",
          6152 => x"528a5182",
          6153 => x"b9fc3f83",
          6154 => x"f4ec0851",
          6155 => x"81de893f",
          6156 => x"800b84e2",
          6157 => x"c834800b",
          6158 => x"84e2c434",
          6159 => x"7b84bb84",
          6160 => x"0cb53d0d",
          6161 => x"04935377",
          6162 => x"52745181",
          6163 => x"caa83f84",
          6164 => x"bb840882",
          6165 => x"d53884bb",
          6166 => x"8408973d",
          6167 => x"5c5d83f4",
          6168 => x"ec085380",
          6169 => x"f8527a51",
          6170 => x"82b7e93f",
          6171 => x"84bb8408",
          6172 => x"5a84bb84",
          6173 => x"087b2e09",
          6174 => x"8106e8f5",
          6175 => x"3884bb84",
          6176 => x"0851ffa5",
          6177 => x"a33f84bb",
          6178 => x"84085780",
          6179 => x"0b84bb84",
          6180 => x"082580fb",
          6181 => x"3884bb84",
          6182 => x"08ff0570",
          6183 => x"1b575780",
          6184 => x"76347681",
          6185 => x"ff0683f4",
          6186 => x"f4337010",
          6187 => x"1083f49c",
          6188 => x"05700858",
          6189 => x"41575974",
          6190 => x"818a3875",
          6191 => x"822b87fc",
          6192 => x"0683f49c",
          6193 => x"05811a70",
          6194 => x"53575f80",
          6195 => x"dafb3f84",
          6196 => x"bb84087f",
          6197 => x"0c83f4f4",
          6198 => x"33701010",
          6199 => x"83f49c05",
          6200 => x"70085456",
          6201 => x"83e39452",
          6202 => x"59ff929c",
          6203 => x"3f83f4f4",
          6204 => x"33701010",
          6205 => x"83f49c05",
          6206 => x"70085741",
          6207 => x"4274a038",
          6208 => x"811d7081",
          6209 => x"ff065e56",
          6210 => x"937d2783",
          6211 => x"38805d76",
          6212 => x"ff2e0981",
          6213 => x"06fec738",
          6214 => x"77e7dc38",
          6215 => x"f8d03975",
          6216 => x"53795274",
          6217 => x"51ffa4c2",
          6218 => x"3f83f4f4",
          6219 => x"33810570",
          6220 => x"81ff065b",
          6221 => x"56937a27",
          6222 => x"80e03880",
          6223 => x"0b83f4f4",
          6224 => x"34ffbd39",
          6225 => x"745180d4",
          6226 => x"903f83f4",
          6227 => x"f4337082",
          6228 => x"2b87fc06",
          6229 => x"83f49c05",
          6230 => x"811b7054",
          6231 => x"52405680",
          6232 => x"d9e73f84",
          6233 => x"bb84087f",
          6234 => x"0c83f4f4",
          6235 => x"33701010",
          6236 => x"83f49c05",
          6237 => x"70085456",
          6238 => x"83e39452",
          6239 => x"59ff9188",
          6240 => x"3f83f4f4",
          6241 => x"33701010",
          6242 => x"83f49c05",
          6243 => x"70085741",
          6244 => x"4274802e",
          6245 => x"feea38ff",
          6246 => x"86397583",
          6247 => x"f4f434fe",
          6248 => x"df397583",
          6249 => x"f4f434f0",
          6250 => x"f13983e2",
          6251 => x"d451ff9d",
          6252 => x"c23f77e6",
          6253 => x"c238f7b6",
          6254 => x"39f23d0d",
          6255 => x"0280c305",
          6256 => x"33028405",
          6257 => x"80c70533",
          6258 => x"5b537283",
          6259 => x"26818d38",
          6260 => x"72812e81",
          6261 => x"8b388173",
          6262 => x"25839e38",
          6263 => x"72822e82",
          6264 => x"a83886c7",
          6265 => x"a0805986",
          6266 => x"c7b08070",
          6267 => x"5e578056",
          6268 => x"9fa05879",
          6269 => x"762e9038",
          6270 => x"7583fab4",
          6271 => x"347583fa",
          6272 => x"b5347583",
          6273 => x"fab22383",
          6274 => x"fab03370",
          6275 => x"982b7190",
          6276 => x"2b077188",
          6277 => x"2b077107",
          6278 => x"7a7f5656",
          6279 => x"565b7877",
          6280 => x"27943880",
          6281 => x"74708405",
          6282 => x"560c7473",
          6283 => x"70840555",
          6284 => x"0c767426",
          6285 => x"ee387578",
          6286 => x"27a23883",
          6287 => x"fab03384",
          6288 => x"99d61779",
          6289 => x"78315555",
          6290 => x"55a00be0",
          6291 => x"e0153474",
          6292 => x"74708105",
          6293 => x"5634ff13",
          6294 => x"5372ee38",
          6295 => x"903d0d04",
          6296 => x"86c7a080",
          6297 => x"0b83fab4",
          6298 => x"33701010",
          6299 => x"1183fab5",
          6300 => x"33719029",
          6301 => x"1174055b",
          6302 => x"41584059",
          6303 => x"86c7b080",
          6304 => x"0b84b8f8",
          6305 => x"337081ff",
          6306 => x"0684b8f7",
          6307 => x"337081ff",
          6308 => x"0683fab2",
          6309 => x"227083ff",
          6310 => x"ff067075",
          6311 => x"295d595d",
          6312 => x"585e575b",
          6313 => x"5d737326",
          6314 => x"87387274",
          6315 => x"31752956",
          6316 => x"7981ff06",
          6317 => x"7e81ff06",
          6318 => x"7c81ff06",
          6319 => x"7a83ffff",
          6320 => x"066281ff",
          6321 => x"06707529",
          6322 => x"145d4257",
          6323 => x"575b5c74",
          6324 => x"74268f38",
          6325 => x"83fab433",
          6326 => x"74763105",
          6327 => x"707d291b",
          6328 => x"595f7683",
          6329 => x"065c7b80",
          6330 => x"2efe9c38",
          6331 => x"787d5553",
          6332 => x"727726fe",
          6333 => x"c1388073",
          6334 => x"70810555",
          6335 => x"3483fab0",
          6336 => x"33747081",
          6337 => x"055634e8",
          6338 => x"3986c7a0",
          6339 => x"805986c7",
          6340 => x"b0807084",
          6341 => x"b8f83370",
          6342 => x"81ff0684",
          6343 => x"b8f73370",
          6344 => x"81ff0683",
          6345 => x"fab22270",
          6346 => x"74295d5b",
          6347 => x"5d575e56",
          6348 => x"5e577478",
          6349 => x"2781df38",
          6350 => x"7381ff06",
          6351 => x"7381ff06",
          6352 => x"71712918",
          6353 => x"5a545479",
          6354 => x"802efdbb",
          6355 => x"38800b83",
          6356 => x"fab43480",
          6357 => x"0b83fab5",
          6358 => x"3483fab0",
          6359 => x"3370982b",
          6360 => x"71902b07",
          6361 => x"71882b07",
          6362 => x"71077a7f",
          6363 => x"5656565b",
          6364 => x"767926fd",
          6365 => x"ae38fdbe",
          6366 => x"3972fce6",
          6367 => x"3883fab4",
          6368 => x"337081ff",
          6369 => x"06701010",
          6370 => x"1183fab5",
          6371 => x"33719029",
          6372 => x"1186c7a0",
          6373 => x"80115e57",
          6374 => x"5b56565f",
          6375 => x"86c7b080",
          6376 => x"701484b8",
          6377 => x"f8337081",
          6378 => x"ff0684b8",
          6379 => x"f7337081",
          6380 => x"ff0683fa",
          6381 => x"b2227083",
          6382 => x"ffff067c",
          6383 => x"75296005",
          6384 => x"5e5a415f",
          6385 => x"585f405e",
          6386 => x"57797326",
          6387 => x"8b38727a",
          6388 => x"3115707d",
          6389 => x"29195753",
          6390 => x"7d81ff06",
          6391 => x"7481ff06",
          6392 => x"7171297d",
          6393 => x"83ffff06",
          6394 => x"6281ff06",
          6395 => x"70752958",
          6396 => x"5f5b5c5d",
          6397 => x"557b7826",
          6398 => x"85387775",
          6399 => x"29537973",
          6400 => x"31167983",
          6401 => x"065b5879",
          6402 => x"fde23876",
          6403 => x"83065c7b",
          6404 => x"fdda38fb",
          6405 => x"f2397478",
          6406 => x"317b2956",
          6407 => x"fe9a39fb",
          6408 => x"3d0d878e",
          6409 => x"808c53ff",
          6410 => x"8a733487",
          6411 => x"73348573",
          6412 => x"34817334",
          6413 => x"878e809c",
          6414 => x"5580f475",
          6415 => x"34ffb075",
          6416 => x"34878e80",
          6417 => x"98568076",
          6418 => x"34807634",
          6419 => x"878e8094",
          6420 => x"548a7434",
          6421 => x"807434ff",
          6422 => x"80753481",
          6423 => x"528351fa",
          6424 => x"d83f86c0",
          6425 => x"87e07008",
          6426 => x"545481f8",
          6427 => x"5686c081",
          6428 => x"f8737706",
          6429 => x"84075455",
          6430 => x"72753473",
          6431 => x"087080ff",
          6432 => x"0680c007",
          6433 => x"51537275",
          6434 => x"3486c087",
          6435 => x"cc087077",
          6436 => x"06810751",
          6437 => x"537286c0",
          6438 => x"81f33473",
          6439 => x"0881f706",
          6440 => x"88075372",
          6441 => x"753480d0",
          6442 => x"0b84b8f8",
          6443 => x"34800b84",
          6444 => x"bb840c87",
          6445 => x"3d0d0484",
          6446 => x"b8f83384",
          6447 => x"bb840c04",
          6448 => x"f73d0d02",
          6449 => x"af053302",
          6450 => x"8405b305",
          6451 => x"3384b8f7",
          6452 => x"335b5956",
          6453 => x"81537579",
          6454 => x"2682da38",
          6455 => x"84b8f833",
          6456 => x"83fab533",
          6457 => x"83fab433",
          6458 => x"72712912",
          6459 => x"86c7a080",
          6460 => x"1183fab2",
          6461 => x"225f5157",
          6462 => x"59717c29",
          6463 => x"057083ff",
          6464 => x"ff0683f9",
          6465 => x"8a335357",
          6466 => x"58537281",
          6467 => x"2e83c438",
          6468 => x"83fab222",
          6469 => x"76055574",
          6470 => x"83fab223",
          6471 => x"83fab433",
          6472 => x"76057081",
          6473 => x"ff067a81",
          6474 => x"ff06555b",
          6475 => x"55727a26",
          6476 => x"828c38ff",
          6477 => x"19537283",
          6478 => x"fab43483",
          6479 => x"fab22270",
          6480 => x"83ffff06",
          6481 => x"84b8f633",
          6482 => x"5c555779",
          6483 => x"74268289",
          6484 => x"3884b8f8",
          6485 => x"33767129",
          6486 => x"54588054",
          6487 => x"729f9f26",
          6488 => x"ac388499",
          6489 => x"d6701454",
          6490 => x"55e0e013",
          6491 => x"33e0e016",
          6492 => x"34727081",
          6493 => x"05543375",
          6494 => x"70810557",
          6495 => x"34811454",
          6496 => x"84b8f573",
          6497 => x"27e33873",
          6498 => x"9f9f26a1",
          6499 => x"3883fab0",
          6500 => x"338499d6",
          6501 => x"155455a0",
          6502 => x"0be0e014",
          6503 => x"34747370",
          6504 => x"81055534",
          6505 => x"8114549f",
          6506 => x"9f7427eb",
          6507 => x"3884b8f6",
          6508 => x"33ff0556",
          6509 => x"7583fab2",
          6510 => x"23755778",
          6511 => x"81ff0677",
          6512 => x"83ffff06",
          6513 => x"54547373",
          6514 => x"2681fd38",
          6515 => x"72743181",
          6516 => x"0584b8f8",
          6517 => x"33717129",
          6518 => x"58555775",
          6519 => x"5586c7a0",
          6520 => x"805886c7",
          6521 => x"b0807981",
          6522 => x"ff067581",
          6523 => x"ff067171",
          6524 => x"29195c5c",
          6525 => x"54577579",
          6526 => x"27b93884",
          6527 => x"99d61654",
          6528 => x"e0e01433",
          6529 => x"5384b980",
          6530 => x"13337870",
          6531 => x"81055a34",
          6532 => x"73708105",
          6533 => x"55337770",
          6534 => x"81055934",
          6535 => x"811584b8",
          6536 => x"f83384b8",
          6537 => x"f7337171",
          6538 => x"2919565c",
          6539 => x"5a557275",
          6540 => x"26ce3880",
          6541 => x"537284bb",
          6542 => x"840c8b3d",
          6543 => x"0d047483",
          6544 => x"fab43483",
          6545 => x"fab22270",
          6546 => x"83ffff06",
          6547 => x"84b8f633",
          6548 => x"5c555773",
          6549 => x"7a27fdf9",
          6550 => x"3877802e",
          6551 => x"fedd3878",
          6552 => x"81ff06ff",
          6553 => x"0583fab4",
          6554 => x"33565372",
          6555 => x"752e0981",
          6556 => x"06fec838",
          6557 => x"73763181",
          6558 => x"0584b8f8",
          6559 => x"33717129",
          6560 => x"78722911",
          6561 => x"56525954",
          6562 => x"737327fe",
          6563 => x"ae3883fa",
          6564 => x"b0338499",
          6565 => x"d6157476",
          6566 => x"31555656",
          6567 => x"a00be0e0",
          6568 => x"16347575",
          6569 => x"70810557",
          6570 => x"34ff1353",
          6571 => x"72802efe",
          6572 => x"8a38a00b",
          6573 => x"e0e01634",
          6574 => x"75757081",
          6575 => x"055734ff",
          6576 => x"135372d8",
          6577 => x"38fdf439",
          6578 => x"800b84b8",
          6579 => x"f8335556",
          6580 => x"fe893983",
          6581 => x"fab61533",
          6582 => x"5984b980",
          6583 => x"19337434",
          6584 => x"84b8f733",
          6585 => x"59fca939",
          6586 => x"fc3d0d76",
          6587 => x"0284059f",
          6588 => x"05335351",
          6589 => x"7086269b",
          6590 => x"38701010",
          6591 => x"83c4fc05",
          6592 => x"51700804",
          6593 => x"84b8f833",
          6594 => x"51717127",
          6595 => x"86387183",
          6596 => x"fab53480",
          6597 => x"0b84bb84",
          6598 => x"0c863d0d",
          6599 => x"04800b83",
          6600 => x"fab53483",
          6601 => x"fab43370",
          6602 => x"81ff0654",
          6603 => x"5272802e",
          6604 => x"e238ff12",
          6605 => x"517083fa",
          6606 => x"b434800b",
          6607 => x"84bb840c",
          6608 => x"863d0d04",
          6609 => x"83fab433",
          6610 => x"70733170",
          6611 => x"09709f2c",
          6612 => x"72065455",
          6613 => x"53547083",
          6614 => x"fab434de",
          6615 => x"3983fab4",
          6616 => x"33720584",
          6617 => x"b8f733ff",
          6618 => x"11555651",
          6619 => x"70752583",
          6620 => x"38705372",
          6621 => x"83fab434",
          6622 => x"800b84bb",
          6623 => x"840c863d",
          6624 => x"0d0483fa",
          6625 => x"b5337073",
          6626 => x"31700970",
          6627 => x"9f2c7206",
          6628 => x"54565355",
          6629 => x"7083fab5",
          6630 => x"34800b84",
          6631 => x"bb840c86",
          6632 => x"3d0d0483",
          6633 => x"fab53372",
          6634 => x"0584b8f8",
          6635 => x"33ff1155",
          6636 => x"55517074",
          6637 => x"25833870",
          6638 => x"537283fa",
          6639 => x"b534800b",
          6640 => x"84bb840c",
          6641 => x"863d0d04",
          6642 => x"800b83fa",
          6643 => x"b53483fa",
          6644 => x"b43384b8",
          6645 => x"f733ff05",
          6646 => x"56527175",
          6647 => x"25feb438",
          6648 => x"81125170",
          6649 => x"83fab434",
          6650 => x"fed039ff",
          6651 => x"3d0d028f",
          6652 => x"05335170",
          6653 => x"b126b338",
          6654 => x"70101083",
          6655 => x"c5980551",
          6656 => x"70080483",
          6657 => x"fab03370",
          6658 => x"80f00671",
          6659 => x"842b80f0",
          6660 => x"06707284",
          6661 => x"2a075152",
          6662 => x"53517180",
          6663 => x"f02e0981",
          6664 => x"069c3880",
          6665 => x"f20b83fa",
          6666 => x"b034800b",
          6667 => x"84bb840c",
          6668 => x"833d0d04",
          6669 => x"83fab033",
          6670 => x"819f0690",
          6671 => x"07517083",
          6672 => x"fab03480",
          6673 => x"0b84bb84",
          6674 => x"0c833d0d",
          6675 => x"0483fab0",
          6676 => x"3380f007",
          6677 => x"517083fa",
          6678 => x"b034e839",
          6679 => x"83fab033",
          6680 => x"81fe0686",
          6681 => x"07517083",
          6682 => x"fab034d7",
          6683 => x"3980f10b",
          6684 => x"83fab034",
          6685 => x"800b84bb",
          6686 => x"840c833d",
          6687 => x"0d0483fa",
          6688 => x"b03381fc",
          6689 => x"06840751",
          6690 => x"7083fab0",
          6691 => x"34ffb439",
          6692 => x"83fab033",
          6693 => x"87075170",
          6694 => x"83fab034",
          6695 => x"ffa53983",
          6696 => x"fab03381",
          6697 => x"fd068507",
          6698 => x"517083fa",
          6699 => x"b034ff93",
          6700 => x"3983fab0",
          6701 => x"3381fb06",
          6702 => x"83075170",
          6703 => x"83fab034",
          6704 => x"ff813983",
          6705 => x"fab03381",
          6706 => x"f9068107",
          6707 => x"517083fa",
          6708 => x"b034feef",
          6709 => x"3983fab0",
          6710 => x"3381f806",
          6711 => x"517083fa",
          6712 => x"b034fedf",
          6713 => x"3983fab0",
          6714 => x"3381df06",
          6715 => x"80d00751",
          6716 => x"7083fab0",
          6717 => x"34fecc39",
          6718 => x"83fab033",
          6719 => x"81bf06b0",
          6720 => x"07517083",
          6721 => x"fab034fe",
          6722 => x"ba3983fa",
          6723 => x"b03381ef",
          6724 => x"0680e007",
          6725 => x"517083fa",
          6726 => x"b034fea7",
          6727 => x"3983fab0",
          6728 => x"3381cf06",
          6729 => x"80c00751",
          6730 => x"7083fab0",
          6731 => x"34fe9439",
          6732 => x"83fab033",
          6733 => x"81af06a0",
          6734 => x"07517083",
          6735 => x"fab034fe",
          6736 => x"823983fa",
          6737 => x"b033818f",
          6738 => x"06517083",
          6739 => x"fab034fd",
          6740 => x"f23983fa",
          6741 => x"b03381fa",
          6742 => x"06820751",
          6743 => x"7083fab0",
          6744 => x"34fde039",
          6745 => x"f33d0d02",
          6746 => x"bf053302",
          6747 => x"840580c3",
          6748 => x"053383fa",
          6749 => x"b43383fa",
          6750 => x"b33383fa",
          6751 => x"b53384b8",
          6752 => x"fa334341",
          6753 => x"5f5d5b59",
          6754 => x"78822e82",
          6755 => x"a1387882",
          6756 => x"24a53878",
          6757 => x"812e8182",
          6758 => x"387d84b8",
          6759 => x"fa34800b",
          6760 => x"84b8fc34",
          6761 => x"7a83fab4",
          6762 => x"347b83fa",
          6763 => x"b2237c83",
          6764 => x"fab5348f",
          6765 => x"3d0d0478",
          6766 => x"832e0981",
          6767 => x"06db3880",
          6768 => x"0b84b8fa",
          6769 => x"34810b84",
          6770 => x"b8fc3482",
          6771 => x"0b83fab4",
          6772 => x"34a80b83",
          6773 => x"fab53482",
          6774 => x"0b83fab2",
          6775 => x"23795884",
          6776 => x"b8f83357",
          6777 => x"84b8f733",
          6778 => x"5684b8f6",
          6779 => x"33557b54",
          6780 => x"7c537a52",
          6781 => x"83e4f851",
          6782 => x"ff808d3f",
          6783 => x"7d84b8fa",
          6784 => x"34800b84",
          6785 => x"b8fc347a",
          6786 => x"83fab434",
          6787 => x"7b83fab2",
          6788 => x"237c83fa",
          6789 => x"b5348f3d",
          6790 => x"0d04800b",
          6791 => x"84b8fa34",
          6792 => x"810b84b8",
          6793 => x"fc34800b",
          6794 => x"83fab434",
          6795 => x"a80b83fa",
          6796 => x"b534800b",
          6797 => x"83fab223",
          6798 => x"84ba8733",
          6799 => x"5884ba86",
          6800 => x"335784ba",
          6801 => x"85335679",
          6802 => x"557b547c",
          6803 => x"537a5283",
          6804 => x"e59451fe",
          6805 => x"ffb23f80",
          6806 => x"0b84ba85",
          6807 => x"335a5a79",
          6808 => x"7927a538",
          6809 => x"791084ba",
          6810 => x"d8057022",
          6811 => x"535983e5",
          6812 => x"ac51feff",
          6813 => x"933f811a",
          6814 => x"7081ff06",
          6815 => x"84ba8533",
          6816 => x"525b5978",
          6817 => x"7a26dd38",
          6818 => x"83d3b451",
          6819 => x"fefef93f",
          6820 => x"7d84b8fa",
          6821 => x"34800b84",
          6822 => x"b8fc347a",
          6823 => x"83fab434",
          6824 => x"7b83fab2",
          6825 => x"237c83fa",
          6826 => x"b5348f3d",
          6827 => x"0d04800b",
          6828 => x"84b8fa34",
          6829 => x"810b84b8",
          6830 => x"fc34810b",
          6831 => x"83fab434",
          6832 => x"a80b83fa",
          6833 => x"b534810b",
          6834 => x"83fab223",
          6835 => x"83f8e851",
          6836 => x"ff90d53f",
          6837 => x"84bb8408",
          6838 => x"5283e5b0",
          6839 => x"51fefea8",
          6840 => x"3f805983",
          6841 => x"f8e851ff",
          6842 => x"90be3f78",
          6843 => x"84bb8408",
          6844 => x"27fda638",
          6845 => x"83f8e819",
          6846 => x"335283e5",
          6847 => x"b851fefe",
          6848 => x"873f8119",
          6849 => x"7081ff06",
          6850 => x"5a5ad839",
          6851 => x"f93d0d7a",
          6852 => x"028405a7",
          6853 => x"053384b8",
          6854 => x"f83383fa",
          6855 => x"b53383fa",
          6856 => x"b4337271",
          6857 => x"291286c7",
          6858 => x"a0801183",
          6859 => x"fab22253",
          6860 => x"51595c71",
          6861 => x"7c290570",
          6862 => x"83ffff06",
          6863 => x"83f98a33",
          6864 => x"52595155",
          6865 => x"57577281",
          6866 => x"2e81e938",
          6867 => x"75892e81",
          6868 => x"f9387589",
          6869 => x"2481b938",
          6870 => x"75812e83",
          6871 => x"85387588",
          6872 => x"2e82d538",
          6873 => x"84b8f833",
          6874 => x"83fab433",
          6875 => x"83fab533",
          6876 => x"72722905",
          6877 => x"55565484",
          6878 => x"b9801633",
          6879 => x"86c7a080",
          6880 => x"143484b8",
          6881 => x"f83383fa",
          6882 => x"b53383fa",
          6883 => x"b2227271",
          6884 => x"29125a5a",
          6885 => x"56537583",
          6886 => x"fab61834",
          6887 => x"83fab433",
          6888 => x"73712916",
          6889 => x"585483fa",
          6890 => x"b03386c7",
          6891 => x"b0801834",
          6892 => x"84b8f833",
          6893 => x"7081ff06",
          6894 => x"83fab222",
          6895 => x"83fab533",
          6896 => x"72722911",
          6897 => x"575b5755",
          6898 => x"5783fab0",
          6899 => x"338499d6",
          6900 => x"14348118",
          6901 => x"7081ff06",
          6902 => x"59557378",
          6903 => x"26819938",
          6904 => x"84b8f933",
          6905 => x"587781ea",
          6906 => x"38ff1753",
          6907 => x"7283fab5",
          6908 => x"3484b8fb",
          6909 => x"33537280",
          6910 => x"2e8c3884",
          6911 => x"b8fc3357",
          6912 => x"76802e80",
          6913 => x"fb38800b",
          6914 => x"84bb840c",
          6915 => x"893d0d04",
          6916 => x"758d2e97",
          6917 => x"38758d24",
          6918 => x"80f73875",
          6919 => x"8a2e0981",
          6920 => x"06fec138",
          6921 => x"81528151",
          6922 => x"f1963f80",
          6923 => x"0b83fab5",
          6924 => x"34ffbe39",
          6925 => x"83fab615",
          6926 => x"335384b9",
          6927 => x"80133374",
          6928 => x"3475892e",
          6929 => x"098106fe",
          6930 => x"89388053",
          6931 => x"7652a051",
          6932 => x"fdba3f81",
          6933 => x"137081ff",
          6934 => x"06545472",
          6935 => x"8326ff91",
          6936 => x"387652a0",
          6937 => x"51fda53f",
          6938 => x"81137081",
          6939 => x"ff065454",
          6940 => x"837327d8",
          6941 => x"38fefa39",
          6942 => x"7483fab5",
          6943 => x"34fef239",
          6944 => x"75528351",
          6945 => x"f9de3f80",
          6946 => x"0b84bb84",
          6947 => x"0c893d0d",
          6948 => x"047580ff",
          6949 => x"2e098106",
          6950 => x"fdca3883",
          6951 => x"fab53370",
          6952 => x"81ff0655",
          6953 => x"ff055373",
          6954 => x"83387353",
          6955 => x"7283fab5",
          6956 => x"347652a0",
          6957 => x"51fcd53f",
          6958 => x"83fab533",
          6959 => x"7081ff06",
          6960 => x"55ff0553",
          6961 => x"73fea538",
          6962 => x"73537283",
          6963 => x"fab534fe",
          6964 => x"a039800b",
          6965 => x"83fab534",
          6966 => x"81528151",
          6967 => x"efe23ffe",
          6968 => x"90398052",
          6969 => x"7551efd8",
          6970 => x"3ffe8639",
          6971 => x"e63d0d02",
          6972 => x"80f30533",
          6973 => x"84ba8008",
          6974 => x"57597581",
          6975 => x"2e81b838",
          6976 => x"75822e83",
          6977 => x"8238788a",
          6978 => x"2e84b538",
          6979 => x"788a2482",
          6980 => x"d1387888",
          6981 => x"2e84b938",
          6982 => x"78892e88",
          6983 => x"8f3884b8",
          6984 => x"f83383fa",
          6985 => x"b43383fa",
          6986 => x"b5337272",
          6987 => x"2905585e",
          6988 => x"5c84b980",
          6989 => x"193386c7",
          6990 => x"a0801734",
          6991 => x"84b8f833",
          6992 => x"83fab533",
          6993 => x"83fab222",
          6994 => x"72712912",
          6995 => x"5a5a4240",
          6996 => x"7883fab6",
          6997 => x"183483fa",
          6998 => x"b4336071",
          6999 => x"29620540",
          7000 => x"5a83fab0",
          7001 => x"337f86c7",
          7002 => x"b0800534",
          7003 => x"84b8f833",
          7004 => x"7081ff06",
          7005 => x"83fab222",
          7006 => x"83fab533",
          7007 => x"72722911",
          7008 => x"42405d58",
          7009 => x"5983fab0",
          7010 => x"338499d6",
          7011 => x"1f34811d",
          7012 => x"7081ff06",
          7013 => x"42587661",
          7014 => x"2681b838",
          7015 => x"84b8f933",
          7016 => x"5a7986f1",
          7017 => x"38ff1956",
          7018 => x"7583fab5",
          7019 => x"34800b84",
          7020 => x"bb840c9c",
          7021 => x"3d0d0478",
          7022 => x"b72e848a",
          7023 => x"38b77925",
          7024 => x"81fd3878",
          7025 => x"b82e9bb3",
          7026 => x"387880db",
          7027 => x"2e89cc38",
          7028 => x"800b84ba",
          7029 => x"800c84b8",
          7030 => x"f83383fa",
          7031 => x"b43383fa",
          7032 => x"b5337272",
          7033 => x"29055e40",
          7034 => x"4084b980",
          7035 => x"193386c7",
          7036 => x"a0801d34",
          7037 => x"84b8f833",
          7038 => x"83fab533",
          7039 => x"83fab222",
          7040 => x"72712912",
          7041 => x"415f5956",
          7042 => x"7883fab6",
          7043 => x"1f3483fa",
          7044 => x"b4337671",
          7045 => x"29195b57",
          7046 => x"83fab033",
          7047 => x"86c7b080",
          7048 => x"1b3484b8",
          7049 => x"f8337081",
          7050 => x"ff0683fa",
          7051 => x"b22283fa",
          7052 => x"b5337272",
          7053 => x"29114442",
          7054 => x"43585983",
          7055 => x"fab03360",
          7056 => x"8499d605",
          7057 => x"34811f58",
          7058 => x"7781ff06",
          7059 => x"41607727",
          7060 => x"feca3877",
          7061 => x"83fab534",
          7062 => x"800b84bb",
          7063 => x"840c9c3d",
          7064 => x"0d04789b",
          7065 => x"2e82b738",
          7066 => x"789b2483",
          7067 => x"8138788d",
          7068 => x"2e098106",
          7069 => x"fda83880",
          7070 => x"0b83fab5",
          7071 => x"34800b84",
          7072 => x"bb840c9c",
          7073 => x"3d0d0478",
          7074 => x"9b2e82aa",
          7075 => x"38d01956",
          7076 => x"75892684",
          7077 => x"d03884ba",
          7078 => x"84338111",
          7079 => x"59577784",
          7080 => x"ba843478",
          7081 => x"84ba8818",
          7082 => x"347781ff",
          7083 => x"0659800b",
          7084 => x"84ba881a",
          7085 => x"34800b84",
          7086 => x"bb840c9c",
          7087 => x"3d0d0478",
          7088 => x"9b2efde9",
          7089 => x"38800b84",
          7090 => x"ba800c84",
          7091 => x"b8f83383",
          7092 => x"fab43383",
          7093 => x"fab53372",
          7094 => x"7229055e",
          7095 => x"404084b9",
          7096 => x"80193386",
          7097 => x"c7a0801d",
          7098 => x"3484b8f8",
          7099 => x"3383fab5",
          7100 => x"3383fab2",
          7101 => x"22727129",
          7102 => x"12415f59",
          7103 => x"567883fa",
          7104 => x"b61f3483",
          7105 => x"fab43376",
          7106 => x"7129195b",
          7107 => x"5783fab0",
          7108 => x"3386c7b0",
          7109 => x"801b3484",
          7110 => x"b8f83370",
          7111 => x"81ff0683",
          7112 => x"fab22283",
          7113 => x"fab53372",
          7114 => x"72291144",
          7115 => x"42435859",
          7116 => x"83fab033",
          7117 => x"608499d6",
          7118 => x"0534811f",
          7119 => x"58fe8939",
          7120 => x"81528151",
          7121 => x"eafa3f80",
          7122 => x"0b83fab5",
          7123 => x"34feae39",
          7124 => x"84b8f833",
          7125 => x"83fab533",
          7126 => x"7081ff06",
          7127 => x"83fab433",
          7128 => x"73712912",
          7129 => x"86c7a080",
          7130 => x"0583fab2",
          7131 => x"2240515d",
          7132 => x"727e2905",
          7133 => x"7083ffff",
          7134 => x"0683f98a",
          7135 => x"335a5159",
          7136 => x"5a5c7581",
          7137 => x"2e86a438",
          7138 => x"7881ff06",
          7139 => x"ff1a5757",
          7140 => x"76fc9538",
          7141 => x"76567583",
          7142 => x"fab534fc",
          7143 => x"9039800b",
          7144 => x"84ba8434",
          7145 => x"800b84ba",
          7146 => x"8534800b",
          7147 => x"84ba8634",
          7148 => x"800b84ba",
          7149 => x"8734810b",
          7150 => x"84ba800c",
          7151 => x"800b84bb",
          7152 => x"840c9c3d",
          7153 => x"0d0483fa",
          7154 => x"b43384ba",
          7155 => x"ec3483fa",
          7156 => x"b53384ba",
          7157 => x"ed3483fa",
          7158 => x"b33384ba",
          7159 => x"ee34800b",
          7160 => x"84ba800c",
          7161 => x"800b84bb",
          7162 => x"840c9c3d",
          7163 => x"0d047880",
          7164 => x"ff2e0981",
          7165 => x"06faa738",
          7166 => x"83fab433",
          7167 => x"84b8f833",
          7168 => x"7081ff06",
          7169 => x"83fab533",
          7170 => x"7081ff06",
          7171 => x"72752911",
          7172 => x"86c7a080",
          7173 => x"0583fab2",
          7174 => x"225c4072",
          7175 => x"7b290570",
          7176 => x"83ffff06",
          7177 => x"83f98a33",
          7178 => x"445c435c",
          7179 => x"425b5c7d",
          7180 => x"812e85fe",
          7181 => x"387881ff",
          7182 => x"06ff1a58",
          7183 => x"56758338",
          7184 => x"75577683",
          7185 => x"fab5347b",
          7186 => x"81ff067a",
          7187 => x"81ff0678",
          7188 => x"81ff0672",
          7189 => x"7229055f",
          7190 => x"405b84b9",
          7191 => x"a03386c7",
          7192 => x"a0801e34",
          7193 => x"84b8f833",
          7194 => x"83fab533",
          7195 => x"83fab222",
          7196 => x"72712912",
          7197 => x"5a5e4240",
          7198 => x"a00b83fa",
          7199 => x"b6183483",
          7200 => x"fab43360",
          7201 => x"71296205",
          7202 => x"5a5683fa",
          7203 => x"b03386c7",
          7204 => x"b0801a34",
          7205 => x"84b8f833",
          7206 => x"7081ff06",
          7207 => x"83fab222",
          7208 => x"83fab533",
          7209 => x"72722911",
          7210 => x"435d5a5e",
          7211 => x"5983fab0",
          7212 => x"337f8499",
          7213 => x"d6053481",
          7214 => x"1a7081ff",
          7215 => x"065c587c",
          7216 => x"7b2695ea",
          7217 => x"3884b8f9",
          7218 => x"335a7996",
          7219 => x"d038ff19",
          7220 => x"587783fa",
          7221 => x"b53483fa",
          7222 => x"b5337081",
          7223 => x"ff0658ff",
          7224 => x"0556fdac",
          7225 => x"3978bb2e",
          7226 => x"95d83878",
          7227 => x"bd2e83d7",
          7228 => x"3878bf2e",
          7229 => x"95a83884",
          7230 => x"ba84335f",
          7231 => x"7e83f938",
          7232 => x"ffbf1956",
          7233 => x"75b42684",
          7234 => x"c8387510",
          7235 => x"1083c6e0",
          7236 => x"05587708",
          7237 => x"04800b83",
          7238 => x"fab53480",
          7239 => x"528151e7",
          7240 => x"9f3f800b",
          7241 => x"84bb840c",
          7242 => x"9c3d0d04",
          7243 => x"83fab433",
          7244 => x"84b8f833",
          7245 => x"7081ff06",
          7246 => x"83fab533",
          7247 => x"7081ff06",
          7248 => x"72752911",
          7249 => x"86c7a080",
          7250 => x"0583fab2",
          7251 => x"225c4172",
          7252 => x"7b290570",
          7253 => x"83ffff06",
          7254 => x"83f98a33",
          7255 => x"4653455c",
          7256 => x"595b5b7f",
          7257 => x"812e82ef",
          7258 => x"38805c7a",
          7259 => x"81ff067a",
          7260 => x"81ff067a",
          7261 => x"81ff0672",
          7262 => x"7229055c",
          7263 => x"584084b9",
          7264 => x"a03386c7",
          7265 => x"a0801b34",
          7266 => x"84b8f833",
          7267 => x"83fab533",
          7268 => x"83fab222",
          7269 => x"72712912",
          7270 => x"5e415e56",
          7271 => x"a00b83fa",
          7272 => x"b61c3483",
          7273 => x"fab43376",
          7274 => x"71291e5a",
          7275 => x"5e83fab0",
          7276 => x"3386c7b0",
          7277 => x"801a3484",
          7278 => x"b8f83370",
          7279 => x"81ff0683",
          7280 => x"fab22283",
          7281 => x"fab53372",
          7282 => x"7229115b",
          7283 => x"445a4059",
          7284 => x"83fab033",
          7285 => x"8499d618",
          7286 => x"34608105",
          7287 => x"7081ff06",
          7288 => x"5b587e7a",
          7289 => x"2681ac38",
          7290 => x"84b8f933",
          7291 => x"587792fb",
          7292 => x"38ff1956",
          7293 => x"7583fab5",
          7294 => x"34811c70",
          7295 => x"81ff065d",
          7296 => x"597b8326",
          7297 => x"f7a73883",
          7298 => x"fab43384",
          7299 => x"b8f83383",
          7300 => x"fab53372",
          7301 => x"81ff0672",
          7302 => x"81ff0672",
          7303 => x"81ff0672",
          7304 => x"72290554",
          7305 => x"5b435b5b",
          7306 => x"5b84b9a0",
          7307 => x"3386c7a0",
          7308 => x"801b3484",
          7309 => x"b8f83383",
          7310 => x"fab53383",
          7311 => x"fab22272",
          7312 => x"7129125e",
          7313 => x"415e56a0",
          7314 => x"0b83fab6",
          7315 => x"1c3483fa",
          7316 => x"b4337671",
          7317 => x"291e5a5e",
          7318 => x"83fab033",
          7319 => x"86c7b080",
          7320 => x"1a3484b8",
          7321 => x"f8337081",
          7322 => x"ff0683fa",
          7323 => x"b22283fa",
          7324 => x"b5337272",
          7325 => x"29115b44",
          7326 => x"5a405983",
          7327 => x"fab03384",
          7328 => x"99d61834",
          7329 => x"60810570",
          7330 => x"81ff065b",
          7331 => x"58797f27",
          7332 => x"fed63877",
          7333 => x"83fab534",
          7334 => x"fedf3982",
          7335 => x"0b84ba80",
          7336 => x"0c800b84",
          7337 => x"bb840c9c",
          7338 => x"3d0d0483",
          7339 => x"fab61733",
          7340 => x"5984b980",
          7341 => x"19337a34",
          7342 => x"83fab533",
          7343 => x"7081ff06",
          7344 => x"58ff0556",
          7345 => x"f9ca3981",
          7346 => x"0b84ba86",
          7347 => x"34800b84",
          7348 => x"bb840c9c",
          7349 => x"3d0d0483",
          7350 => x"fab61733",
          7351 => x"5b84b980",
          7352 => x"1b337c34",
          7353 => x"83fab433",
          7354 => x"84b8f833",
          7355 => x"83fab533",
          7356 => x"5b5b5b80",
          7357 => x"5cfcf439",
          7358 => x"84ba8842",
          7359 => x"9c3ddc11",
          7360 => x"53d80551",
          7361 => x"ff88ff3f",
          7362 => x"84bb8408",
          7363 => x"802efbf0",
          7364 => x"3884ba85",
          7365 => x"33811157",
          7366 => x"5a7584ba",
          7367 => x"85347910",
          7368 => x"83fe0641",
          7369 => x"0280ca05",
          7370 => x"226184ba",
          7371 => x"d80523fb",
          7372 => x"cf3983fa",
          7373 => x"b617335c",
          7374 => x"84b9801c",
          7375 => x"337b3483",
          7376 => x"fab43384",
          7377 => x"b8f83383",
          7378 => x"fab5335b",
          7379 => x"5b5cf9e5",
          7380 => x"3984b8f8",
          7381 => x"3383fab4",
          7382 => x"3383fab5",
          7383 => x"33727229",
          7384 => x"05415d5b",
          7385 => x"84b98019",
          7386 => x"337f86c7",
          7387 => x"a0800534",
          7388 => x"84b8f833",
          7389 => x"83fab533",
          7390 => x"83fab222",
          7391 => x"72712912",
          7392 => x"5a435b56",
          7393 => x"7883fab6",
          7394 => x"183483fa",
          7395 => x"b4337671",
          7396 => x"291b415e",
          7397 => x"83fab033",
          7398 => x"6086c7b0",
          7399 => x"80053484",
          7400 => x"b8f83370",
          7401 => x"81ff0683",
          7402 => x"fab22283",
          7403 => x"fab53372",
          7404 => x"72291141",
          7405 => x"5f5a425a",
          7406 => x"83fab033",
          7407 => x"8499d61e",
          7408 => x"34811c70",
          7409 => x"81ff065c",
          7410 => x"58607b26",
          7411 => x"90a23884",
          7412 => x"b8f93358",
          7413 => x"7790e238",
          7414 => x"ff1a5675",
          7415 => x"83fab534",
          7416 => x"800b84ba",
          7417 => x"800c84b8",
          7418 => x"fb33407f",
          7419 => x"802ef3bd",
          7420 => x"3884b8fc",
          7421 => x"335675f3",
          7422 => x"b4387852",
          7423 => x"8151eae4",
          7424 => x"3f800b84",
          7425 => x"bb840c9c",
          7426 => x"3d0d0484",
          7427 => x"baec3383",
          7428 => x"fab43484",
          7429 => x"baed3383",
          7430 => x"fab53484",
          7431 => x"baee3357",
          7432 => x"7683fab2",
          7433 => x"23ffb939",
          7434 => x"83fab433",
          7435 => x"84baec34",
          7436 => x"83fab533",
          7437 => x"84baed34",
          7438 => x"83fab333",
          7439 => x"84baee34",
          7440 => x"ff9e3984",
          7441 => x"ba85335b",
          7442 => x"7a802eff",
          7443 => x"933884ba",
          7444 => x"d8225d7c",
          7445 => x"862e0981",
          7446 => x"06ff8538",
          7447 => x"83fab533",
          7448 => x"81055583",
          7449 => x"fab43381",
          7450 => x"05549b53",
          7451 => x"83e5c052",
          7452 => x"943d7052",
          7453 => x"57feecb0",
          7454 => x"3f7651fe",
          7455 => x"fdaa3f84",
          7456 => x"bb840881",
          7457 => x"ff0683f9",
          7458 => x"88335776",
          7459 => x"054160a0",
          7460 => x"24fecd38",
          7461 => x"765283f8",
          7462 => x"e851fefb",
          7463 => x"f53ffec0",
          7464 => x"39800b84",
          7465 => x"ba85335b",
          7466 => x"587981ff",
          7467 => x"065b777b",
          7468 => x"27fead38",
          7469 => x"771084ba",
          7470 => x"d8058111",
          7471 => x"33574175",
          7472 => x"b1268aa5",
          7473 => x"38751010",
          7474 => x"83c8b405",
          7475 => x"5f7e0804",
          7476 => x"84ba8533",
          7477 => x"5e7d802e",
          7478 => x"8fa43883",
          7479 => x"fab43384",
          7480 => x"bad93371",
          7481 => x"71317009",
          7482 => x"709f2c72",
          7483 => x"065a4259",
          7484 => x"5e5c7583",
          7485 => x"fab434fd",
          7486 => x"e73984ba",
          7487 => x"85335675",
          7488 => x"802e8ee7",
          7489 => x"3884bad9",
          7490 => x"33ff0570",
          7491 => x"81ff0684",
          7492 => x"b8f8335d",
          7493 => x"575f757b",
          7494 => x"27fdc538",
          7495 => x"7583fab5",
          7496 => x"34fdbd39",
          7497 => x"800b83fa",
          7498 => x"b53483fa",
          7499 => x"b4337081",
          7500 => x"ff065d57",
          7501 => x"7b802efd",
          7502 => x"a738ff17",
          7503 => x"567583fa",
          7504 => x"b434fd9c",
          7505 => x"39800b83",
          7506 => x"fab53483",
          7507 => x"fab43384",
          7508 => x"b8f733ff",
          7509 => x"05575776",
          7510 => x"7625fd84",
          7511 => x"38811756",
          7512 => x"7583fab4",
          7513 => x"34fcf939",
          7514 => x"84ba8533",
          7515 => x"407f802e",
          7516 => x"8de03883",
          7517 => x"fab53384",
          7518 => x"bad93371",
          7519 => x"71317009",
          7520 => x"709f2c72",
          7521 => x"065a4159",
          7522 => x"425a7583",
          7523 => x"fab534fc",
          7524 => x"cf3984ba",
          7525 => x"85335b7a",
          7526 => x"802efcc4",
          7527 => x"3884bad8",
          7528 => x"22416099",
          7529 => x"2e098106",
          7530 => x"fcb63884",
          7531 => x"b8f83383",
          7532 => x"fab53383",
          7533 => x"fab43372",
          7534 => x"71291286",
          7535 => x"c7a08011",
          7536 => x"83fab222",
          7537 => x"43515a58",
          7538 => x"71602905",
          7539 => x"7083ffff",
          7540 => x"0683f988",
          7541 => x"0887fffe",
          7542 => x"8006425a",
          7543 => x"5d5d7e84",
          7544 => x"82802e92",
          7545 => x"bf38800b",
          7546 => x"83f98934",
          7547 => x"fbf23984",
          7548 => x"ba85335a",
          7549 => x"79802efb",
          7550 => x"e73884ba",
          7551 => x"d8225877",
          7552 => x"992e0981",
          7553 => x"06fbd938",
          7554 => x"810b83f9",
          7555 => x"8934fbd0",
          7556 => x"3984ba85",
          7557 => x"33567580",
          7558 => x"2e90be38",
          7559 => x"84bad933",
          7560 => x"83fab533",
          7561 => x"5d7c0584",
          7562 => x"b8f833ff",
          7563 => x"11595e56",
          7564 => x"757d2583",
          7565 => x"38755776",
          7566 => x"83fab534",
          7567 => x"fba23984",
          7568 => x"ba853357",
          7569 => x"76802e8c",
          7570 => x"c83884ba",
          7571 => x"d93383fa",
          7572 => x"b4334261",
          7573 => x"0584b8f7",
          7574 => x"33ff1159",
          7575 => x"41567560",
          7576 => x"25833875",
          7577 => x"577683fa",
          7578 => x"b434faf4",
          7579 => x"3983e5cc",
          7580 => x"51fee794",
          7581 => x"3f800b84",
          7582 => x"ba853357",
          7583 => x"57767627",
          7584 => x"8bc73876",
          7585 => x"1084bad8",
          7586 => x"05702253",
          7587 => x"5a83e5ac",
          7588 => x"51fee6f4",
          7589 => x"3f811770",
          7590 => x"81ff0684",
          7591 => x"ba853358",
          7592 => x"5858da39",
          7593 => x"820b84ba",
          7594 => x"85335f57",
          7595 => x"7d802e8d",
          7596 => x"3884bad8",
          7597 => x"22567583",
          7598 => x"26833875",
          7599 => x"57815276",
          7600 => x"81ff0651",
          7601 => x"d5f33ffa",
          7602 => x"973984ba",
          7603 => x"85335781",
          7604 => x"77278eb7",
          7605 => x"3884badb",
          7606 => x"33ff0570",
          7607 => x"81ff0684",
          7608 => x"bad933ff",
          7609 => x"057081ff",
          7610 => x"0684b8f7",
          7611 => x"337081ff",
          7612 => x"06ff1140",
          7613 => x"43525b59",
          7614 => x"5c5c777e",
          7615 => x"27833877",
          7616 => x"5a7983fa",
          7617 => x"b2237681",
          7618 => x"ff06ff18",
          7619 => x"585f777f",
          7620 => x"27833877",
          7621 => x"577683fa",
          7622 => x"b43484b8",
          7623 => x"f833ff11",
          7624 => x"57407a60",
          7625 => x"27f9b438",
          7626 => x"7a567583",
          7627 => x"fab534f9",
          7628 => x"af3984ba",
          7629 => x"85335f7e",
          7630 => x"802e8aef",
          7631 => x"3884bad9",
          7632 => x"3384b8f7",
          7633 => x"33405b7a",
          7634 => x"7f26f994",
          7635 => x"3883fab4",
          7636 => x"3384b8f8",
          7637 => x"337081ff",
          7638 => x"0683fab5",
          7639 => x"33717429",
          7640 => x"1186c7a0",
          7641 => x"800583fa",
          7642 => x"b2225f40",
          7643 => x"717e2905",
          7644 => x"7083ffff",
          7645 => x"0683f98a",
          7646 => x"33465259",
          7647 => x"595f5d60",
          7648 => x"812e84f0",
          7649 => x"387983ff",
          7650 => x"ff06707c",
          7651 => x"315d5780",
          7652 => x"7c248efe",
          7653 => x"3884b8f7",
          7654 => x"33567676",
          7655 => x"278ed638",
          7656 => x"ff165675",
          7657 => x"83fab223",
          7658 => x"7c81ff06",
          7659 => x"707c3141",
          7660 => x"57806024",
          7661 => x"8ee53884",
          7662 => x"b8f73356",
          7663 => x"7676278d",
          7664 => x"ee38ff16",
          7665 => x"567583fa",
          7666 => x"b4347e81",
          7667 => x"ff0683fa",
          7668 => x"b2225757",
          7669 => x"805a7676",
          7670 => x"26903875",
          7671 => x"77318105",
          7672 => x"7e81ff06",
          7673 => x"7171295c",
          7674 => x"5e5b7958",
          7675 => x"86c7a080",
          7676 => x"5b86c7b0",
          7677 => x"807f81ff",
          7678 => x"067f81ff",
          7679 => x"06717129",
          7680 => x"1d425842",
          7681 => x"5c797f27",
          7682 => x"f7d63884",
          7683 => x"99d61a57",
          7684 => x"e0e01733",
          7685 => x"5f84b980",
          7686 => x"1f337b70",
          7687 => x"81055d34",
          7688 => x"76708105",
          7689 => x"58337c70",
          7690 => x"81055e34",
          7691 => x"811884b8",
          7692 => x"f83384b8",
          7693 => x"f7337171",
          7694 => x"291d4340",
          7695 => x"5e587760",
          7696 => x"27f79d38",
          7697 => x"e0e01733",
          7698 => x"5f84b980",
          7699 => x"1f337b70",
          7700 => x"81055d34",
          7701 => x"76708105",
          7702 => x"58337c70",
          7703 => x"81055e34",
          7704 => x"811884b8",
          7705 => x"f83384b8",
          7706 => x"f7337171",
          7707 => x"291d4340",
          7708 => x"5e587f78",
          7709 => x"26ff9938",
          7710 => x"f6e63984",
          7711 => x"ba853356",
          7712 => x"75802e87",
          7713 => x"e0388052",
          7714 => x"84bad933",
          7715 => x"51d8b13f",
          7716 => x"f6ce3980",
          7717 => x"0b84b8f8",
          7718 => x"33ff1184",
          7719 => x"ba85335d",
          7720 => x"59405879",
          7721 => x"782e9438",
          7722 => x"84bad822",
          7723 => x"5675782e",
          7724 => x"0981068b",
          7725 => x"be3883fa",
          7726 => x"b5335876",
          7727 => x"81ff0683",
          7728 => x"fab43379",
          7729 => x"435c5c76",
          7730 => x"ff2e81ed",
          7731 => x"3884b8f7",
          7732 => x"33407a60",
          7733 => x"26f68938",
          7734 => x"7e81ff06",
          7735 => x"56607626",
          7736 => x"f5fe387b",
          7737 => x"7626617d",
          7738 => x"27075776",
          7739 => x"f5f2387a",
          7740 => x"10101b70",
          7741 => x"90296205",
          7742 => x"86c7a080",
          7743 => x"11701f5d",
          7744 => x"5a86c7b0",
          7745 => x"80057983",
          7746 => x"0658515d",
          7747 => x"758bac38",
          7748 => x"79830657",
          7749 => x"768ba438",
          7750 => x"83fab033",
          7751 => x"70982b71",
          7752 => x"902b0771",
          7753 => x"882b0771",
          7754 => x"07797f59",
          7755 => x"525f5777",
          7756 => x"7a279e38",
          7757 => x"80777084",
          7758 => x"05590c7d",
          7759 => x"76708405",
          7760 => x"580c7977",
          7761 => x"26ee3884",
          7762 => x"b8f83384",
          7763 => x"b8f73341",
          7764 => x"5f7e81ff",
          7765 => x"066081ff",
          7766 => x"0683fab2",
          7767 => x"227d7329",
          7768 => x"64055959",
          7769 => x"595a7777",
          7770 => x"268c3876",
          7771 => x"78311b70",
          7772 => x"7b296205",
          7773 => x"57407576",
          7774 => x"1d575776",
          7775 => x"7626f4e0",
          7776 => x"3883fab0",
          7777 => x"338499d6",
          7778 => x"18595aa0",
          7779 => x"0be0e019",
          7780 => x"34797870",
          7781 => x"81055a34",
          7782 => x"81175776",
          7783 => x"7626f4c0",
          7784 => x"38a00be0",
          7785 => x"e0193479",
          7786 => x"78708105",
          7787 => x"5a348117",
          7788 => x"57757727",
          7789 => x"d638f4a8",
          7790 => x"39ff1f70",
          7791 => x"81ff065d",
          7792 => x"58fe8a39",
          7793 => x"83fab033",
          7794 => x"7080f006",
          7795 => x"71842b80",
          7796 => x"f0067184",
          7797 => x"2a07585d",
          7798 => x"577b80f0",
          7799 => x"2e098106",
          7800 => x"be3880f2",
          7801 => x"0b83fab0",
          7802 => x"34811870",
          7803 => x"81ff0659",
          7804 => x"56f5b639",
          7805 => x"83fab617",
          7806 => x"335e84b9",
          7807 => x"801e337c",
          7808 => x"3483fab4",
          7809 => x"3384b8f8",
          7810 => x"3383fab2",
          7811 => x"2284b8f7",
          7812 => x"33425c5f",
          7813 => x"5dfaee39",
          7814 => x"83fab033",
          7815 => x"87075675",
          7816 => x"83fab034",
          7817 => x"81187081",
          7818 => x"ff065956",
          7819 => x"f4fb3983",
          7820 => x"fab03381",
          7821 => x"fd068507",
          7822 => x"567583fa",
          7823 => x"b034e539",
          7824 => x"83fab033",
          7825 => x"81fb0683",
          7826 => x"07567583",
          7827 => x"fab034d4",
          7828 => x"3983fab0",
          7829 => x"3381f906",
          7830 => x"81075675",
          7831 => x"83fab034",
          7832 => x"c33983fa",
          7833 => x"b033819f",
          7834 => x"06900756",
          7835 => x"7583fab0",
          7836 => x"34ffb139",
          7837 => x"80f10b83",
          7838 => x"fab03481",
          7839 => x"187081ff",
          7840 => x"065956f4",
          7841 => x"a43983fa",
          7842 => x"b033818f",
          7843 => x"06567583",
          7844 => x"fab034ff",
          7845 => x"8f3983fa",
          7846 => x"b033819f",
          7847 => x"06900756",
          7848 => x"7583fab0",
          7849 => x"34fefd39",
          7850 => x"83fab033",
          7851 => x"81ef0680",
          7852 => x"e0075675",
          7853 => x"83fab034",
          7854 => x"feea3983",
          7855 => x"fab03381",
          7856 => x"cf0680c0",
          7857 => x"07567583",
          7858 => x"fab034fe",
          7859 => x"d73983fa",
          7860 => x"b03381af",
          7861 => x"06a00756",
          7862 => x"7583fab0",
          7863 => x"34fec539",
          7864 => x"83fab033",
          7865 => x"81fe0686",
          7866 => x"07567583",
          7867 => x"fab034fe",
          7868 => x"b33983fa",
          7869 => x"b03381fc",
          7870 => x"06840756",
          7871 => x"7583fab0",
          7872 => x"34fea139",
          7873 => x"83fab033",
          7874 => x"81fa0682",
          7875 => x"07567583",
          7876 => x"fab034fe",
          7877 => x"8f3983fa",
          7878 => x"b03381f8",
          7879 => x"06567583",
          7880 => x"fab034fd",
          7881 => x"ff3983fa",
          7882 => x"b03380f0",
          7883 => x"07567583",
          7884 => x"fab034fd",
          7885 => x"ef3983fa",
          7886 => x"b03380f0",
          7887 => x"07567583",
          7888 => x"fab034fd",
          7889 => x"df3983fa",
          7890 => x"b03381df",
          7891 => x"0680d007",
          7892 => x"567583fa",
          7893 => x"b034fdcc",
          7894 => x"3983fab0",
          7895 => x"3381bf06",
          7896 => x"b0075675",
          7897 => x"83fab034",
          7898 => x"fdba3980",
          7899 => x"0b83fab5",
          7900 => x"34805281",
          7901 => x"51d2c93f",
          7902 => x"ecff3984",
          7903 => x"baec3383",
          7904 => x"fab43484",
          7905 => x"baed3383",
          7906 => x"fab53484",
          7907 => x"baee3359",
          7908 => x"7883fab2",
          7909 => x"23800b84",
          7910 => x"ba800ce8",
          7911 => x"c739810b",
          7912 => x"84ba8734",
          7913 => x"800b84bb",
          7914 => x"840c9c3d",
          7915 => x"0d047783",
          7916 => x"fab53483",
          7917 => x"fab53370",
          7918 => x"81ff0658",
          7919 => x"ff0556e7",
          7920 => x"cf3984ba",
          7921 => x"88429c3d",
          7922 => x"dc1153d8",
          7923 => x"0551fef7",
          7924 => x"b53f84bb",
          7925 => x"8408a138",
          7926 => x"84bb8408",
          7927 => x"84ba800c",
          7928 => x"800b84ba",
          7929 => x"8434800b",
          7930 => x"84bb840c",
          7931 => x"9c3d0d04",
          7932 => x"7783fab5",
          7933 => x"34efe939",
          7934 => x"84ba8533",
          7935 => x"81115c5c",
          7936 => x"7a84ba85",
          7937 => x"347b1083",
          7938 => x"fe065d02",
          7939 => x"80ca0522",
          7940 => x"84bad81e",
          7941 => x"23800b84",
          7942 => x"ba8434ca",
          7943 => x"39800b83",
          7944 => x"fab53480",
          7945 => x"528151d1",
          7946 => x"973f83fa",
          7947 => x"b5337081",
          7948 => x"ff0658ff",
          7949 => x"0556e6d8",
          7950 => x"39800b83",
          7951 => x"fab53480",
          7952 => x"528151d0",
          7953 => x"fb3fef98",
          7954 => x"398a51fe",
          7955 => x"ea903fef",
          7956 => x"8f3983fa",
          7957 => x"b533ff05",
          7958 => x"7009709f",
          7959 => x"2c720658",
          7960 => x"5f57f2a6",
          7961 => x"39755281",
          7962 => x"51d93984",
          7963 => x"b8f83340",
          7964 => x"756027ee",
          7965 => x"eb387583",
          7966 => x"fab534ee",
          7967 => x"e33983fa",
          7968 => x"b433ff05",
          7969 => x"7009709f",
          7970 => x"2c720658",
          7971 => x"4057f0e2",
          7972 => x"3983fab4",
          7973 => x"33810584",
          7974 => x"b8f733ff",
          7975 => x"11595956",
          7976 => x"757825f3",
          7977 => x"c0387557",
          7978 => x"f3bb3984",
          7979 => x"b8f73370",
          7980 => x"81ff0658",
          7981 => x"5c817726",
          7982 => x"eea63883",
          7983 => x"fab43384",
          7984 => x"b8f83370",
          7985 => x"81ff0683",
          7986 => x"fab53371",
          7987 => x"74291186",
          7988 => x"c7a08005",
          7989 => x"83fab222",
          7990 => x"5f5f717e",
          7991 => x"29057083",
          7992 => x"ffff0683",
          7993 => x"f98a335d",
          7994 => x"5b44425f",
          7995 => x"5d77812e",
          7996 => x"81f53879",
          7997 => x"83ffff06",
          7998 => x"ff115c57",
          7999 => x"807b2484",
          8000 => x"893884b8",
          8001 => x"f7335676",
          8002 => x"76278398",
          8003 => x"38ff1656",
          8004 => x"7583fab2",
          8005 => x"237c81ff",
          8006 => x"06ff1157",
          8007 => x"57807624",
          8008 => x"83df3884",
          8009 => x"b8f73356",
          8010 => x"76762782",
          8011 => x"ec38ff16",
          8012 => x"567583fa",
          8013 => x"b4347b81",
          8014 => x"ff0683fa",
          8015 => x"b2225757",
          8016 => x"805a7676",
          8017 => x"26903875",
          8018 => x"77318105",
          8019 => x"7e81ff06",
          8020 => x"7171295c",
          8021 => x"5e5f7958",
          8022 => x"86c7a080",
          8023 => x"5b86c7b0",
          8024 => x"807c81ff",
          8025 => x"067f81ff",
          8026 => x"06717129",
          8027 => x"1d414242",
          8028 => x"5d797e27",
          8029 => x"ecea3884",
          8030 => x"99d61a57",
          8031 => x"e0e01733",
          8032 => x"5e84b980",
          8033 => x"1e337b70",
          8034 => x"81055d34",
          8035 => x"76708105",
          8036 => x"58337d70",
          8037 => x"81055f34",
          8038 => x"811884b8",
          8039 => x"f83384b8",
          8040 => x"f7337171",
          8041 => x"291d5941",
          8042 => x"5d587776",
          8043 => x"27ecb138",
          8044 => x"e0e01733",
          8045 => x"5e84b980",
          8046 => x"1e337b70",
          8047 => x"81055d34",
          8048 => x"76708105",
          8049 => x"58337d70",
          8050 => x"81055f34",
          8051 => x"811884b8",
          8052 => x"f83384b8",
          8053 => x"f7337171",
          8054 => x"291d5941",
          8055 => x"5d587578",
          8056 => x"26ff9938",
          8057 => x"ebfa3983",
          8058 => x"fab61733",
          8059 => x"5c84b980",
          8060 => x"1c337b34",
          8061 => x"83fab433",
          8062 => x"84b8f833",
          8063 => x"83fab222",
          8064 => x"84b8f733",
          8065 => x"5f5c5f5d",
          8066 => x"fde93976",
          8067 => x"ebd23884",
          8068 => x"b8f73370",
          8069 => x"81ff06ff",
          8070 => x"115c4258",
          8071 => x"76612783",
          8072 => x"38765a79",
          8073 => x"83fab223",
          8074 => x"7781ff06",
          8075 => x"ff19585a",
          8076 => x"807a2783",
          8077 => x"38805776",
          8078 => x"83fab434",
          8079 => x"84b8f833",
          8080 => x"7081ff06",
          8081 => x"ff125259",
          8082 => x"56807827",
          8083 => x"eb8d3880",
          8084 => x"567583fa",
          8085 => x"b534eb88",
          8086 => x"3983fab5",
          8087 => x"33810584",
          8088 => x"b8f833ff",
          8089 => x"11594056",
          8090 => x"757f25ef",
          8091 => x"ca387557",
          8092 => x"efc53975",
          8093 => x"812e0981",
          8094 => x"06f4c038",
          8095 => x"83fab533",
          8096 => x"7081ff06",
          8097 => x"83fab433",
          8098 => x"7a445d5d",
          8099 => x"5776ff2e",
          8100 => x"098106f4",
          8101 => x"b838f6a1",
          8102 => x"39ff1d56",
          8103 => x"7583fab4",
          8104 => x"34fd9339",
          8105 => x"ff1a5675",
          8106 => x"83fab223",
          8107 => x"fce7397c",
          8108 => x"7b315675",
          8109 => x"83fab434",
          8110 => x"f2903977",
          8111 => x"7d585677",
          8112 => x"7a26f58d",
          8113 => x"38807670",
          8114 => x"81055834",
          8115 => x"83fab033",
          8116 => x"77708105",
          8117 => x"5934757a",
          8118 => x"26f4ec38",
          8119 => x"80767081",
          8120 => x"05583483",
          8121 => x"fab03377",
          8122 => x"70810559",
          8123 => x"34797627",
          8124 => x"d438f4d3",
          8125 => x"39797b31",
          8126 => x"567583fa",
          8127 => x"b223f1a8",
          8128 => x"39800b83",
          8129 => x"fab434fc",
          8130 => x"ad397e83",
          8131 => x"fab223fc",
          8132 => x"8439800b",
          8133 => x"83fab223",
          8134 => x"f18e3980",
          8135 => x"0b83fab4",
          8136 => x"34f1a739",
          8137 => x"83fab618",
          8138 => x"335a84b9",
          8139 => x"801a3377",
          8140 => x"34800b83",
          8141 => x"f98934e9",
          8142 => x"a739fd3d",
          8143 => x"0d029705",
          8144 => x"3384b8fa",
          8145 => x"33545472",
          8146 => x"802e9038",
          8147 => x"7351db9c",
          8148 => x"3f800b84",
          8149 => x"bb840c85",
          8150 => x"3d0d0476",
          8151 => x"527351d7",
          8152 => x"ab3f800b",
          8153 => x"84bb840c",
          8154 => x"853d0d04",
          8155 => x"f33d0d02",
          8156 => x"bf05335c",
          8157 => x"ff0b83f9",
          8158 => x"88337081",
          8159 => x"ff0683f8",
          8160 => x"e8113358",
          8161 => x"55555974",
          8162 => x"802e80d6",
          8163 => x"38811456",
          8164 => x"7583f988",
          8165 => x"34745978",
          8166 => x"84bb840c",
          8167 => x"8f3d0d04",
          8168 => x"83f8e408",
          8169 => x"54825373",
          8170 => x"802e9138",
          8171 => x"73733270",
          8172 => x"30710770",
          8173 => x"09709f2a",
          8174 => x"565d5e58",
          8175 => x"7283f8e4",
          8176 => x"0cff5980",
          8177 => x"547b812e",
          8178 => x"09810683",
          8179 => x"387b547b",
          8180 => x"83327030",
          8181 => x"70802576",
          8182 => x"075c5c5d",
          8183 => x"79802e85",
          8184 => x"c43884b8",
          8185 => x"f83383fa",
          8186 => x"b53383fa",
          8187 => x"b4337271",
          8188 => x"291286c7",
          8189 => x"a0800583",
          8190 => x"fab2225b",
          8191 => x"595d7179",
          8192 => x"29057083",
          8193 => x"ffff0683",
          8194 => x"f9893358",
          8195 => x"59555874",
          8196 => x"812e838c",
          8197 => x"3881f054",
          8198 => x"73878e80",
          8199 => x"8034800b",
          8200 => x"87c09888",
          8201 => x"0c87c098",
          8202 => x"88085675",
          8203 => x"802ef638",
          8204 => x"878e8084",
          8205 => x"08577683",
          8206 => x"f6b41534",
          8207 => x"81147081",
          8208 => x"ff065555",
          8209 => x"81f97427",
          8210 => x"cf388054",
          8211 => x"83f8a414",
          8212 => x"337081ff",
          8213 => x"0683f8ae",
          8214 => x"16335854",
          8215 => x"5572762e",
          8216 => x"85c13872",
          8217 => x"81ff2e86",
          8218 => x"b4387483",
          8219 => x"f8b81534",
          8220 => x"7581ff06",
          8221 => x"5a7981ff",
          8222 => x"2e85cd38",
          8223 => x"7583f8c2",
          8224 => x"153483f8",
          8225 => x"a4143383",
          8226 => x"f8ae1534",
          8227 => x"81147081",
          8228 => x"ff06555e",
          8229 => x"897427ff",
          8230 => x"b33883f8",
          8231 => x"ac337098",
          8232 => x"2b708025",
          8233 => x"58565475",
          8234 => x"83f8dc34",
          8235 => x"7381ff06",
          8236 => x"70862a81",
          8237 => x"32708106",
          8238 => x"51545872",
          8239 => x"802e85e7",
          8240 => x"38810b83",
          8241 => x"f8dd3473",
          8242 => x"09810653",
          8243 => x"72802e85",
          8244 => x"e438810b",
          8245 => x"83f8de34",
          8246 => x"800b83f8",
          8247 => x"dd3383f8",
          8248 => x"e40883f8",
          8249 => x"de337083",
          8250 => x"f8e03383",
          8251 => x"f8df335d",
          8252 => x"5d425e5c",
          8253 => x"5e5683f8",
          8254 => x"b8163355",
          8255 => x"7481ff2e",
          8256 => x"8d3883f8",
          8257 => x"cc163354",
          8258 => x"73802e82",
          8259 => x"823883f8",
          8260 => x"c2163353",
          8261 => x"7281ff2e",
          8262 => x"8b3883f8",
          8263 => x"cc163354",
          8264 => x"7381ec38",
          8265 => x"7481ff06",
          8266 => x"547381ff",
          8267 => x"2e8d3883",
          8268 => x"f8cc1633",
          8269 => x"5372812e",
          8270 => x"81da3874",
          8271 => x"81ff0653",
          8272 => x"7281ff2e",
          8273 => x"848c3883",
          8274 => x"f8cc1633",
          8275 => x"54817427",
          8276 => x"84803883",
          8277 => x"f8d80887",
          8278 => x"e80587c0",
          8279 => x"989c0854",
          8280 => x"54737327",
          8281 => x"83ec3881",
          8282 => x"0b87c098",
          8283 => x"9c0883f8",
          8284 => x"d80c5881",
          8285 => x"167081ff",
          8286 => x"06575489",
          8287 => x"7627fef6",
          8288 => x"387683f8",
          8289 => x"df347783",
          8290 => x"f8e034fe",
          8291 => x"9e195372",
          8292 => x"9c26828b",
          8293 => x"38721010",
          8294 => x"83c9fc05",
          8295 => x"5a790804",
          8296 => x"83f98c08",
          8297 => x"5473802e",
          8298 => x"913883f4",
          8299 => x"1487c098",
          8300 => x"9c085e5e",
          8301 => x"7d7d27fc",
          8302 => x"dc38800b",
          8303 => x"83f98a33",
          8304 => x"54547281",
          8305 => x"2e833874",
          8306 => x"547383f9",
          8307 => x"8a3487c0",
          8308 => x"989c0883",
          8309 => x"f98c0c73",
          8310 => x"81ff0658",
          8311 => x"77812e94",
          8312 => x"3883fab6",
          8313 => x"17335484",
          8314 => x"b9801433",
          8315 => x"763481f0",
          8316 => x"54fca539",
          8317 => x"83f8e408",
          8318 => x"5372802e",
          8319 => x"829c3872",
          8320 => x"812e83f4",
          8321 => x"3880c376",
          8322 => x"3481f054",
          8323 => x"fc8a3980",
          8324 => x"58fee039",
          8325 => x"80745657",
          8326 => x"83597c81",
          8327 => x"2e9b3879",
          8328 => x"772e0981",
          8329 => x"0683b438",
          8330 => x"7d812e80",
          8331 => x"ed387981",
          8332 => x"2e80d738",
          8333 => x"7981ff06",
          8334 => x"59877727",
          8335 => x"75982b54",
          8336 => x"54728025",
          8337 => x"a1387380",
          8338 => x"2e9c3881",
          8339 => x"177081ff",
          8340 => x"06761081",
          8341 => x"fe068772",
          8342 => x"2771982b",
          8343 => x"57535758",
          8344 => x"54807324",
          8345 => x"e1387810",
          8346 => x"10107910",
          8347 => x"05761183",
          8348 => x"2b780583",
          8349 => x"f5940570",
          8350 => x"335b5654",
          8351 => x"7887c098",
          8352 => x"9c0883f8",
          8353 => x"d80c57fd",
          8354 => x"ea398059",
          8355 => x"7d812eff",
          8356 => x"a8387981",
          8357 => x"ff0659ff",
          8358 => x"a0398259",
          8359 => x"ff9b3978",
          8360 => x"ff2efa9f",
          8361 => x"38800b84",
          8362 => x"b8fa3354",
          8363 => x"5472812e",
          8364 => x"83e8387b",
          8365 => x"82327030",
          8366 => x"70802576",
          8367 => x"07405956",
          8368 => x"7d8a387b",
          8369 => x"832e0981",
          8370 => x"06f9cc38",
          8371 => x"78ff2ef9",
          8372 => x"c6388053",
          8373 => x"72101010",
          8374 => x"83f99005",
          8375 => x"70335d54",
          8376 => x"787c2e83",
          8377 => x"ba388113",
          8378 => x"7081ff06",
          8379 => x"54579373",
          8380 => x"27e23884",
          8381 => x"b8fb3353",
          8382 => x"72802ef9",
          8383 => x"9a3884b8",
          8384 => x"fc335574",
          8385 => x"f9913878",
          8386 => x"81ff0652",
          8387 => x"8251ccd4",
          8388 => x"3f7884bb",
          8389 => x"840c8f3d",
          8390 => x"0d04be76",
          8391 => x"3481f054",
          8392 => x"f9f63972",
          8393 => x"81ff2e92",
          8394 => x"3883f8cc",
          8395 => x"14338105",
          8396 => x"5b7a83f8",
          8397 => x"cc1534fa",
          8398 => x"c939800b",
          8399 => x"83f8cc15",
          8400 => x"34ff0b83",
          8401 => x"f8b81534",
          8402 => x"ff0b83f8",
          8403 => x"c21534fa",
          8404 => x"b1397481",
          8405 => x"ff065372",
          8406 => x"81ff2efc",
          8407 => x"963883f8",
          8408 => x"cc163355",
          8409 => x"817527fc",
          8410 => x"8a387781",
          8411 => x"ff065473",
          8412 => x"812e0981",
          8413 => x"06fbfc38",
          8414 => x"83f8d808",
          8415 => x"81fa0587",
          8416 => x"c0989c08",
          8417 => x"54557473",
          8418 => x"27fbe838",
          8419 => x"87c0989c",
          8420 => x"0883f8d8",
          8421 => x"0c7681ff",
          8422 => x"0659fbd7",
          8423 => x"39ff0b83",
          8424 => x"f8b81534",
          8425 => x"f9ca3972",
          8426 => x"83f8dd34",
          8427 => x"73098106",
          8428 => x"5372fa9e",
          8429 => x"387283f8",
          8430 => x"de34800b",
          8431 => x"83f8dd33",
          8432 => x"83f8e408",
          8433 => x"83f8de33",
          8434 => x"7083f8e0",
          8435 => x"3383f8df",
          8436 => x"335d5d42",
          8437 => x"5e5c5e56",
          8438 => x"fa9c3979",
          8439 => x"822e0981",
          8440 => x"06fccb38",
          8441 => x"7a597a81",
          8442 => x"2efcce38",
          8443 => x"79812e09",
          8444 => x"8106fcc0",
          8445 => x"38fd9339",
          8446 => x"ef763481",
          8447 => x"f054f898",
          8448 => x"39800b84",
          8449 => x"b8fb3357",
          8450 => x"54758338",
          8451 => x"81547384",
          8452 => x"b8fb34ff",
          8453 => x"59f7ac39",
          8454 => x"800b84b8",
          8455 => x"fa335854",
          8456 => x"76833881",
          8457 => x"547384b8",
          8458 => x"fa34ff59",
          8459 => x"f7953981",
          8460 => x"5383f8e4",
          8461 => x"08842ef7",
          8462 => x"8338840b",
          8463 => x"83f8e40c",
          8464 => x"f6ff3984",
          8465 => x"b8f73370",
          8466 => x"81ff06ff",
          8467 => x"11575a54",
          8468 => x"80792783",
          8469 => x"38805574",
          8470 => x"83fab223",
          8471 => x"7381ff06",
          8472 => x"ff155553",
          8473 => x"80732783",
          8474 => x"38805473",
          8475 => x"83fab434",
          8476 => x"84b8f833",
          8477 => x"7081ff06",
          8478 => x"56ff0553",
          8479 => x"80752783",
          8480 => x"38805372",
          8481 => x"83fab534",
          8482 => x"ff59f6b7",
          8483 => x"39815283",
          8484 => x"51ffbaa5",
          8485 => x"3fff59f6",
          8486 => x"aa397254",
          8487 => x"fc953984",
          8488 => x"14085283",
          8489 => x"f8e851fe",
          8490 => x"dd9d3f81",
          8491 => x"0b83f988",
          8492 => x"3483f8e8",
          8493 => x"3359fcbb",
          8494 => x"39803d0d",
          8495 => x"8151f5ac",
          8496 => x"3f823d0d",
          8497 => x"04fa3d0d",
          8498 => x"800b83f5",
          8499 => x"90085357",
          8500 => x"02a30533",
          8501 => x"82133483",
          8502 => x"f5900851",
          8503 => x"80e07134",
          8504 => x"850b83f5",
          8505 => x"90085556",
          8506 => x"fe0b8115",
          8507 => x"34800b87",
          8508 => x"9080e834",
          8509 => x"87c0989c",
          8510 => x"0883f590",
          8511 => x"085580ce",
          8512 => x"90055387",
          8513 => x"c0989c08",
          8514 => x"5287c098",
          8515 => x"9c085170",
          8516 => x"722ef638",
          8517 => x"81143387",
          8518 => x"c0989c08",
          8519 => x"56527473",
          8520 => x"27873871",
          8521 => x"81fe2edb",
          8522 => x"3887c098",
          8523 => x"a40851ff",
          8524 => x"55707327",
          8525 => x"80c83871",
          8526 => x"5571ff2e",
          8527 => x"80c03887",
          8528 => x"c0989c08",
          8529 => x"80ce9005",
          8530 => x"5387c098",
          8531 => x"9c085287",
          8532 => x"c0989c08",
          8533 => x"5574722e",
          8534 => x"f6388114",
          8535 => x"3387c098",
          8536 => x"9c085252",
          8537 => x"70732787",
          8538 => x"387181ff",
          8539 => x"2edb3887",
          8540 => x"c098a408",
          8541 => x"55727526",
          8542 => x"8338ff52",
          8543 => x"7155ff16",
          8544 => x"7081ff06",
          8545 => x"57537580",
          8546 => x"2e983874",
          8547 => x"81ff0652",
          8548 => x"71fed538",
          8549 => x"74ff2e8a",
          8550 => x"387684bb",
          8551 => x"840c883d",
          8552 => x"0d04810b",
          8553 => x"84bb840c",
          8554 => x"883d0d04",
          8555 => x"fa3d0d79",
          8556 => x"028405a3",
          8557 => x"05335652",
          8558 => x"800b83f5",
          8559 => x"90087388",
          8560 => x"2b87fc80",
          8561 => x"80067075",
          8562 => x"982a0751",
          8563 => x"55555771",
          8564 => x"83153472",
          8565 => x"902a5170",
          8566 => x"84153471",
          8567 => x"902a5675",
          8568 => x"85153472",
          8569 => x"86153483",
          8570 => x"f5900852",
          8571 => x"74821334",
          8572 => x"83f59008",
          8573 => x"5180e171",
          8574 => x"34850b83",
          8575 => x"f5900855",
          8576 => x"56fe0b81",
          8577 => x"1534800b",
          8578 => x"879080e8",
          8579 => x"3487c098",
          8580 => x"9c0883f5",
          8581 => x"90085580",
          8582 => x"ce900553",
          8583 => x"87c0989c",
          8584 => x"085287c0",
          8585 => x"989c0851",
          8586 => x"70722ef6",
          8587 => x"38811433",
          8588 => x"87c0989c",
          8589 => x"08565274",
          8590 => x"73278738",
          8591 => x"7181fe2e",
          8592 => x"db3887c0",
          8593 => x"98a40851",
          8594 => x"ff557073",
          8595 => x"2780c838",
          8596 => x"715571ff",
          8597 => x"2e80c038",
          8598 => x"87c0989c",
          8599 => x"0880ce90",
          8600 => x"055387c0",
          8601 => x"989c0852",
          8602 => x"87c0989c",
          8603 => x"08557472",
          8604 => x"2ef63881",
          8605 => x"143387c0",
          8606 => x"989c0852",
          8607 => x"52707327",
          8608 => x"87387181",
          8609 => x"ff2edb38",
          8610 => x"87c098a4",
          8611 => x"08557275",
          8612 => x"268338ff",
          8613 => x"527155ff",
          8614 => x"167081ff",
          8615 => x"06575375",
          8616 => x"802e80c7",
          8617 => x"387481ff",
          8618 => x"065271fe",
          8619 => x"d4387451",
          8620 => x"7081ff06",
          8621 => x"5675aa38",
          8622 => x"80c6147b",
          8623 => x"84801155",
          8624 => x"52527073",
          8625 => x"27923871",
          8626 => x"70810553",
          8627 => x"33717081",
          8628 => x"05533472",
          8629 => x"7126f038",
          8630 => x"7684bb84",
          8631 => x"0c883d0d",
          8632 => x"04810b84",
          8633 => x"bb840c88",
          8634 => x"3d0d04ff",
          8635 => x"51c239fa",
          8636 => x"3d0d7902",
          8637 => x"8405a305",
          8638 => x"33565680",
          8639 => x"0b83f590",
          8640 => x"0877882b",
          8641 => x"87fc8080",
          8642 => x"06707998",
          8643 => x"2a075155",
          8644 => x"55577583",
          8645 => x"15347290",
          8646 => x"2a517084",
          8647 => x"15347590",
          8648 => x"2a527185",
          8649 => x"15347286",
          8650 => x"15347a83",
          8651 => x"f5900880",
          8652 => x"c6118480",
          8653 => x"13565455",
          8654 => x"51707327",
          8655 => x"97387070",
          8656 => x"81055233",
          8657 => x"72708105",
          8658 => x"54347271",
          8659 => x"26f03883",
          8660 => x"f5900854",
          8661 => x"74821534",
          8662 => x"83f59008",
          8663 => x"5580e275",
          8664 => x"34850b83",
          8665 => x"f5900855",
          8666 => x"56fe0b81",
          8667 => x"1534800b",
          8668 => x"879080e8",
          8669 => x"3487c098",
          8670 => x"9c0883f5",
          8671 => x"90085580",
          8672 => x"ce900553",
          8673 => x"87c0989c",
          8674 => x"085287c0",
          8675 => x"989c0851",
          8676 => x"70722ef6",
          8677 => x"38811433",
          8678 => x"87c0989c",
          8679 => x"08565274",
          8680 => x"73278738",
          8681 => x"7181fe2e",
          8682 => x"db3887c0",
          8683 => x"98a40851",
          8684 => x"ff557073",
          8685 => x"2780c838",
          8686 => x"715571ff",
          8687 => x"2e80c038",
          8688 => x"87c0989c",
          8689 => x"0880ce90",
          8690 => x"055387c0",
          8691 => x"989c0852",
          8692 => x"87c0989c",
          8693 => x"08557472",
          8694 => x"2ef63881",
          8695 => x"143387c0",
          8696 => x"989c0852",
          8697 => x"52707327",
          8698 => x"87387181",
          8699 => x"ff2edb38",
          8700 => x"87c098a4",
          8701 => x"08557275",
          8702 => x"268338ff",
          8703 => x"527155ff",
          8704 => x"167081ff",
          8705 => x"06575375",
          8706 => x"802ea138",
          8707 => x"7481ff06",
          8708 => x"5271fed5",
          8709 => x"38745170",
          8710 => x"81ff0654",
          8711 => x"73802e83",
          8712 => x"38815776",
          8713 => x"84bb840c",
          8714 => x"883d0d04",
          8715 => x"ff51e839",
          8716 => x"fb3d0d83",
          8717 => x"f5900851",
          8718 => x"80d07134",
          8719 => x"850b83f5",
          8720 => x"90085656",
          8721 => x"fe0b8116",
          8722 => x"34800b87",
          8723 => x"9080e834",
          8724 => x"87c0989c",
          8725 => x"0883f590",
          8726 => x"085680ce",
          8727 => x"90055487",
          8728 => x"c0989c08",
          8729 => x"5287c098",
          8730 => x"9c085372",
          8731 => x"722ef638",
          8732 => x"81153387",
          8733 => x"c0989c08",
          8734 => x"52527074",
          8735 => x"27873871",
          8736 => x"81fe2edb",
          8737 => x"3887c098",
          8738 => x"a40851ff",
          8739 => x"53707427",
          8740 => x"80c83871",
          8741 => x"5371ff2e",
          8742 => x"80c03887",
          8743 => x"c0989c08",
          8744 => x"80ce9005",
          8745 => x"5387c098",
          8746 => x"9c085287",
          8747 => x"c0989c08",
          8748 => x"5170722e",
          8749 => x"f6388115",
          8750 => x"3387c098",
          8751 => x"9c085552",
          8752 => x"73732787",
          8753 => x"387181ff",
          8754 => x"2edb3887",
          8755 => x"c098a408",
          8756 => x"51727126",
          8757 => x"8338ff52",
          8758 => x"7153ff16",
          8759 => x"7081ff06",
          8760 => x"57527580",
          8761 => x"2e8a3872",
          8762 => x"81ff0654",
          8763 => x"73fed538",
          8764 => x"ff39803d",
          8765 => x"0d83e688",
          8766 => x"51fecef7",
          8767 => x"3f823d0d",
          8768 => x"04f93d0d",
          8769 => x"84baf408",
          8770 => x"7a713183",
          8771 => x"2a7083ff",
          8772 => x"ff067083",
          8773 => x"2b731170",
          8774 => x"33811233",
          8775 => x"718b2b71",
          8776 => x"832b0777",
          8777 => x"11703381",
          8778 => x"12337198",
          8779 => x"2b71902b",
          8780 => x"075c5441",
          8781 => x"53535d57",
          8782 => x"59525657",
          8783 => x"53807124",
          8784 => x"81af3872",
          8785 => x"16821133",
          8786 => x"83123371",
          8787 => x"8b2b7183",
          8788 => x"2b077605",
          8789 => x"70338112",
          8790 => x"3371982b",
          8791 => x"71902b07",
          8792 => x"57535c52",
          8793 => x"59565280",
          8794 => x"7124839e",
          8795 => x"38841333",
          8796 => x"85143371",
          8797 => x"8b2b7183",
          8798 => x"2b077505",
          8799 => x"76882a52",
          8800 => x"54565774",
          8801 => x"86133473",
          8802 => x"81ff0654",
          8803 => x"73871334",
          8804 => x"84baf408",
          8805 => x"70178412",
          8806 => x"33851333",
          8807 => x"71882b07",
          8808 => x"70882a5c",
          8809 => x"55595451",
          8810 => x"77841434",
          8811 => x"71851434",
          8812 => x"84baf408",
          8813 => x"1652800b",
          8814 => x"86133480",
          8815 => x"0b871334",
          8816 => x"84baf408",
          8817 => x"53748414",
          8818 => x"34738514",
          8819 => x"3484baf4",
          8820 => x"08167033",
          8821 => x"81123371",
          8822 => x"882b0782",
          8823 => x"80800770",
          8824 => x"882a5858",
          8825 => x"52527472",
          8826 => x"34758113",
          8827 => x"34893d0d",
          8828 => x"04861233",
          8829 => x"87133371",
          8830 => x"8b2b7183",
          8831 => x"2b077511",
          8832 => x"84163385",
          8833 => x"17337188",
          8834 => x"2b077088",
          8835 => x"2a585854",
          8836 => x"51535858",
          8837 => x"71841234",
          8838 => x"72851234",
          8839 => x"84baf408",
          8840 => x"70168411",
          8841 => x"33851233",
          8842 => x"718b2b71",
          8843 => x"832b0756",
          8844 => x"5a5a5272",
          8845 => x"05861233",
          8846 => x"87133371",
          8847 => x"882b0770",
          8848 => x"882a5255",
          8849 => x"59527786",
          8850 => x"13347287",
          8851 => x"133484ba",
          8852 => x"f4081570",
          8853 => x"33811233",
          8854 => x"71882b07",
          8855 => x"81ffff06",
          8856 => x"70882a5a",
          8857 => x"5a545276",
          8858 => x"72347781",
          8859 => x"133484ba",
          8860 => x"f4087017",
          8861 => x"70338112",
          8862 => x"33718b2b",
          8863 => x"71832b07",
          8864 => x"74057033",
          8865 => x"81123371",
          8866 => x"882b0770",
          8867 => x"832b8fff",
          8868 => x"f8067705",
          8869 => x"7b882a54",
          8870 => x"5253545c",
          8871 => x"5a575452",
          8872 => x"77821434",
          8873 => x"73831434",
          8874 => x"84baf408",
          8875 => x"70177033",
          8876 => x"81123371",
          8877 => x"8b2b7183",
          8878 => x"2b077405",
          8879 => x"70338112",
          8880 => x"3371882b",
          8881 => x"0781ffff",
          8882 => x"0670882a",
          8883 => x"5f525355",
          8884 => x"5a575452",
          8885 => x"77733470",
          8886 => x"81143484",
          8887 => x"baf40870",
          8888 => x"17821133",
          8889 => x"83123371",
          8890 => x"8b2b7183",
          8891 => x"2b077405",
          8892 => x"70338112",
          8893 => x"3371982b",
          8894 => x"71902b07",
          8895 => x"58535d52",
          8896 => x"5a575353",
          8897 => x"708025fc",
          8898 => x"e4387133",
          8899 => x"81133371",
          8900 => x"882b0782",
          8901 => x"80800770",
          8902 => x"882a5959",
          8903 => x"54767534",
          8904 => x"77811634",
          8905 => x"84baf408",
          8906 => x"70177033",
          8907 => x"81123371",
          8908 => x"8b2b7183",
          8909 => x"2b077405",
          8910 => x"82143383",
          8911 => x"15337188",
          8912 => x"2b077088",
          8913 => x"2a575c5c",
          8914 => x"52585652",
          8915 => x"53728215",
          8916 => x"34758315",
          8917 => x"34893d0d",
          8918 => x"04f93d0d",
          8919 => x"7984baf4",
          8920 => x"08585876",
          8921 => x"802e8f38",
          8922 => x"77802e86",
          8923 => x"387751fb",
          8924 => x"903f893d",
          8925 => x"0d0484ff",
          8926 => x"f40b84ba",
          8927 => x"f40ca080",
          8928 => x"0b84baf0",
          8929 => x"23828080",
          8930 => x"53765284",
          8931 => x"fff451fe",
          8932 => x"d1ed3f84",
          8933 => x"baf40855",
          8934 => x"76753481",
          8935 => x"0b811634",
          8936 => x"84baf408",
          8937 => x"54768415",
          8938 => x"34810b85",
          8939 => x"153484ba",
          8940 => x"f4085676",
          8941 => x"86173481",
          8942 => x"0b871734",
          8943 => x"84baf408",
          8944 => x"84baf022",
          8945 => x"ff05fe80",
          8946 => x"80077083",
          8947 => x"ffff0670",
          8948 => x"882a5851",
          8949 => x"55567488",
          8950 => x"17347389",
          8951 => x"173484ba",
          8952 => x"f0227010",
          8953 => x"101084ba",
          8954 => x"f40805f8",
          8955 => x"05555576",
          8956 => x"82153481",
          8957 => x"0b831534",
          8958 => x"feee39f7",
          8959 => x"3d0d7b52",
          8960 => x"80538151",
          8961 => x"8472278e",
          8962 => x"38fb1283",
          8963 => x"2a820570",
          8964 => x"83ffff06",
          8965 => x"51517083",
          8966 => x"ffff0684",
          8967 => x"baf40884",
          8968 => x"11338512",
          8969 => x"3371882b",
          8970 => x"07705259",
          8971 => x"5a585581",
          8972 => x"ffff5475",
          8973 => x"802e80cc",
          8974 => x"38751010",
          8975 => x"10177033",
          8976 => x"81123371",
          8977 => x"882b0770",
          8978 => x"81ffff06",
          8979 => x"79317083",
          8980 => x"ffff0670",
          8981 => x"7a275653",
          8982 => x"5c5c5452",
          8983 => x"7274278a",
          8984 => x"3870802e",
          8985 => x"85387573",
          8986 => x"55588412",
          8987 => x"33851333",
          8988 => x"71882b07",
          8989 => x"575a75c1",
          8990 => x"387381ff",
          8991 => x"ff2e8538",
          8992 => x"77745456",
          8993 => x"8076832b",
          8994 => x"78117033",
          8995 => x"81123371",
          8996 => x"882b0770",
          8997 => x"81ffff06",
          8998 => x"56565d56",
          8999 => x"59597079",
          9000 => x"2e833881",
          9001 => x"59805174",
          9002 => x"7326828d",
          9003 => x"38785178",
          9004 => x"802e8285",
          9005 => x"3872752e",
          9006 => x"82883874",
          9007 => x"1670832b",
          9008 => x"78117482",
          9009 => x"80800770",
          9010 => x"882a5b5c",
          9011 => x"56565a76",
          9012 => x"74347881",
          9013 => x"153484ba",
          9014 => x"f4081576",
          9015 => x"882a5353",
          9016 => x"71821434",
          9017 => x"75831434",
          9018 => x"84baf408",
          9019 => x"70197033",
          9020 => x"81123371",
          9021 => x"882b0770",
          9022 => x"832b8fff",
          9023 => x"f8067405",
          9024 => x"7e83ffff",
          9025 => x"0670882a",
          9026 => x"5c585357",
          9027 => x"59525275",
          9028 => x"82123472",
          9029 => x"81ff0653",
          9030 => x"72831234",
          9031 => x"84baf408",
          9032 => x"18547574",
          9033 => x"34728115",
          9034 => x"3484baf4",
          9035 => x"08701986",
          9036 => x"11338712",
          9037 => x"33718b2b",
          9038 => x"71832b07",
          9039 => x"7405585c",
          9040 => x"5c535775",
          9041 => x"84153472",
          9042 => x"85153484",
          9043 => x"baf40870",
          9044 => x"16557805",
          9045 => x"86113387",
          9046 => x"12337188",
          9047 => x"2b077088",
          9048 => x"2a545458",
          9049 => x"59708615",
          9050 => x"34718715",
          9051 => x"3484baf4",
          9052 => x"08701984",
          9053 => x"11338512",
          9054 => x"33718b2b",
          9055 => x"71832b07",
          9056 => x"7405585a",
          9057 => x"5c5a5275",
          9058 => x"86153472",
          9059 => x"87153484",
          9060 => x"baf40870",
          9061 => x"16557805",
          9062 => x"84113385",
          9063 => x"12337188",
          9064 => x"2b077088",
          9065 => x"2a545c57",
          9066 => x"59708415",
          9067 => x"34798515",
          9068 => x"3484baf4",
          9069 => x"08188405",
          9070 => x"517084bb",
          9071 => x"840c8b3d",
          9072 => x"0d048614",
          9073 => x"33871533",
          9074 => x"718b2b71",
          9075 => x"832b0779",
          9076 => x"05841733",
          9077 => x"85183371",
          9078 => x"882b0770",
          9079 => x"882a5a5b",
          9080 => x"59535452",
          9081 => x"74841234",
          9082 => x"76851234",
          9083 => x"84baf408",
          9084 => x"70198411",
          9085 => x"33851233",
          9086 => x"718b2b71",
          9087 => x"832b0774",
          9088 => x"05861433",
          9089 => x"87153371",
          9090 => x"882b0770",
          9091 => x"882a585d",
          9092 => x"5f52565b",
          9093 => x"57527086",
          9094 => x"1a347687",
          9095 => x"1a3484ba",
          9096 => x"f4081870",
          9097 => x"33811233",
          9098 => x"71882b07",
          9099 => x"81ffff06",
          9100 => x"70882a59",
          9101 => x"57545775",
          9102 => x"77347481",
          9103 => x"183484ba",
          9104 => x"f4081884",
          9105 => x"0551fef1",
          9106 => x"39f93d0d",
          9107 => x"7984baf4",
          9108 => x"08585876",
          9109 => x"802ea038",
          9110 => x"7754778a",
          9111 => x"387384bb",
          9112 => x"840c893d",
          9113 => x"0d047751",
          9114 => x"fb913f84",
          9115 => x"bb840884",
          9116 => x"bb840c89",
          9117 => x"3d0d0484",
          9118 => x"fff40b84",
          9119 => x"baf40ca0",
          9120 => x"800b84ba",
          9121 => x"f0238280",
          9122 => x"80537652",
          9123 => x"84fff451",
          9124 => x"fecbec3f",
          9125 => x"84baf408",
          9126 => x"55767534",
          9127 => x"810b8116",
          9128 => x"3484baf4",
          9129 => x"08547684",
          9130 => x"1534810b",
          9131 => x"85153484",
          9132 => x"baf40856",
          9133 => x"76861734",
          9134 => x"810b8717",
          9135 => x"3484baf4",
          9136 => x"0884baf0",
          9137 => x"22ff05fe",
          9138 => x"80800770",
          9139 => x"83ffff06",
          9140 => x"70882a58",
          9141 => x"51555674",
          9142 => x"88173473",
          9143 => x"89173484",
          9144 => x"baf02270",
          9145 => x"10101084",
          9146 => x"baf40805",
          9147 => x"f8055555",
          9148 => x"76821534",
          9149 => x"810b8315",
          9150 => x"34775477",
          9151 => x"802efedd",
          9152 => x"38fee339",
          9153 => x"ed3d0d65",
          9154 => x"67415f80",
          9155 => x"7084baf4",
          9156 => x"08594541",
          9157 => x"76612e84",
          9158 => x"aa387e80",
          9159 => x"2e85af38",
          9160 => x"7f802e88",
          9161 => x"d7388154",
          9162 => x"8460278f",
          9163 => x"387ffb05",
          9164 => x"832a8205",
          9165 => x"7083ffff",
          9166 => x"06555873",
          9167 => x"83ffff06",
          9168 => x"7f783183",
          9169 => x"2a7083ff",
          9170 => x"ff067083",
          9171 => x"2b7a1170",
          9172 => x"33811233",
          9173 => x"71882b07",
          9174 => x"70753170",
          9175 => x"83ffff06",
          9176 => x"70101010",
          9177 => x"fc057383",
          9178 => x"2b611170",
          9179 => x"33811233",
          9180 => x"71882b07",
          9181 => x"70902b70",
          9182 => x"902c5342",
          9183 => x"45464453",
          9184 => x"5443445c",
          9185 => x"4859525e",
          9186 => x"5f42807a",
          9187 => x"2485fd38",
          9188 => x"82153383",
          9189 => x"16337188",
          9190 => x"2b077010",
          9191 => x"10101970",
          9192 => x"33811233",
          9193 => x"71982b71",
          9194 => x"902b0753",
          9195 => x"5c535656",
          9196 => x"56807424",
          9197 => x"85c9387a",
          9198 => x"622782f6",
          9199 => x"38631b58",
          9200 => x"77622e87",
          9201 => x"a2386080",
          9202 => x"2e85f938",
          9203 => x"601b5877",
          9204 => x"622587be",
          9205 => x"38631859",
          9206 => x"61792492",
          9207 => x"f738761e",
          9208 => x"70338112",
          9209 => x"33718b2b",
          9210 => x"71832b07",
          9211 => x"7a117033",
          9212 => x"81123371",
          9213 => x"982b7190",
          9214 => x"2b074743",
          9215 => x"59525357",
          9216 => x"5b588060",
          9217 => x"248cba38",
          9218 => x"761e8211",
          9219 => x"33831233",
          9220 => x"718b2b71",
          9221 => x"832b077a",
          9222 => x"11861133",
          9223 => x"87123371",
          9224 => x"8b2b7183",
          9225 => x"2b077e05",
          9226 => x"84143385",
          9227 => x"15337188",
          9228 => x"2b077088",
          9229 => x"2a595748",
          9230 => x"525b4158",
          9231 => x"535c5956",
          9232 => x"77841d34",
          9233 => x"79851d34",
          9234 => x"84baf408",
          9235 => x"70178411",
          9236 => x"33851233",
          9237 => x"718b2b71",
          9238 => x"832b0774",
          9239 => x"05861433",
          9240 => x"87153371",
          9241 => x"882b0770",
          9242 => x"882a5f42",
          9243 => x"5e524057",
          9244 => x"41577786",
          9245 => x"16347b87",
          9246 => x"163484ba",
          9247 => x"f4081670",
          9248 => x"33811233",
          9249 => x"71882b07",
          9250 => x"81ffff06",
          9251 => x"70882a5a",
          9252 => x"5c5e5976",
          9253 => x"79347981",
          9254 => x"1a3484ba",
          9255 => x"f408701f",
          9256 => x"82113383",
          9257 => x"1233718b",
          9258 => x"2b71832b",
          9259 => x"07740573",
          9260 => x"33811533",
          9261 => x"71882b07",
          9262 => x"70882a41",
          9263 => x"5c455d5f",
          9264 => x"5a555579",
          9265 => x"79347581",
          9266 => x"1a3484ba",
          9267 => x"f408701f",
          9268 => x"70338112",
          9269 => x"33718b2b",
          9270 => x"71832b07",
          9271 => x"74058214",
          9272 => x"33831533",
          9273 => x"71882b07",
          9274 => x"70882a41",
          9275 => x"5c455d5f",
          9276 => x"5a555579",
          9277 => x"821a3475",
          9278 => x"831a3484",
          9279 => x"baf40870",
          9280 => x"1f821133",
          9281 => x"83123371",
          9282 => x"882b0766",
          9283 => x"57625670",
          9284 => x"832b4252",
          9285 => x"5a5d7e05",
          9286 => x"840551fe",
          9287 => x"c3a43f84",
          9288 => x"baf4081e",
          9289 => x"84056165",
          9290 => x"051c7083",
          9291 => x"ffff065d",
          9292 => x"445f7a62",
          9293 => x"2681b638",
          9294 => x"7e547384",
          9295 => x"bb840c95",
          9296 => x"3d0d0484",
          9297 => x"fff40b84",
          9298 => x"baf40ca0",
          9299 => x"800b84ba",
          9300 => x"f0238280",
          9301 => x"80536052",
          9302 => x"84fff451",
          9303 => x"fec6a03f",
          9304 => x"84baf408",
          9305 => x"5e607e34",
          9306 => x"810b811f",
          9307 => x"3484baf4",
          9308 => x"085d6084",
          9309 => x"1e34810b",
          9310 => x"851e3484",
          9311 => x"baf4085c",
          9312 => x"60861d34",
          9313 => x"810b871d",
          9314 => x"3484baf4",
          9315 => x"0884baf0",
          9316 => x"22ff05fe",
          9317 => x"80800770",
          9318 => x"83ffff06",
          9319 => x"70882a5c",
          9320 => x"5a5b5778",
          9321 => x"88183477",
          9322 => x"89183484",
          9323 => x"baf02270",
          9324 => x"10101084",
          9325 => x"baf40805",
          9326 => x"f8055556",
          9327 => x"60821534",
          9328 => x"810b8315",
          9329 => x"3484baf4",
          9330 => x"08577efa",
          9331 => x"d3387680",
          9332 => x"2e828c38",
          9333 => x"7e547f80",
          9334 => x"2efedf38",
          9335 => x"7f51f49b",
          9336 => x"3f84bb84",
          9337 => x"0884bb84",
          9338 => x"0c953d0d",
          9339 => x"04611c84",
          9340 => x"baf40871",
          9341 => x"832b7111",
          9342 => x"5e447f05",
          9343 => x"70338112",
          9344 => x"3371882b",
          9345 => x"0781ffff",
          9346 => x"0670882a",
          9347 => x"48445b5e",
          9348 => x"40637b34",
          9349 => x"60811c34",
          9350 => x"6184baf4",
          9351 => x"08057c88",
          9352 => x"2a575875",
          9353 => x"8219347b",
          9354 => x"83193484",
          9355 => x"baf40870",
          9356 => x"1f703381",
          9357 => x"12337188",
          9358 => x"2b077083",
          9359 => x"2b8ffff8",
          9360 => x"06740564",
          9361 => x"83ffff06",
          9362 => x"70882a4a",
          9363 => x"5c47575e",
          9364 => x"5b5d6363",
          9365 => x"82053476",
          9366 => x"81ff0641",
          9367 => x"60638305",
          9368 => x"3484baf4",
          9369 => x"081e5b63",
          9370 => x"7b346081",
          9371 => x"1c346184",
          9372 => x"baf40805",
          9373 => x"840551ed",
          9374 => x"883f7e54",
          9375 => x"fdbc397b",
          9376 => x"75317083",
          9377 => x"ffff0642",
          9378 => x"54faac39",
          9379 => x"7781ffff",
          9380 => x"06763170",
          9381 => x"83ffff06",
          9382 => x"82173383",
          9383 => x"18337188",
          9384 => x"2b077010",
          9385 => x"10101b70",
          9386 => x"33811233",
          9387 => x"71982b71",
          9388 => x"902b0753",
          9389 => x"5e535458",
          9390 => x"58455473",
          9391 => x"8025f9f7",
          9392 => x"38ffbc39",
          9393 => x"617824fa",
          9394 => x"8338807a",
          9395 => x"248b8f38",
          9396 => x"7783ffff",
          9397 => x"065b617b",
          9398 => x"27fcdd38",
          9399 => x"fe8f3984",
          9400 => x"fff40b84",
          9401 => x"baf40ca0",
          9402 => x"800b84ba",
          9403 => x"f0238280",
          9404 => x"80537e52",
          9405 => x"84fff451",
          9406 => x"fec3843f",
          9407 => x"84baf408",
          9408 => x"5a7e7a34",
          9409 => x"810b811b",
          9410 => x"3484baf4",
          9411 => x"08597e84",
          9412 => x"1a34810b",
          9413 => x"851a3484",
          9414 => x"baf40858",
          9415 => x"7e861934",
          9416 => x"810b8719",
          9417 => x"3484baf4",
          9418 => x"0884baf0",
          9419 => x"22ff05fe",
          9420 => x"80800770",
          9421 => x"83ffff06",
          9422 => x"70882a58",
          9423 => x"56574474",
          9424 => x"64880534",
          9425 => x"73648905",
          9426 => x"3484baf0",
          9427 => x"22701010",
          9428 => x"1084baf4",
          9429 => x"0805f805",
          9430 => x"42437e61",
          9431 => x"82053481",
          9432 => x"61830534",
          9433 => x"fcee3980",
          9434 => x"7a2483de",
          9435 => x"386183ff",
          9436 => x"ff065b61",
          9437 => x"7b27fbc0",
          9438 => x"38fcf239",
          9439 => x"76802e82",
          9440 => x"bd387e51",
          9441 => x"eafb3f7f",
          9442 => x"547384bb",
          9443 => x"840c953d",
          9444 => x"0d04761e",
          9445 => x"82113383",
          9446 => x"1233718b",
          9447 => x"2b71832b",
          9448 => x"077a1186",
          9449 => x"11338712",
          9450 => x"33718b2b",
          9451 => x"71832b07",
          9452 => x"7e058414",
          9453 => x"33851533",
          9454 => x"71882b07",
          9455 => x"70882a43",
          9456 => x"4445565b",
          9457 => x"4658535c",
          9458 => x"45567864",
          9459 => x"8405347a",
          9460 => x"64850534",
          9461 => x"84baf408",
          9462 => x"70178411",
          9463 => x"33851233",
          9464 => x"718b2b71",
          9465 => x"832b0774",
          9466 => x"05861433",
          9467 => x"87153371",
          9468 => x"882b0770",
          9469 => x"882a5b41",
          9470 => x"42485d59",
          9471 => x"5d417364",
          9472 => x"8605347a",
          9473 => x"64870534",
          9474 => x"84baf408",
          9475 => x"16703381",
          9476 => x"12337188",
          9477 => x"2b0781ff",
          9478 => x"ff067088",
          9479 => x"2a5f5c5a",
          9480 => x"5d7b7d34",
          9481 => x"79811e34",
          9482 => x"84baf408",
          9483 => x"701f8211",
          9484 => x"33831233",
          9485 => x"718b2b71",
          9486 => x"832b0774",
          9487 => x"05733381",
          9488 => x"15337188",
          9489 => x"2b077088",
          9490 => x"2a5e5c5e",
          9491 => x"40435745",
          9492 => x"54767c34",
          9493 => x"75811d34",
          9494 => x"84baf408",
          9495 => x"701f7033",
          9496 => x"81123371",
          9497 => x"8b2b7183",
          9498 => x"2b077405",
          9499 => x"82143383",
          9500 => x"15337188",
          9501 => x"2b077088",
          9502 => x"2a404740",
          9503 => x"5b405c55",
          9504 => x"55788218",
          9505 => x"34608318",
          9506 => x"3484baf4",
          9507 => x"08701f82",
          9508 => x"11338312",
          9509 => x"3371882b",
          9510 => x"07665762",
          9511 => x"5670832b",
          9512 => x"4252585d",
          9513 => x"7e058405",
          9514 => x"51febc96",
          9515 => x"3f84baf4",
          9516 => x"081e8405",
          9517 => x"7883ffff",
          9518 => x"065c5ffc",
          9519 => x"993984ff",
          9520 => x"f40b84ba",
          9521 => x"f40ca080",
          9522 => x"0b84baf0",
          9523 => x"23828080",
          9524 => x"537f5284",
          9525 => x"fff451fe",
          9526 => x"bfa53f84",
          9527 => x"baf40856",
          9528 => x"7f763481",
          9529 => x"0b811734",
          9530 => x"84baf408",
          9531 => x"557f8416",
          9532 => x"34810b85",
          9533 => x"163484ba",
          9534 => x"f408547f",
          9535 => x"86153481",
          9536 => x"0b871534",
          9537 => x"84baf408",
          9538 => x"84baf022",
          9539 => x"ff05fe80",
          9540 => x"80077083",
          9541 => x"ffff0670",
          9542 => x"882a4543",
          9543 => x"445e6188",
          9544 => x"1f346089",
          9545 => x"1f3484ba",
          9546 => x"f0227010",
          9547 => x"101084ba",
          9548 => x"f40805f8",
          9549 => x"055c5d7f",
          9550 => x"821c3481",
          9551 => x"0b831c34",
          9552 => x"7e51e7bd",
          9553 => x"3f7f54fc",
          9554 => x"c0398619",
          9555 => x"33871a33",
          9556 => x"718b2b71",
          9557 => x"832b0779",
          9558 => x"05841c33",
          9559 => x"851d3371",
          9560 => x"882b0770",
          9561 => x"882a5c48",
          9562 => x"5e435955",
          9563 => x"76618405",
          9564 => x"34636185",
          9565 => x"053484ba",
          9566 => x"f408701e",
          9567 => x"84113385",
          9568 => x"1233718b",
          9569 => x"2b71832b",
          9570 => x"07740586",
          9571 => x"14338715",
          9572 => x"3371882b",
          9573 => x"0770882a",
          9574 => x"415f4848",
          9575 => x"59565940",
          9576 => x"79648605",
          9577 => x"34786487",
          9578 => x"053484ba",
          9579 => x"f4081d70",
          9580 => x"33811233",
          9581 => x"71882b07",
          9582 => x"81ffff06",
          9583 => x"70882a59",
          9584 => x"42585875",
          9585 => x"78347f81",
          9586 => x"193484ba",
          9587 => x"f408701f",
          9588 => x"70338112",
          9589 => x"33718b2b",
          9590 => x"71832b07",
          9591 => x"74057033",
          9592 => x"81123371",
          9593 => x"882b0770",
          9594 => x"832b8fff",
          9595 => x"f8067705",
          9596 => x"63882a48",
          9597 => x"5d5d5a5d",
          9598 => x"405d4441",
          9599 => x"7f821734",
          9600 => x"7b831734",
          9601 => x"84baf408",
          9602 => x"701f7033",
          9603 => x"81123371",
          9604 => x"8b2b7183",
          9605 => x"2b077405",
          9606 => x"70338112",
          9607 => x"3371882b",
          9608 => x"0781ffff",
          9609 => x"0670882a",
          9610 => x"485d5e5e",
          9611 => x"465a415b",
          9612 => x"60603476",
          9613 => x"60810534",
          9614 => x"6183ffff",
          9615 => x"065bfab3",
          9616 => x"39861533",
          9617 => x"87163371",
          9618 => x"8b2b7183",
          9619 => x"2b077905",
          9620 => x"84183385",
          9621 => x"19337188",
          9622 => x"2b077088",
          9623 => x"2a5e5e5a",
          9624 => x"52415d78",
          9625 => x"841e3479",
          9626 => x"851e3484",
          9627 => x"baf40870",
          9628 => x"19841133",
          9629 => x"85123371",
          9630 => x"8b2b7183",
          9631 => x"2b077405",
          9632 => x"86143387",
          9633 => x"15337188",
          9634 => x"2b077088",
          9635 => x"2a44565e",
          9636 => x"525a4255",
          9637 => x"567c6086",
          9638 => x"05347560",
          9639 => x"87053484",
          9640 => x"baf40818",
          9641 => x"70338112",
          9642 => x"3371882b",
          9643 => x"0781ffff",
          9644 => x"0670882a",
          9645 => x"5b5b5855",
          9646 => x"77753478",
          9647 => x"81163484",
          9648 => x"baf40870",
          9649 => x"1f703381",
          9650 => x"1233718b",
          9651 => x"2b71832b",
          9652 => x"07740570",
          9653 => x"33811233",
          9654 => x"71882b07",
          9655 => x"70832b8f",
          9656 => x"fff80677",
          9657 => x"0563882a",
          9658 => x"56545f5f",
          9659 => x"5859425e",
          9660 => x"557f8217",
          9661 => x"347b8317",
          9662 => x"3484baf4",
          9663 => x"08701f70",
          9664 => x"33811233",
          9665 => x"718b2b71",
          9666 => x"832b0774",
          9667 => x"05703381",
          9668 => x"12337188",
          9669 => x"2b0781ff",
          9670 => x"ff067088",
          9671 => x"2a5d545e",
          9672 => x"585b595d",
          9673 => x"55757c34",
          9674 => x"76811d34",
          9675 => x"84baf408",
          9676 => x"701f8211",
          9677 => x"33831233",
          9678 => x"718b2b71",
          9679 => x"832b0774",
          9680 => x"11861133",
          9681 => x"87123371",
          9682 => x"8b2b7183",
          9683 => x"2b077805",
          9684 => x"84143385",
          9685 => x"15337188",
          9686 => x"2b077088",
          9687 => x"2a595749",
          9688 => x"525c4259",
          9689 => x"535d5a57",
          9690 => x"5777841d",
          9691 => x"3479851d",
          9692 => x"3484baf4",
          9693 => x"08701784",
          9694 => x"11338512",
          9695 => x"33718b2b",
          9696 => x"71832b07",
          9697 => x"74058614",
          9698 => x"33871533",
          9699 => x"71882b07",
          9700 => x"70882a5f",
          9701 => x"425e5240",
          9702 => x"57415777",
          9703 => x"8616347b",
          9704 => x"87163484",
          9705 => x"baf40816",
          9706 => x"70338112",
          9707 => x"3371882b",
          9708 => x"0781ffff",
          9709 => x"0670882a",
          9710 => x"5a5c5e59",
          9711 => x"76793479",
          9712 => x"811a3484",
          9713 => x"baf40870",
          9714 => x"1f821133",
          9715 => x"83123371",
          9716 => x"8b2b7183",
          9717 => x"2b077405",
          9718 => x"73338115",
          9719 => x"3371882b",
          9720 => x"0770882a",
          9721 => x"415c455d",
          9722 => x"5f5a5555",
          9723 => x"79793475",
          9724 => x"811a3484",
          9725 => x"baf40870",
          9726 => x"1f703381",
          9727 => x"1233718b",
          9728 => x"2b71832b",
          9729 => x"07740582",
          9730 => x"14338315",
          9731 => x"3371882b",
          9732 => x"0770882a",
          9733 => x"415c455d",
          9734 => x"5f5a5555",
          9735 => x"79821a34",
          9736 => x"75831a34",
          9737 => x"84baf408",
          9738 => x"701f8211",
          9739 => x"33831233",
          9740 => x"71882b07",
          9741 => x"66576256",
          9742 => x"70832b42",
          9743 => x"525a5d7e",
          9744 => x"05840551",
          9745 => x"feb4fb3f",
          9746 => x"84baf408",
          9747 => x"1e840561",
          9748 => x"65051c70",
          9749 => x"83ffff06",
          9750 => x"5d445ff1",
          9751 => x"d5398619",
          9752 => x"33871a33",
          9753 => x"718b2b71",
          9754 => x"832b0779",
          9755 => x"05841c33",
          9756 => x"851d3371",
          9757 => x"882b0770",
          9758 => x"882a4048",
          9759 => x"5d434155",
          9760 => x"7a618405",
          9761 => x"34636185",
          9762 => x"053484ba",
          9763 => x"f408701e",
          9764 => x"84113385",
          9765 => x"1233718b",
          9766 => x"2b71832b",
          9767 => x"07740586",
          9768 => x"14338715",
          9769 => x"3371882b",
          9770 => x"0770882a",
          9771 => x"5b415f48",
          9772 => x"5c594156",
          9773 => x"73648605",
          9774 => x"347a6487",
          9775 => x"053484ba",
          9776 => x"f4081d70",
          9777 => x"33811233",
          9778 => x"71882b07",
          9779 => x"81ffff06",
          9780 => x"70882a5c",
          9781 => x"5f425578",
          9782 => x"75347c81",
          9783 => x"163484ba",
          9784 => x"f408701f",
          9785 => x"70338112",
          9786 => x"33718b2b",
          9787 => x"71832b07",
          9788 => x"74057033",
          9789 => x"81123371",
          9790 => x"882b0770",
          9791 => x"832b8fff",
          9792 => x"f8067705",
          9793 => x"63882a5d",
          9794 => x"445c4958",
          9795 => x"5e455840",
          9796 => x"74821e34",
          9797 => x"7b831e34",
          9798 => x"84baf408",
          9799 => x"701f7033",
          9800 => x"81123371",
          9801 => x"8b2b7183",
          9802 => x"2b077405",
          9803 => x"70338112",
          9804 => x"3371882b",
          9805 => x"0781ffff",
          9806 => x"0670882a",
          9807 => x"475f4958",
          9808 => x"46595e5b",
          9809 => x"7f7d3478",
          9810 => x"811e3477",
          9811 => x"83ffff06",
          9812 => x"5bf38339",
          9813 => x"7e605254",
          9814 => x"e5a13f84",
          9815 => x"bb84085f",
          9816 => x"84bb8408",
          9817 => x"802e9338",
          9818 => x"62537352",
          9819 => x"84bb8408",
          9820 => x"51feb3f6",
          9821 => x"3f7351df",
          9822 => x"883f615b",
          9823 => x"617b27ef",
          9824 => x"b738f0e9",
          9825 => x"39f93d0d",
          9826 => x"7a7a2984",
          9827 => x"baf40858",
          9828 => x"5876802e",
          9829 => x"b7387754",
          9830 => x"778a3873",
          9831 => x"84bb840c",
          9832 => x"893d0d04",
          9833 => x"7751e4d3",
          9834 => x"3f84bb84",
          9835 => x"085484bb",
          9836 => x"8408802e",
          9837 => x"e6387753",
          9838 => x"805284bb",
          9839 => x"840851fe",
          9840 => x"b5bd3f73",
          9841 => x"84bb840c",
          9842 => x"893d0d04",
          9843 => x"84fff40b",
          9844 => x"84baf40c",
          9845 => x"a0800b84",
          9846 => x"baf02382",
          9847 => x"80805376",
          9848 => x"5284fff4",
          9849 => x"51feb597",
          9850 => x"3f84baf4",
          9851 => x"08557675",
          9852 => x"34810b81",
          9853 => x"163484ba",
          9854 => x"f4085476",
          9855 => x"84153481",
          9856 => x"0b851534",
          9857 => x"84baf408",
          9858 => x"56768617",
          9859 => x"34810b87",
          9860 => x"173484ba",
          9861 => x"f40884ba",
          9862 => x"f022ff05",
          9863 => x"fe808007",
          9864 => x"7083ffff",
          9865 => x"0670882a",
          9866 => x"58515556",
          9867 => x"74881734",
          9868 => x"73891734",
          9869 => x"84baf022",
          9870 => x"70101010",
          9871 => x"84baf408",
          9872 => x"05f80555",
          9873 => x"55768215",
          9874 => x"34810b83",
          9875 => x"15347754",
          9876 => x"77802efe",
          9877 => x"c638fecc",
          9878 => x"39ff3d0d",
          9879 => x"028f0533",
          9880 => x"51815270",
          9881 => x"72268738",
          9882 => x"84bb8011",
          9883 => x"33527184",
          9884 => x"bb840c83",
          9885 => x"3d0d04fe",
          9886 => x"3d0d0293",
          9887 => x"05335283",
          9888 => x"53718126",
          9889 => x"9d387151",
          9890 => x"d4bb3f84",
          9891 => x"bb840881",
          9892 => x"ff065372",
          9893 => x"87387284",
          9894 => x"bb801334",
          9895 => x"84bb8012",
          9896 => x"33537284",
          9897 => x"bb840c84",
          9898 => x"3d0d04f7",
          9899 => x"3d0d7c7e",
          9900 => x"60028c05",
          9901 => x"af05335a",
          9902 => x"5c575981",
          9903 => x"54767426",
          9904 => x"873884bb",
          9905 => x"80173354",
          9906 => x"73810654",
          9907 => x"835573bd",
          9908 => x"38735885",
          9909 => x"0b87c098",
          9910 => x"8c0c7853",
          9911 => x"75527651",
          9912 => x"d5ca3f84",
          9913 => x"bb840881",
          9914 => x"ff065574",
          9915 => x"802ea738",
          9916 => x"87c0988c",
          9917 => x"085473e2",
          9918 => x"38797826",
          9919 => x"d63874fc",
          9920 => x"80800654",
          9921 => x"73802e83",
          9922 => x"38815473",
          9923 => x"557484bb",
          9924 => x"840c8b3d",
          9925 => x"0d048480",
          9926 => x"16811970",
          9927 => x"81ff065a",
          9928 => x"55567978",
          9929 => x"26ffac38",
          9930 => x"d539f73d",
          9931 => x"0d7c7e60",
          9932 => x"028c05af",
          9933 => x"05335a5c",
          9934 => x"57598154",
          9935 => x"76742687",
          9936 => x"3884bb80",
          9937 => x"17335473",
          9938 => x"81065483",
          9939 => x"5573bd38",
          9940 => x"7358850b",
          9941 => x"87c0988c",
          9942 => x"0c785375",
          9943 => x"527651d7",
          9944 => x"8e3f84bb",
          9945 => x"840881ff",
          9946 => x"06557480",
          9947 => x"2ea73887",
          9948 => x"c0988c08",
          9949 => x"5473e238",
          9950 => x"797826d6",
          9951 => x"3874fc80",
          9952 => x"80065473",
          9953 => x"802e8338",
          9954 => x"81547355",
          9955 => x"7484bb84",
          9956 => x"0c8b3d0d",
          9957 => x"04848016",
          9958 => x"81197081",
          9959 => x"ff065a55",
          9960 => x"56797826",
          9961 => x"ffac38d5",
          9962 => x"39fc3d0d",
          9963 => x"78028405",
          9964 => x"9b053302",
          9965 => x"88059f05",
          9966 => x"33535355",
          9967 => x"81537173",
          9968 => x"26873884",
          9969 => x"bb801233",
          9970 => x"53728106",
          9971 => x"54835373",
          9972 => x"9b38850b",
          9973 => x"87c0988c",
          9974 => x"0c815370",
          9975 => x"732e9638",
          9976 => x"727125ad",
          9977 => x"3870832e",
          9978 => x"9a388453",
          9979 => x"7284bb84",
          9980 => x"0c863d0d",
          9981 => x"0488800a",
          9982 => x"750c7384",
          9983 => x"bb840c86",
          9984 => x"3d0d0481",
          9985 => x"80750c80",
          9986 => x"0b84bb84",
          9987 => x"0c863d0d",
          9988 => x"0471842b",
          9989 => x"87c0928c",
          9990 => x"11535470",
          9991 => x"cd387108",
          9992 => x"70812a81",
          9993 => x"06515170",
          9994 => x"802e8a38",
          9995 => x"87c0988c",
          9996 => x"085574ea",
          9997 => x"3887c098",
          9998 => x"8c085170",
          9999 => x"ca388172",
         10000 => x"0c87c092",
         10001 => x"8c145271",
         10002 => x"08820654",
         10003 => x"73802eff",
         10004 => x"9b387108",
         10005 => x"82065473",
         10006 => x"ee38ff90",
         10007 => x"39f63d0d",
         10008 => x"7c58800b",
         10009 => x"83193371",
         10010 => x"5b565774",
         10011 => x"772e0981",
         10012 => x"06a83877",
         10013 => x"33567583",
         10014 => x"2e818738",
         10015 => x"80538052",
         10016 => x"81183351",
         10017 => x"fea33f84",
         10018 => x"bb840880",
         10019 => x"2e833881",
         10020 => x"597884bb",
         10021 => x"840c8c3d",
         10022 => x"0d048154",
         10023 => x"b4180853",
         10024 => x"b8187053",
         10025 => x"81193352",
         10026 => x"5afcff3f",
         10027 => x"815984bb",
         10028 => x"8408772e",
         10029 => x"098106d9",
         10030 => x"3884bb84",
         10031 => x"08831934",
         10032 => x"b4180870",
         10033 => x"a81a0831",
         10034 => x"a01a0884",
         10035 => x"bb84085c",
         10036 => x"58565b74",
         10037 => x"7627ff9b",
         10038 => x"38821833",
         10039 => x"5574822e",
         10040 => x"098106ff",
         10041 => x"8e388154",
         10042 => x"751b5379",
         10043 => x"52811833",
         10044 => x"51fcb73f",
         10045 => x"76783357",
         10046 => x"5975832e",
         10047 => x"098106fe",
         10048 => x"fb388418",
         10049 => x"33577681",
         10050 => x"2e098106",
         10051 => x"feee38b8",
         10052 => x"185a8480",
         10053 => x"7a565780",
         10054 => x"75708105",
         10055 => x"5734ff17",
         10056 => x"5776f438",
         10057 => x"80d50b84",
         10058 => x"b61934ff",
         10059 => x"aa0b84b7",
         10060 => x"193480d2",
         10061 => x"7a3480d2",
         10062 => x"0bb91934",
         10063 => x"80e10bba",
         10064 => x"193480c1",
         10065 => x"0bbb1934",
         10066 => x"80f20b84",
         10067 => x"9c193480",
         10068 => x"f20b849d",
         10069 => x"193480c1",
         10070 => x"0b849e19",
         10071 => x"3480e10b",
         10072 => x"849f1934",
         10073 => x"94180855",
         10074 => x"7484a019",
         10075 => x"3474882a",
         10076 => x"5b7a84a1",
         10077 => x"19347490",
         10078 => x"2a567584",
         10079 => x"a2193474",
         10080 => x"982a5b7a",
         10081 => x"84a31934",
         10082 => x"9018085b",
         10083 => x"7a84a419",
         10084 => x"347a882a",
         10085 => x"557484a5",
         10086 => x"19347a90",
         10087 => x"2a567584",
         10088 => x"a619347a",
         10089 => x"982a5574",
         10090 => x"84a71934",
         10091 => x"a4180881",
         10092 => x"0570b41a",
         10093 => x"0c5b8154",
         10094 => x"7a537952",
         10095 => x"81183351",
         10096 => x"fae83f76",
         10097 => x"84193480",
         10098 => x"53805281",
         10099 => x"183351fb",
         10100 => x"d83f84bb",
         10101 => x"8408802e",
         10102 => x"fdb738fd",
         10103 => x"b239f33d",
         10104 => x"0d606070",
         10105 => x"08595656",
         10106 => x"81762788",
         10107 => x"389c1708",
         10108 => x"76268c38",
         10109 => x"81587784",
         10110 => x"bb840c8f",
         10111 => x"3d0d04ff",
         10112 => x"77335658",
         10113 => x"74822e81",
         10114 => x"cc387482",
         10115 => x"2482a538",
         10116 => x"74812e09",
         10117 => x"8106dd38",
         10118 => x"75812a16",
         10119 => x"70892aa8",
         10120 => x"1908055a",
         10121 => x"5a805bb4",
         10122 => x"1708792e",
         10123 => x"b0388317",
         10124 => x"335c7b7b",
         10125 => x"2e098106",
         10126 => x"83de3881",
         10127 => x"547853b8",
         10128 => x"17528117",
         10129 => x"3351f8e3",
         10130 => x"3f84bb84",
         10131 => x"08802e85",
         10132 => x"38ff5981",
         10133 => x"5b78b418",
         10134 => x"0c7aff9a",
         10135 => x"387983ff",
         10136 => x"0617b811",
         10137 => x"33811c70",
         10138 => x"892aa81b",
         10139 => x"0805535d",
         10140 => x"5d59b417",
         10141 => x"08792eb5",
         10142 => x"38800b83",
         10143 => x"1833715c",
         10144 => x"565d747d",
         10145 => x"2e098106",
         10146 => x"84b53881",
         10147 => x"547853b8",
         10148 => x"17528117",
         10149 => x"3351f893",
         10150 => x"3f84bb84",
         10151 => x"08802e85",
         10152 => x"38ff5981",
         10153 => x"5a78b418",
         10154 => x"0c79feca",
         10155 => x"387a83ff",
         10156 => x"0617b811",
         10157 => x"3370882b",
         10158 => x"7e077881",
         10159 => x"0671842a",
         10160 => x"535d5959",
         10161 => x"5d79feae",
         10162 => x"38769fff",
         10163 => x"0684bb84",
         10164 => x"0c8f3d0d",
         10165 => x"0475882a",
         10166 => x"a8180805",
         10167 => x"59b41708",
         10168 => x"792eb538",
         10169 => x"800b8318",
         10170 => x"33715c5d",
         10171 => x"5b7b7b2e",
         10172 => x"09810681",
         10173 => x"c2388154",
         10174 => x"7853b817",
         10175 => x"52811733",
         10176 => x"51f7a83f",
         10177 => x"84bb8408",
         10178 => x"802e8538",
         10179 => x"ff59815a",
         10180 => x"78b4180c",
         10181 => x"79fddf38",
         10182 => x"751083fe",
         10183 => x"067705b8",
         10184 => x"05811133",
         10185 => x"71337188",
         10186 => x"2b0784bb",
         10187 => x"840c575b",
         10188 => x"8f3d0d04",
         10189 => x"74832e09",
         10190 => x"8106fdb8",
         10191 => x"3875872a",
         10192 => x"a8180805",
         10193 => x"59b41708",
         10194 => x"792eb538",
         10195 => x"800b8318",
         10196 => x"33715c5e",
         10197 => x"5b7c7b2e",
         10198 => x"09810682",
         10199 => x"81388154",
         10200 => x"7853b817",
         10201 => x"52811733",
         10202 => x"51f6c03f",
         10203 => x"84bb8408",
         10204 => x"802e8538",
         10205 => x"ff59815a",
         10206 => x"78b4180c",
         10207 => x"79fcf738",
         10208 => x"75822b83",
         10209 => x"fc067705",
         10210 => x"b8058311",
         10211 => x"33821233",
         10212 => x"71902b71",
         10213 => x"882b0781",
         10214 => x"14337072",
         10215 => x"07882b75",
         10216 => x"337180ff",
         10217 => x"fffe8006",
         10218 => x"0784bb84",
         10219 => x"0c415c5e",
         10220 => x"595a568f",
         10221 => x"3d0d0481",
         10222 => x"54b41708",
         10223 => x"53b81770",
         10224 => x"53811833",
         10225 => x"525cf6e2",
         10226 => x"3f815a84",
         10227 => x"bb84087b",
         10228 => x"2e098106",
         10229 => x"febe3884",
         10230 => x"bb840883",
         10231 => x"1834b417",
         10232 => x"08a81808",
         10233 => x"3184bb84",
         10234 => x"085b5e7d",
         10235 => x"a0180827",
         10236 => x"fe843882",
         10237 => x"17335574",
         10238 => x"822e0981",
         10239 => x"06fdf738",
         10240 => x"8154b417",
         10241 => x"08a01808",
         10242 => x"05537b52",
         10243 => x"81173351",
         10244 => x"f6983f7a",
         10245 => x"5afddf39",
         10246 => x"8154b417",
         10247 => x"0853b817",
         10248 => x"70538118",
         10249 => x"33525cf6",
         10250 => x"813f84bb",
         10251 => x"84087b2e",
         10252 => x"09810682",
         10253 => x"813884bb",
         10254 => x"84088318",
         10255 => x"34b41708",
         10256 => x"a8180831",
         10257 => x"5d7ca018",
         10258 => x"08278b38",
         10259 => x"8217335e",
         10260 => x"7d822e81",
         10261 => x"cb3884bb",
         10262 => x"84085bfb",
         10263 => x"de398154",
         10264 => x"b4170853",
         10265 => x"b8177053",
         10266 => x"81183352",
         10267 => x"5cf5bb3f",
         10268 => x"815a84bb",
         10269 => x"84087b2e",
         10270 => x"098106fd",
         10271 => x"ff3884bb",
         10272 => x"84088318",
         10273 => x"34b41708",
         10274 => x"a8180831",
         10275 => x"84bb8408",
         10276 => x"5b5e7da0",
         10277 => x"180827fd",
         10278 => x"c5388217",
         10279 => x"33557482",
         10280 => x"2e098106",
         10281 => x"fdb83881",
         10282 => x"54b41708",
         10283 => x"a0180805",
         10284 => x"537b5281",
         10285 => x"173351f4",
         10286 => x"f13f7a5a",
         10287 => x"fda03981",
         10288 => x"54b41708",
         10289 => x"53b81770",
         10290 => x"53811833",
         10291 => x"525ef4da",
         10292 => x"3f815a84",
         10293 => x"bb84087d",
         10294 => x"2e098106",
         10295 => x"fbcb3884",
         10296 => x"bb840883",
         10297 => x"1834b417",
         10298 => x"08a81808",
         10299 => x"3184bb84",
         10300 => x"085b5574",
         10301 => x"a0180827",
         10302 => x"fb913882",
         10303 => x"17335574",
         10304 => x"822e0981",
         10305 => x"06fb8438",
         10306 => x"8154b417",
         10307 => x"08a01808",
         10308 => x"05537d52",
         10309 => x"81173351",
         10310 => x"f4903f7c",
         10311 => x"5afaec39",
         10312 => x"8154b417",
         10313 => x"08a01808",
         10314 => x"05537b52",
         10315 => x"81173351",
         10316 => x"f3f83ffa",
         10317 => x"8639815b",
         10318 => x"7af9bb38",
         10319 => x"fa9f39f2",
         10320 => x"3d0d6062",
         10321 => x"645d5759",
         10322 => x"82588176",
         10323 => x"279c3875",
         10324 => x"9c1a0827",
         10325 => x"95387833",
         10326 => x"5574782e",
         10327 => x"96387478",
         10328 => x"24818038",
         10329 => x"74812e82",
         10330 => x"8a387784",
         10331 => x"bb840c90",
         10332 => x"3d0d0475",
         10333 => x"882aa81a",
         10334 => x"08055880",
         10335 => x"0bb41a08",
         10336 => x"585c7678",
         10337 => x"2e86b638",
         10338 => x"8319337c",
         10339 => x"5b5d7c7c",
         10340 => x"2e098106",
         10341 => x"83fa3881",
         10342 => x"547753b8",
         10343 => x"19528119",
         10344 => x"3351f287",
         10345 => x"3f84bb84",
         10346 => x"08802e85",
         10347 => x"38ff5881",
         10348 => x"5a77b41a",
         10349 => x"0c795879",
         10350 => x"ffb03875",
         10351 => x"1083fe06",
         10352 => x"79057b83",
         10353 => x"ffff0658",
         10354 => x"5e76b81f",
         10355 => x"3476882a",
         10356 => x"5a79b91f",
         10357 => x"34810b83",
         10358 => x"1a347784",
         10359 => x"bb840c90",
         10360 => x"3d0d0474",
         10361 => x"832e0981",
         10362 => x"06feff38",
         10363 => x"75872aa8",
         10364 => x"1a080558",
         10365 => x"800bb41a",
         10366 => x"08585c76",
         10367 => x"782e85e1",
         10368 => x"38831933",
         10369 => x"7c5b5d7c",
         10370 => x"7c2e0981",
         10371 => x"0684bd38",
         10372 => x"81547753",
         10373 => x"b8195281",
         10374 => x"193351f1",
         10375 => x"8e3f84bb",
         10376 => x"8408802e",
         10377 => x"8538ff58",
         10378 => x"815a77b4",
         10379 => x"1a0c7958",
         10380 => x"79feb738",
         10381 => x"75822b83",
         10382 => x"fc067905",
         10383 => x"b8118311",
         10384 => x"3370982b",
         10385 => x"8f0a067e",
         10386 => x"f00a0607",
         10387 => x"41575e5c",
         10388 => x"7d7d347d",
         10389 => x"882a5675",
         10390 => x"b91d347d",
         10391 => x"902a5a79",
         10392 => x"ba1d347d",
         10393 => x"982a5b7a",
         10394 => x"bb1d3481",
         10395 => x"0b831a34",
         10396 => x"fee83975",
         10397 => x"812a1670",
         10398 => x"892aa81b",
         10399 => x"0805b41b",
         10400 => x"0859595a",
         10401 => x"76782eb7",
         10402 => x"38800b83",
         10403 => x"1a33715e",
         10404 => x"565d747d",
         10405 => x"2e098106",
         10406 => x"82d43881",
         10407 => x"547753b8",
         10408 => x"19528119",
         10409 => x"3351f083",
         10410 => x"3f84bb84",
         10411 => x"08802e85",
         10412 => x"38ff5881",
         10413 => x"5c77b41a",
         10414 => x"0c7b587b",
         10415 => x"fdac3879",
         10416 => x"83ff0619",
         10417 => x"b805811b",
         10418 => x"7781065f",
         10419 => x"5f577a55",
         10420 => x"7c802e8f",
         10421 => x"387a842b",
         10422 => x"9ff00677",
         10423 => x"338f0671",
         10424 => x"07565a74",
         10425 => x"7734810b",
         10426 => x"831a347d",
         10427 => x"892aa81a",
         10428 => x"08055680",
         10429 => x"0bb41a08",
         10430 => x"565f7476",
         10431 => x"2e83dd38",
         10432 => x"81547453",
         10433 => x"b8197053",
         10434 => x"811a3352",
         10435 => x"57f09b3f",
         10436 => x"815884bb",
         10437 => x"84087f2e",
         10438 => x"09810680",
         10439 => x"c73884bb",
         10440 => x"8408831a",
         10441 => x"34b41908",
         10442 => x"70a81b08",
         10443 => x"31a01b08",
         10444 => x"84bb8408",
         10445 => x"5b5c565c",
         10446 => x"747a278b",
         10447 => x"38821933",
         10448 => x"5574822e",
         10449 => x"82e43881",
         10450 => x"54755376",
         10451 => x"52811933",
         10452 => x"51eed83f",
         10453 => x"84bb8408",
         10454 => x"802e8538",
         10455 => x"ff568158",
         10456 => x"75b41a0c",
         10457 => x"77fc8338",
         10458 => x"7d83ff06",
         10459 => x"19b8057b",
         10460 => x"842a5656",
         10461 => x"7c8f387a",
         10462 => x"882a7633",
         10463 => x"81f00671",
         10464 => x"8f060756",
         10465 => x"5c747634",
         10466 => x"810b831a",
         10467 => x"34fccb39",
         10468 => x"81547653",
         10469 => x"b8197053",
         10470 => x"811a3352",
         10471 => x"5def8b3f",
         10472 => x"815a84bb",
         10473 => x"84087c2e",
         10474 => x"098106fc",
         10475 => x"883884bb",
         10476 => x"8408831a",
         10477 => x"34b41908",
         10478 => x"70a81b08",
         10479 => x"31a01b08",
         10480 => x"84bb8408",
         10481 => x"5d59405e",
         10482 => x"7e7727fb",
         10483 => x"ca388219",
         10484 => x"33557482",
         10485 => x"2e098106",
         10486 => x"fbbd3881",
         10487 => x"54761e53",
         10488 => x"7c528119",
         10489 => x"3351eec2",
         10490 => x"3f7b5afb",
         10491 => x"aa398154",
         10492 => x"7653b819",
         10493 => x"7053811a",
         10494 => x"335257ee",
         10495 => x"ad3f815c",
         10496 => x"84bb8408",
         10497 => x"7d2e0981",
         10498 => x"06fdae38",
         10499 => x"84bb8408",
         10500 => x"831a34b4",
         10501 => x"190870a8",
         10502 => x"1b0831a0",
         10503 => x"1b0884bb",
         10504 => x"84085f40",
         10505 => x"565f747e",
         10506 => x"27fcf038",
         10507 => x"82193355",
         10508 => x"74822e09",
         10509 => x"8106fce3",
         10510 => x"3881547d",
         10511 => x"1f537652",
         10512 => x"81193351",
         10513 => x"ede43f7c",
         10514 => x"5cfcd039",
         10515 => x"81547653",
         10516 => x"b8197053",
         10517 => x"811a3352",
         10518 => x"57edcf3f",
         10519 => x"815a84bb",
         10520 => x"84087c2e",
         10521 => x"098106fb",
         10522 => x"c53884bb",
         10523 => x"8408831a",
         10524 => x"34b41908",
         10525 => x"70a81b08",
         10526 => x"31a01b08",
         10527 => x"84bb8408",
         10528 => x"5d5f405e",
         10529 => x"7e7d27fb",
         10530 => x"87388219",
         10531 => x"33557482",
         10532 => x"2e098106",
         10533 => x"fafa3881",
         10534 => x"547c1e53",
         10535 => x"76528119",
         10536 => x"3351ed86",
         10537 => x"3f7b5afa",
         10538 => x"e7398154",
         10539 => x"791c5376",
         10540 => x"52811933",
         10541 => x"51ecf33f",
         10542 => x"7e58fd8b",
         10543 => x"397b7610",
         10544 => x"83fe067a",
         10545 => x"057c83ff",
         10546 => x"ff06595f",
         10547 => x"5876b81f",
         10548 => x"3476882a",
         10549 => x"5a79b91f",
         10550 => x"34f9fa39",
         10551 => x"7e58fd88",
         10552 => x"397b7682",
         10553 => x"2b83fc06",
         10554 => x"7a05b811",
         10555 => x"83113370",
         10556 => x"982b8f0a",
         10557 => x"067ff00a",
         10558 => x"06074258",
         10559 => x"5f5d587d",
         10560 => x"7d347d88",
         10561 => x"2a5675b9",
         10562 => x"1d347d90",
         10563 => x"2a5a79ba",
         10564 => x"1d347d98",
         10565 => x"2a5b7abb",
         10566 => x"1d34facf",
         10567 => x"39f63d0d",
         10568 => x"7c7e7108",
         10569 => x"5b5c5a7a",
         10570 => x"818a3890",
         10571 => x"19085776",
         10572 => x"802e80f4",
         10573 => x"38769c1a",
         10574 => x"082780ec",
         10575 => x"38941908",
         10576 => x"70565473",
         10577 => x"802e80d7",
         10578 => x"38767b2e",
         10579 => x"81933876",
         10580 => x"56811656",
         10581 => x"9c190876",
         10582 => x"26893882",
         10583 => x"56757726",
         10584 => x"82b23875",
         10585 => x"527951f0",
         10586 => x"f53f84bb",
         10587 => x"8408802e",
         10588 => x"81d03880",
         10589 => x"5884bb84",
         10590 => x"08812eb1",
         10591 => x"3884bb84",
         10592 => x"08097030",
         10593 => x"70720780",
         10594 => x"25707b07",
         10595 => x"51515555",
         10596 => x"7382aa38",
         10597 => x"75772e09",
         10598 => x"8106ffb5",
         10599 => x"38735574",
         10600 => x"84bb840c",
         10601 => x"8c3d0d04",
         10602 => x"8157ff91",
         10603 => x"3984bb84",
         10604 => x"0858ca39",
         10605 => x"7a527951",
         10606 => x"f0a43f81",
         10607 => x"557484bb",
         10608 => x"840827db",
         10609 => x"3884bb84",
         10610 => x"085584bb",
         10611 => x"8408ff2e",
         10612 => x"ce389c19",
         10613 => x"0884bb84",
         10614 => x"0826c438",
         10615 => x"7a57fedd",
         10616 => x"39811b56",
         10617 => x"9c190876",
         10618 => x"26833882",
         10619 => x"56755279",
         10620 => x"51efeb3f",
         10621 => x"805884bb",
         10622 => x"8408812e",
         10623 => x"81a03884",
         10624 => x"bb840809",
         10625 => x"70307072",
         10626 => x"07802570",
         10627 => x"7b0784bb",
         10628 => x"84085451",
         10629 => x"51555573",
         10630 => x"ff853884",
         10631 => x"bb840880",
         10632 => x"2e9a3890",
         10633 => x"19085481",
         10634 => x"7427fea3",
         10635 => x"38739c1a",
         10636 => x"0827fe9b",
         10637 => x"38737057",
         10638 => x"57fe9639",
         10639 => x"75802efe",
         10640 => x"8e38ff53",
         10641 => x"75527851",
         10642 => x"f5f53f84",
         10643 => x"bb840884",
         10644 => x"bb840830",
         10645 => x"7084bb84",
         10646 => x"08078025",
         10647 => x"5658557a",
         10648 => x"80c43874",
         10649 => x"80e33875",
         10650 => x"901a0c9c",
         10651 => x"1908fe05",
         10652 => x"941a0856",
         10653 => x"58747826",
         10654 => x"8638ff15",
         10655 => x"941a0c84",
         10656 => x"19338107",
         10657 => x"5a79841a",
         10658 => x"34755574",
         10659 => x"84bb840c",
         10660 => x"8c3d0d04",
         10661 => x"800b84bb",
         10662 => x"840c8c3d",
         10663 => x"0d0484bb",
         10664 => x"840858fe",
         10665 => x"da397380",
         10666 => x"2effb838",
         10667 => x"75537a52",
         10668 => x"7851f58b",
         10669 => x"3f84bb84",
         10670 => x"0855ffa7",
         10671 => x"3984bb84",
         10672 => x"0884bb84",
         10673 => x"0c8c3d0d",
         10674 => x"04ff5674",
         10675 => x"812effb9",
         10676 => x"388155ff",
         10677 => x"b639f83d",
         10678 => x"0d7a7c71",
         10679 => x"08595558",
         10680 => x"73f0800a",
         10681 => x"2680df38",
         10682 => x"739f0653",
         10683 => x"7280d738",
         10684 => x"7390190c",
         10685 => x"88180855",
         10686 => x"7480df38",
         10687 => x"76335675",
         10688 => x"822680cc",
         10689 => x"3873852a",
         10690 => x"53820b88",
         10691 => x"18225a56",
         10692 => x"727927a9",
         10693 => x"38ac1708",
         10694 => x"98190c74",
         10695 => x"94190c98",
         10696 => x"18085382",
         10697 => x"5672802e",
         10698 => x"94387389",
         10699 => x"2a139819",
         10700 => x"0c7383ff",
         10701 => x"0617b805",
         10702 => x"9c190c80",
         10703 => x"567584bb",
         10704 => x"840c8a3d",
         10705 => x"0d04820b",
         10706 => x"84bb840c",
         10707 => x"8a3d0d04",
         10708 => x"ac170855",
         10709 => x"74802eff",
         10710 => x"ac388a17",
         10711 => x"2270892b",
         10712 => x"57597376",
         10713 => x"27a5389c",
         10714 => x"170853fe",
         10715 => x"15fe1454",
         10716 => x"56805975",
         10717 => x"73278d38",
         10718 => x"8a172276",
         10719 => x"7129b019",
         10720 => x"08055a53",
         10721 => x"7898190c",
         10722 => x"ff913974",
         10723 => x"527751ec",
         10724 => x"cd3f84bb",
         10725 => x"84085584",
         10726 => x"bb8408ff",
         10727 => x"2ea43881",
         10728 => x"0b84bb84",
         10729 => x"0827ff9e",
         10730 => x"389c1708",
         10731 => x"5384bb84",
         10732 => x"087327ff",
         10733 => x"91387376",
         10734 => x"31547376",
         10735 => x"27cd38ff",
         10736 => x"aa39810b",
         10737 => x"84bb840c",
         10738 => x"8a3d0d04",
         10739 => x"f33d0d7f",
         10740 => x"70089012",
         10741 => x"08a0055c",
         10742 => x"5a57f080",
         10743 => x"0a7a2786",
         10744 => x"38800b98",
         10745 => x"180c9817",
         10746 => x"08558456",
         10747 => x"74802eb2",
         10748 => x"387983ff",
         10749 => x"065b7a9d",
         10750 => x"38811594",
         10751 => x"18085758",
         10752 => x"75a93879",
         10753 => x"852a881a",
         10754 => x"22575574",
         10755 => x"762781f5",
         10756 => x"38779818",
         10757 => x"0c799018",
         10758 => x"0c781bb8",
         10759 => x"059c180c",
         10760 => x"80567584",
         10761 => x"bb840c8f",
         10762 => x"3d0d0477",
         10763 => x"98180c8a",
         10764 => x"1922ff05",
         10765 => x"7a892a06",
         10766 => x"5c7bda38",
         10767 => x"75527651",
         10768 => x"eb9c3f84",
         10769 => x"bb84085d",
         10770 => x"8256810b",
         10771 => x"84bb8408",
         10772 => x"27d03881",
         10773 => x"5684bb84",
         10774 => x"08ff2ec6",
         10775 => x"389c1908",
         10776 => x"84bb8408",
         10777 => x"26829138",
         10778 => x"60802e81",
         10779 => x"98389417",
         10780 => x"08527651",
         10781 => x"f9a73f84",
         10782 => x"bb84085d",
         10783 => x"875684bb",
         10784 => x"8408802e",
         10785 => x"ff9c3882",
         10786 => x"5684bb84",
         10787 => x"08812eff",
         10788 => x"91388156",
         10789 => x"84bb8408",
         10790 => x"ff2eff86",
         10791 => x"3884bb84",
         10792 => x"08831a33",
         10793 => x"5f587d80",
         10794 => x"ea38fe18",
         10795 => x"9c1a08fe",
         10796 => x"05595680",
         10797 => x"5c757827",
         10798 => x"8d388a19",
         10799 => x"22767129",
         10800 => x"b01b0805",
         10801 => x"5d5e7bb4",
         10802 => x"1a0cb819",
         10803 => x"58848078",
         10804 => x"57558076",
         10805 => x"70810558",
         10806 => x"34ff1555",
         10807 => x"74f43874",
         10808 => x"568a1922",
         10809 => x"55757527",
         10810 => x"81803881",
         10811 => x"54751c53",
         10812 => x"77528119",
         10813 => x"3351e4b2",
         10814 => x"3f84bb84",
         10815 => x"0880e738",
         10816 => x"811656dd",
         10817 => x"397a9818",
         10818 => x"0c840b84",
         10819 => x"bb840c8f",
         10820 => x"3d0d0475",
         10821 => x"54b41908",
         10822 => x"53b81970",
         10823 => x"53811a33",
         10824 => x"5256e486",
         10825 => x"3f84bb84",
         10826 => x"0880f338",
         10827 => x"84bb8408",
         10828 => x"831a34b4",
         10829 => x"1908a81a",
         10830 => x"08315574",
         10831 => x"a01a0827",
         10832 => x"fee83882",
         10833 => x"19335c7b",
         10834 => x"822e0981",
         10835 => x"06fedb38",
         10836 => x"8154b419",
         10837 => x"08a01a08",
         10838 => x"05537552",
         10839 => x"81193351",
         10840 => x"e3c83ffe",
         10841 => x"c5398a19",
         10842 => x"22557483",
         10843 => x"ffff0655",
         10844 => x"74762e09",
         10845 => x"8106a738",
         10846 => x"7c94180c",
         10847 => x"fe1d9c1a",
         10848 => x"08fe055e",
         10849 => x"56805875",
         10850 => x"7d27fd85",
         10851 => x"388a1922",
         10852 => x"767129b0",
         10853 => x"1b080598",
         10854 => x"190c5cfc",
         10855 => x"f839810b",
         10856 => x"84bb840c",
         10857 => x"8f3d0d04",
         10858 => x"ee3d0d64",
         10859 => x"66415c84",
         10860 => x"7c085a5b",
         10861 => x"81ff7098",
         10862 => x"1e08585e",
         10863 => x"5e75802e",
         10864 => x"82d238b8",
         10865 => x"195f755a",
         10866 => x"8058b419",
         10867 => x"08762e82",
         10868 => x"d1388319",
         10869 => x"33785855",
         10870 => x"74782e09",
         10871 => x"81068194",
         10872 => x"38815475",
         10873 => x"53b81952",
         10874 => x"81193351",
         10875 => x"e1bd3f84",
         10876 => x"bb840880",
         10877 => x"2e8538ff",
         10878 => x"5a815779",
         10879 => x"b41a0c76",
         10880 => x"5b768290",
         10881 => x"389c1c08",
         10882 => x"70335858",
         10883 => x"76802e82",
         10884 => x"81388b18",
         10885 => x"33bf0670",
         10886 => x"81ff065b",
         10887 => x"4160861d",
         10888 => x"347681e5",
         10889 => x"32703078",
         10890 => x"ae327030",
         10891 => x"72802571",
         10892 => x"80250754",
         10893 => x"45455755",
         10894 => x"74933874",
         10895 => x"7adf0643",
         10896 => x"5661882e",
         10897 => x"81bf3875",
         10898 => x"602e8186",
         10899 => x"3881ff5d",
         10900 => x"80527b51",
         10901 => x"faf63f84",
         10902 => x"bb84085b",
         10903 => x"84bb8408",
         10904 => x"81b23898",
         10905 => x"1c085675",
         10906 => x"fedc387a",
         10907 => x"84bb840c",
         10908 => x"943d0d04",
         10909 => x"8154b419",
         10910 => x"08537e52",
         10911 => x"81193351",
         10912 => x"e1a83f81",
         10913 => x"5784bb84",
         10914 => x"08782e09",
         10915 => x"8106feef",
         10916 => x"3884bb84",
         10917 => x"08831a34",
         10918 => x"b41908a8",
         10919 => x"1a083184",
         10920 => x"bb840858",
         10921 => x"5b7aa01a",
         10922 => x"0827feb5",
         10923 => x"38821933",
         10924 => x"4160822e",
         10925 => x"098106fe",
         10926 => x"a8388154",
         10927 => x"b41908a0",
         10928 => x"1a080553",
         10929 => x"7e528119",
         10930 => x"3351e0de",
         10931 => x"3f7757fe",
         10932 => x"9039798f",
         10933 => x"2e098106",
         10934 => x"81e73876",
         10935 => x"862a8106",
         10936 => x"5b7a802e",
         10937 => x"93388d18",
         10938 => x"337781bf",
         10939 => x"0670901f",
         10940 => x"087fac05",
         10941 => x"0c595e5e",
         10942 => x"767d2eab",
         10943 => x"3881ff55",
         10944 => x"745dfecc",
         10945 => x"39815675",
         10946 => x"602e0981",
         10947 => x"06febe38",
         10948 => x"c139845b",
         10949 => x"800b981d",
         10950 => x"0c7a84bb",
         10951 => x"840c943d",
         10952 => x"0d04775b",
         10953 => x"fddf398d",
         10954 => x"1833577d",
         10955 => x"772e0981",
         10956 => x"06cb388c",
         10957 => x"19089b19",
         10958 => x"339a1a33",
         10959 => x"71882b07",
         10960 => x"58564175",
         10961 => x"ffb73877",
         10962 => x"337081bf",
         10963 => x"068d29f3",
         10964 => x"05515a81",
         10965 => x"76585b83",
         10966 => x"e7841733",
         10967 => x"78058111",
         10968 => x"33713371",
         10969 => x"882b0752",
         10970 => x"44567a80",
         10971 => x"2e80c538",
         10972 => x"7981fe26",
         10973 => x"ff873879",
         10974 => x"10610576",
         10975 => x"5c427562",
         10976 => x"23811a5a",
         10977 => x"8117578c",
         10978 => x"7727cc38",
         10979 => x"77337086",
         10980 => x"2a810659",
         10981 => x"5777802e",
         10982 => x"90387981",
         10983 => x"fe26fedd",
         10984 => x"38791061",
         10985 => x"05438063",
         10986 => x"23ff1d70",
         10987 => x"81ff065e",
         10988 => x"41fd9d39",
         10989 => x"7583ffff",
         10990 => x"2eca3881",
         10991 => x"ff55fec0",
         10992 => x"397ca838",
         10993 => x"7c558b57",
         10994 => x"74812a75",
         10995 => x"81802905",
         10996 => x"78708105",
         10997 => x"5a33407f",
         10998 => x"057081ff",
         10999 => x"06ff1959",
         11000 => x"565976e4",
         11001 => x"38747e2e",
         11002 => x"fd8138ff",
         11003 => x"0bac1d0c",
         11004 => x"7a84bb84",
         11005 => x"0c943d0d",
         11006 => x"04ef3d0d",
         11007 => x"6370085c",
         11008 => x"5c80527b",
         11009 => x"51f5cf3f",
         11010 => x"84bb8408",
         11011 => x"5a84bb84",
         11012 => x"08828038",
         11013 => x"81ff7040",
         11014 => x"5dff0bac",
         11015 => x"1d0cb81b",
         11016 => x"5e981c08",
         11017 => x"568058b4",
         11018 => x"1b08762e",
         11019 => x"82cc3883",
         11020 => x"1b337858",
         11021 => x"5574782e",
         11022 => x"09810681",
         11023 => x"df388154",
         11024 => x"7553b81b",
         11025 => x"52811b33",
         11026 => x"51dce03f",
         11027 => x"84bb8408",
         11028 => x"802e8538",
         11029 => x"ff568157",
         11030 => x"75b41c0c",
         11031 => x"765a7681",
         11032 => x"b2389c1c",
         11033 => x"08703358",
         11034 => x"5976802e",
         11035 => x"8499388b",
         11036 => x"1933bf06",
         11037 => x"7081ff06",
         11038 => x"57587786",
         11039 => x"1d347681",
         11040 => x"e52e80f2",
         11041 => x"3875832a",
         11042 => x"81065575",
         11043 => x"8f2e81ef",
         11044 => x"387480e2",
         11045 => x"38758f2e",
         11046 => x"81e5387c",
         11047 => x"aa38787d",
         11048 => x"56588b57",
         11049 => x"74812a75",
         11050 => x"81802905",
         11051 => x"78708105",
         11052 => x"5a335776",
         11053 => x"057081ff",
         11054 => x"06ff1959",
         11055 => x"565d76e4",
         11056 => x"38747f2e",
         11057 => x"80cd38ab",
         11058 => x"1c338106",
         11059 => x"5776a738",
         11060 => x"8b0ba01d",
         11061 => x"59577870",
         11062 => x"81055a33",
         11063 => x"78708105",
         11064 => x"5a337171",
         11065 => x"31ff1a5a",
         11066 => x"58424076",
         11067 => x"802e81dc",
         11068 => x"3875802e",
         11069 => x"e13881ff",
         11070 => x"5dff0bac",
         11071 => x"1d0c8052",
         11072 => x"7b51f5c8",
         11073 => x"3f84bb84",
         11074 => x"085a84bb",
         11075 => x"8408802e",
         11076 => x"fe8f3879",
         11077 => x"84bb840c",
         11078 => x"933d0d04",
         11079 => x"8154b41b",
         11080 => x"08537d52",
         11081 => x"811b3351",
         11082 => x"dc803f81",
         11083 => x"5784bb84",
         11084 => x"08782e09",
         11085 => x"8106fea4",
         11086 => x"3884bb84",
         11087 => x"08831c34",
         11088 => x"b41b08a8",
         11089 => x"1c083184",
         11090 => x"bb840858",
         11091 => x"5978a01c",
         11092 => x"0827fdea",
         11093 => x"38821b33",
         11094 => x"5a79822e",
         11095 => x"098106fd",
         11096 => x"dd388154",
         11097 => x"b41b08a0",
         11098 => x"1c080553",
         11099 => x"7d52811b",
         11100 => x"3351dbb6",
         11101 => x"3f7757fd",
         11102 => x"c539775a",
         11103 => x"fde439ab",
         11104 => x"1c337086",
         11105 => x"2a810642",
         11106 => x"5560fef2",
         11107 => x"3876862a",
         11108 => x"81065a79",
         11109 => x"802e9338",
         11110 => x"8d193377",
         11111 => x"81bf0670",
         11112 => x"901f087f",
         11113 => x"ac050c59",
         11114 => x"5e5f767d",
         11115 => x"2eaf3881",
         11116 => x"ff55745d",
         11117 => x"80527b51",
         11118 => x"f4923f84",
         11119 => x"bb84085a",
         11120 => x"84bb8408",
         11121 => x"802efcd9",
         11122 => x"38fec839",
         11123 => x"75802efe",
         11124 => x"c23881ff",
         11125 => x"5dff0bac",
         11126 => x"1d0cfea2",
         11127 => x"398d1933",
         11128 => x"577e772e",
         11129 => x"098106c7",
         11130 => x"388c1b08",
         11131 => x"9b1a339a",
         11132 => x"1b337188",
         11133 => x"2b075942",
         11134 => x"4076ffb3",
         11135 => x"38783370",
         11136 => x"bf068d29",
         11137 => x"f3055b55",
         11138 => x"81775956",
         11139 => x"83e78418",
         11140 => x"33790581",
         11141 => x"11337133",
         11142 => x"71882b07",
         11143 => x"52425775",
         11144 => x"802e80ed",
         11145 => x"387981fe",
         11146 => x"26ff8438",
         11147 => x"765181a0",
         11148 => x"d13f84bb",
         11149 => x"84087a10",
         11150 => x"61057022",
         11151 => x"5343811b",
         11152 => x"5b5681a0",
         11153 => x"bd3f7584",
         11154 => x"bb84082e",
         11155 => x"098106fe",
         11156 => x"de387656",
         11157 => x"8118588c",
         11158 => x"7827ffb0",
         11159 => x"38783370",
         11160 => x"862a8106",
         11161 => x"56597580",
         11162 => x"2e923874",
         11163 => x"802e8d38",
         11164 => x"79106005",
         11165 => x"70224141",
         11166 => x"7ffeb438",
         11167 => x"ff1d7081",
         11168 => x"ff065e5a",
         11169 => x"feae3984",
         11170 => x"0b84bb84",
         11171 => x"0c933d0d",
         11172 => x"047683ff",
         11173 => x"ff2effbc",
         11174 => x"3881ff55",
         11175 => x"fe9439ea",
         11176 => x"3d0d6870",
         11177 => x"0870ab13",
         11178 => x"3381a006",
         11179 => x"585a5d5e",
         11180 => x"86567485",
         11181 => x"b538748c",
         11182 => x"1d087022",
         11183 => x"57575d74",
         11184 => x"802e8e38",
         11185 => x"811d7010",
         11186 => x"17702251",
         11187 => x"565d74f4",
         11188 => x"38953da0",
         11189 => x"1f5b408c",
         11190 => x"607b5858",
         11191 => x"55757081",
         11192 => x"05573377",
         11193 => x"70810559",
         11194 => x"34ff1555",
         11195 => x"74ef3802",
         11196 => x"80db0533",
         11197 => x"70810658",
         11198 => x"5676802e",
         11199 => x"82aa3880",
         11200 => x"c00bab1f",
         11201 => x"34810b94",
         11202 => x"3d405b8c",
         11203 => x"1c087b58",
         11204 => x"598b7a61",
         11205 => x"5a575577",
         11206 => x"70810559",
         11207 => x"33767081",
         11208 => x"055834ff",
         11209 => x"155574ef",
         11210 => x"38857b27",
         11211 => x"80c2387a",
         11212 => x"79225657",
         11213 => x"74802eb8",
         11214 => x"3874821a",
         11215 => x"5a568f58",
         11216 => x"75810677",
         11217 => x"10077681",
         11218 => x"2a7083ff",
         11219 => x"ff067290",
         11220 => x"2a810644",
         11221 => x"58565760",
         11222 => x"802e8738",
         11223 => x"7684a0a1",
         11224 => x"3257ff18",
         11225 => x"58778025",
         11226 => x"d7387822",
         11227 => x"5574ca38",
         11228 => x"87028405",
         11229 => x"80cf0557",
         11230 => x"5876b007",
         11231 => x"bf0655b9",
         11232 => x"75278438",
         11233 => x"87155574",
         11234 => x"7634ff16",
         11235 => x"ff197884",
         11236 => x"2a595956",
         11237 => x"76e33877",
         11238 => x"1f5980fe",
         11239 => x"7934767a",
         11240 => x"58568078",
         11241 => x"27a03879",
         11242 => x"335574a0",
         11243 => x"2e983881",
         11244 => x"16567578",
         11245 => x"2788a238",
         11246 => x"751a7033",
         11247 => x"565774a0",
         11248 => x"2e098106",
         11249 => x"ea388116",
         11250 => x"56a05577",
         11251 => x"87268e38",
         11252 => x"983d7805",
         11253 => x"ec058119",
         11254 => x"71335759",
         11255 => x"41747734",
         11256 => x"87762787",
         11257 => x"f4387d51",
         11258 => x"f88f3f84",
         11259 => x"bb84088b",
         11260 => x"38811b5b",
         11261 => x"80e37b27",
         11262 => x"fe913887",
         11263 => x"567a80e4",
         11264 => x"2e82e738",
         11265 => x"84bb8408",
         11266 => x"5684bb84",
         11267 => x"08842e09",
         11268 => x"810682d6",
         11269 => x"380280db",
         11270 => x"0533ab1f",
         11271 => x"347d0802",
         11272 => x"840580db",
         11273 => x"05335758",
         11274 => x"75812a81",
         11275 => x"065f815b",
         11276 => x"7e802e90",
         11277 => x"388d528c",
         11278 => x"1d51fe88",
         11279 => x"e83f84bb",
         11280 => x"84081b5b",
         11281 => x"80527d51",
         11282 => x"ed8c3f84",
         11283 => x"bb840856",
         11284 => x"84bb8408",
         11285 => x"81823884",
         11286 => x"bb8408b8",
         11287 => x"195e5998",
         11288 => x"1e085680",
         11289 => x"57b41808",
         11290 => x"762e85f3",
         11291 => x"38831833",
         11292 => x"407f772e",
         11293 => x"09810682",
         11294 => x"a3388154",
         11295 => x"7553b818",
         11296 => x"52811833",
         11297 => x"51d4a43f",
         11298 => x"84bb8408",
         11299 => x"802e8538",
         11300 => x"ff568157",
         11301 => x"75b4190c",
         11302 => x"765676bc",
         11303 => x"389c1e08",
         11304 => x"70335642",
         11305 => x"7481e52e",
         11306 => x"81c93874",
         11307 => x"30708025",
         11308 => x"7807565f",
         11309 => x"74802e81",
         11310 => x"c9388119",
         11311 => x"59787b2e",
         11312 => x"86893881",
         11313 => x"527d51ee",
         11314 => x"833f84bb",
         11315 => x"84085684",
         11316 => x"bb840880",
         11317 => x"2eff8838",
         11318 => x"87587584",
         11319 => x"2e818938",
         11320 => x"75587581",
         11321 => x"8338ff1b",
         11322 => x"407f81f3",
         11323 => x"38981e08",
         11324 => x"57b41c08",
         11325 => x"772eaf38",
         11326 => x"831c3378",
         11327 => x"57407f84",
         11328 => x"82388154",
         11329 => x"7653b81c",
         11330 => x"52811c33",
         11331 => x"51d39c3f",
         11332 => x"84bb8408",
         11333 => x"802e8538",
         11334 => x"ff578156",
         11335 => x"76b41d0c",
         11336 => x"75587580",
         11337 => x"c338a00b",
         11338 => x"9c1f0857",
         11339 => x"55807670",
         11340 => x"81055834",
         11341 => x"ff155574",
         11342 => x"f4388b0b",
         11343 => x"9c1f087b",
         11344 => x"58585575",
         11345 => x"70810557",
         11346 => x"33777081",
         11347 => x"055934ff",
         11348 => x"155574ef",
         11349 => x"389c1e08",
         11350 => x"ab1f3398",
         11351 => x"065e5a7c",
         11352 => x"8c1b3481",
         11353 => x"0b831d34",
         11354 => x"77567584",
         11355 => x"bb840c98",
         11356 => x"3d0d0481",
         11357 => x"75307080",
         11358 => x"25720757",
         11359 => x"405774fe",
         11360 => x"b9387459",
         11361 => x"81527d51",
         11362 => x"ecc23f84",
         11363 => x"bb840856",
         11364 => x"84bb8408",
         11365 => x"802efdc7",
         11366 => x"38febd39",
         11367 => x"8154b418",
         11368 => x"08537c52",
         11369 => x"81183351",
         11370 => x"d3803f84",
         11371 => x"bb840877",
         11372 => x"2e098106",
         11373 => x"83bf3884",
         11374 => x"bb840883",
         11375 => x"1934b418",
         11376 => x"08a81908",
         11377 => x"315574a0",
         11378 => x"1908278b",
         11379 => x"38821833",
         11380 => x"4160822e",
         11381 => x"84ac3884",
         11382 => x"bb840857",
         11383 => x"fd9c397f",
         11384 => x"852b901f",
         11385 => x"08713153",
         11386 => x"587d51e9",
         11387 => x"e93f84bb",
         11388 => x"84085884",
         11389 => x"bb8408fe",
         11390 => x"ef387984",
         11391 => x"bb840856",
         11392 => x"588b5774",
         11393 => x"812a7581",
         11394 => x"80290578",
         11395 => x"7081055a",
         11396 => x"33577605",
         11397 => x"7081ff06",
         11398 => x"ff195956",
         11399 => x"5d76e438",
         11400 => x"7481ff06",
         11401 => x"b81d4341",
         11402 => x"981e0857",
         11403 => x"8056b41c",
         11404 => x"08772eb2",
         11405 => x"38831c33",
         11406 => x"5b7a762e",
         11407 => x"09810682",
         11408 => x"c9388154",
         11409 => x"7653b81c",
         11410 => x"52811c33",
         11411 => x"51d0dc3f",
         11412 => x"84bb8408",
         11413 => x"802e8538",
         11414 => x"ff578156",
         11415 => x"76b41d0c",
         11416 => x"755875fe",
         11417 => x"83388c1c",
         11418 => x"089c1f08",
         11419 => x"6181ff06",
         11420 => x"5f5c5f60",
         11421 => x"8d1c348f",
         11422 => x"0b8b1c34",
         11423 => x"758c1c34",
         11424 => x"759a1c34",
         11425 => x"759b1c34",
         11426 => x"7c8d29f3",
         11427 => x"0576775a",
         11428 => x"58597683",
         11429 => x"ffff2e8b",
         11430 => x"3878101f",
         11431 => x"7022811b",
         11432 => x"5b585683",
         11433 => x"e7841833",
         11434 => x"7b055576",
         11435 => x"75708105",
         11436 => x"57347688",
         11437 => x"2a567575",
         11438 => x"34768538",
         11439 => x"83ffff57",
         11440 => x"8118588c",
         11441 => x"7827cb38",
         11442 => x"7683ffff",
         11443 => x"2e81b338",
         11444 => x"78101f70",
         11445 => x"22585876",
         11446 => x"802e81a6",
         11447 => x"387c7b34",
         11448 => x"810b831d",
         11449 => x"3480527d",
         11450 => x"51e9e13f",
         11451 => x"84bb8408",
         11452 => x"5884bb84",
         11453 => x"08fcf138",
         11454 => x"7fff0540",
         11455 => x"7ffea938",
         11456 => x"fbeb3981",
         11457 => x"54b41c08",
         11458 => x"53b81c70",
         11459 => x"53811d33",
         11460 => x"5259d096",
         11461 => x"3f815684",
         11462 => x"bb8408fc",
         11463 => x"833884bb",
         11464 => x"8408831d",
         11465 => x"34b41c08",
         11466 => x"a81d0831",
         11467 => x"84bb8408",
         11468 => x"574160a0",
         11469 => x"1d0827fb",
         11470 => x"c938821c",
         11471 => x"33426182",
         11472 => x"2e098106",
         11473 => x"fbbc3881",
         11474 => x"54b41c08",
         11475 => x"a01d0805",
         11476 => x"53785281",
         11477 => x"1c3351cf",
         11478 => x"d13f7756",
         11479 => x"fba43976",
         11480 => x"9c1f0870",
         11481 => x"33574356",
         11482 => x"7481e52e",
         11483 => x"098106fa",
         11484 => x"ba38fbff",
         11485 => x"39817057",
         11486 => x"5776802e",
         11487 => x"fa9f38fa",
         11488 => x"d7397c80",
         11489 => x"c0075dfe",
         11490 => x"d4398154",
         11491 => x"b41c0853",
         11492 => x"6152811c",
         11493 => x"3351cf92",
         11494 => x"3f84bb84",
         11495 => x"08762e09",
         11496 => x"8106bc38",
         11497 => x"84bb8408",
         11498 => x"831d34b4",
         11499 => x"1c08a81d",
         11500 => x"08315574",
         11501 => x"a01d0827",
         11502 => x"8a38821c",
         11503 => x"335f7e82",
         11504 => x"2eaa3884",
         11505 => x"bb840856",
         11506 => x"fcf83975",
         11507 => x"ff1c4158",
         11508 => x"7f802efa",
         11509 => x"9838fc87",
         11510 => x"39751a57",
         11511 => x"f7e83981",
         11512 => x"70595675",
         11513 => x"802efcfe",
         11514 => x"38fafd39",
         11515 => x"8154b41c",
         11516 => x"08a01d08",
         11517 => x"05536152",
         11518 => x"811c3351",
         11519 => x"ceac3ffc",
         11520 => x"c1398154",
         11521 => x"b41808a0",
         11522 => x"19080553",
         11523 => x"7c528118",
         11524 => x"3351ce96",
         11525 => x"3ff8e339",
         11526 => x"f33d0d7f",
         11527 => x"61710840",
         11528 => x"5e5c800b",
         11529 => x"961e3498",
         11530 => x"1c08802e",
         11531 => x"82b538ac",
         11532 => x"1c08ff2e",
         11533 => x"80d93880",
         11534 => x"7071608c",
         11535 => x"05087022",
         11536 => x"57585b5c",
         11537 => x"5872782e",
         11538 => x"bc387754",
         11539 => x"74147022",
         11540 => x"811b5b55",
         11541 => x"567a8295",
         11542 => x"3880d080",
         11543 => x"147083ff",
         11544 => x"ff06585a",
         11545 => x"768fff26",
         11546 => x"82833873",
         11547 => x"791a7611",
         11548 => x"70225d58",
         11549 => x"555b79d4",
         11550 => x"387a3070",
         11551 => x"80257030",
         11552 => x"7a065a5c",
         11553 => x"5e7c1894",
         11554 => x"0557800b",
         11555 => x"82183480",
         11556 => x"70891f59",
         11557 => x"57589c1c",
         11558 => x"08167033",
         11559 => x"81185856",
         11560 => x"5374a02e",
         11561 => x"b2387485",
         11562 => x"2e81bc38",
         11563 => x"75893270",
         11564 => x"30707207",
         11565 => x"8025555b",
         11566 => x"54778b26",
         11567 => x"90387280",
         11568 => x"2e8b38ae",
         11569 => x"77708105",
         11570 => x"59348118",
         11571 => x"58747770",
         11572 => x"81055934",
         11573 => x"8118588a",
         11574 => x"7627ffba",
         11575 => x"387c1888",
         11576 => x"0555800b",
         11577 => x"81163496",
         11578 => x"1d335372",
         11579 => x"a5387781",
         11580 => x"f338bf0b",
         11581 => x"961e3481",
         11582 => x"577c1794",
         11583 => x"0556800b",
         11584 => x"8217349c",
         11585 => x"1c088c11",
         11586 => x"33555373",
         11587 => x"89387389",
         11588 => x"1e349c1c",
         11589 => x"08538b13",
         11590 => x"33881e34",
         11591 => x"9c1c089c",
         11592 => x"11831133",
         11593 => x"82123371",
         11594 => x"902b7188",
         11595 => x"2b078114",
         11596 => x"33707207",
         11597 => x"882b7533",
         11598 => x"7107640c",
         11599 => x"59971633",
         11600 => x"96173371",
         11601 => x"882b075f",
         11602 => x"415b405a",
         11603 => x"565b5577",
         11604 => x"861e2399",
         11605 => x"15339816",
         11606 => x"3371882b",
         11607 => x"075d547b",
         11608 => x"841e238f",
         11609 => x"3d0d0481",
         11610 => x"e555fec0",
         11611 => x"39771d96",
         11612 => x"1181ff7a",
         11613 => x"31585b57",
         11614 => x"83b5527a",
         11615 => x"902b7407",
         11616 => x"518190d0",
         11617 => x"3f84bb84",
         11618 => x"0883ffff",
         11619 => x"065581ff",
         11620 => x"7527ad38",
         11621 => x"81762781",
         11622 => x"b3387488",
         11623 => x"2a54737a",
         11624 => x"34749718",
         11625 => x"34827805",
         11626 => x"58800b8c",
         11627 => x"1f08565b",
         11628 => x"78197511",
         11629 => x"70225c57",
         11630 => x"5479fd90",
         11631 => x"38fdba39",
         11632 => x"74307630",
         11633 => x"70780780",
         11634 => x"25728025",
         11635 => x"07585557",
         11636 => x"7580f938",
         11637 => x"747a3481",
         11638 => x"78055880",
         11639 => x"0b8c1f08",
         11640 => x"565bcd39",
         11641 => x"7273891f",
         11642 => x"335a5757",
         11643 => x"77802efe",
         11644 => x"88387c96",
         11645 => x"1e7e5759",
         11646 => x"54891433",
         11647 => x"ffbf115a",
         11648 => x"54789926",
         11649 => x"a4389c1c",
         11650 => x"088c1133",
         11651 => x"545b8876",
         11652 => x"27b43872",
         11653 => x"842a5372",
         11654 => x"81065e7d",
         11655 => x"802e8a38",
         11656 => x"a0147083",
         11657 => x"ffff0655",
         11658 => x"53737870",
         11659 => x"81055a34",
         11660 => x"81168116",
         11661 => x"81197189",
         11662 => x"13335e57",
         11663 => x"59565679",
         11664 => x"ffb738fd",
         11665 => x"b4397283",
         11666 => x"2a53cc39",
         11667 => x"807b3070",
         11668 => x"80257030",
         11669 => x"7306535d",
         11670 => x"5f58fca9",
         11671 => x"39ef3d0d",
         11672 => x"63700870",
         11673 => x"42575c80",
         11674 => x"65703357",
         11675 => x"555374af",
         11676 => x"2e833881",
         11677 => x"537480dc",
         11678 => x"2e81df38",
         11679 => x"72802e81",
         11680 => x"d9389816",
         11681 => x"08881d0c",
         11682 => x"7333963d",
         11683 => x"943d4142",
         11684 => x"559f7527",
         11685 => x"82a73873",
         11686 => x"428c1608",
         11687 => x"58805761",
         11688 => x"70708105",
         11689 => x"52335553",
         11690 => x"7381df38",
         11691 => x"727f0c73",
         11692 => x"ff2e81ec",
         11693 => x"3883ffff",
         11694 => x"74278b38",
         11695 => x"76101856",
         11696 => x"80762381",
         11697 => x"17577383",
         11698 => x"ffff0670",
         11699 => x"af327030",
         11700 => x"9f732771",
         11701 => x"80250757",
         11702 => x"5b5b5573",
         11703 => x"82903874",
         11704 => x"80dc2e82",
         11705 => x"89387480",
         11706 => x"ff26b238",
         11707 => x"83e6a00b",
         11708 => x"83e6a033",
         11709 => x"7081ff06",
         11710 => x"56545673",
         11711 => x"802e81ab",
         11712 => x"3873752e",
         11713 => x"8f388116",
         11714 => x"70337081",
         11715 => x"ff065654",
         11716 => x"5673ee38",
         11717 => x"7281ff06",
         11718 => x"5b7a8184",
         11719 => x"387681fe",
         11720 => x"2680fd38",
         11721 => x"7610185d",
         11722 => x"747d2381",
         11723 => x"17627070",
         11724 => x"81055233",
         11725 => x"56545773",
         11726 => x"802efef0",
         11727 => x"3880cb39",
         11728 => x"817380dc",
         11729 => x"32703070",
         11730 => x"80257307",
         11731 => x"51555855",
         11732 => x"72802ea1",
         11733 => x"38811470",
         11734 => x"46548074",
         11735 => x"33545572",
         11736 => x"af2edd38",
         11737 => x"7280dc32",
         11738 => x"70307080",
         11739 => x"25770751",
         11740 => x"545772e1",
         11741 => x"3872881d",
         11742 => x"0c733396",
         11743 => x"3d943d41",
         11744 => x"4255749f",
         11745 => x"26fe9038",
         11746 => x"b43983b5",
         11747 => x"52735181",
         11748 => x"8dae3f84",
         11749 => x"bb840883",
         11750 => x"ffff0654",
         11751 => x"73fe8d38",
         11752 => x"86547384",
         11753 => x"bb840c93",
         11754 => x"3d0d0483",
         11755 => x"e6a03370",
         11756 => x"81ff065c",
         11757 => x"537a802e",
         11758 => x"fee338e4",
         11759 => x"39ff800b",
         11760 => x"ab1d3480",
         11761 => x"527b51de",
         11762 => x"8d3f84bb",
         11763 => x"840884bb",
         11764 => x"840c933d",
         11765 => x"0d048173",
         11766 => x"80dc3270",
         11767 => x"30708025",
         11768 => x"73074155",
         11769 => x"5a567d80",
         11770 => x"2ea13881",
         11771 => x"14428062",
         11772 => x"70335555",
         11773 => x"5672af2e",
         11774 => x"dd387280",
         11775 => x"dc327030",
         11776 => x"70802578",
         11777 => x"07405459",
         11778 => x"7de13873",
         11779 => x"610c9f75",
         11780 => x"27822b5a",
         11781 => x"76812e84",
         11782 => x"f8387682",
         11783 => x"2e83d138",
         11784 => x"76175976",
         11785 => x"802ea738",
         11786 => x"76177811",
         11787 => x"fe057022",
         11788 => x"70a03270",
         11789 => x"30709f2a",
         11790 => x"5242565f",
         11791 => x"56597cae",
         11792 => x"2e843872",
         11793 => x"8938ff17",
         11794 => x"5776dd38",
         11795 => x"76597719",
         11796 => x"56807623",
         11797 => x"76802efe",
         11798 => x"c7388078",
         11799 => x"227083ff",
         11800 => x"ff067258",
         11801 => x"5d55567a",
         11802 => x"a02e82e6",
         11803 => x"387383ff",
         11804 => x"ff065372",
         11805 => x"ae2e82f1",
         11806 => x"3876802e",
         11807 => x"aa387719",
         11808 => x"fe057022",
         11809 => x"5a5478ae",
         11810 => x"2e9d3876",
         11811 => x"1018fe05",
         11812 => x"54ff1757",
         11813 => x"76802e8f",
         11814 => x"38fe1470",
         11815 => x"225e547c",
         11816 => x"ae2e0981",
         11817 => x"06eb388b",
         11818 => x"0ba01d55",
         11819 => x"53a07470",
         11820 => x"81055634",
         11821 => x"ff135372",
         11822 => x"f4387273",
         11823 => x"5c5e8878",
         11824 => x"16702281",
         11825 => x"19595754",
         11826 => x"5d74802e",
         11827 => x"80ed3874",
         11828 => x"a02e83d0",
         11829 => x"3874ae32",
         11830 => x"70307080",
         11831 => x"25555a54",
         11832 => x"75772e85",
         11833 => x"ce387283",
         11834 => x"bb387259",
         11835 => x"7c7b2683",
         11836 => x"38815975",
         11837 => x"77327030",
         11838 => x"70720780",
         11839 => x"25707c07",
         11840 => x"51515454",
         11841 => x"72802e83",
         11842 => x"e0387c8b",
         11843 => x"2e868338",
         11844 => x"75772e8a",
         11845 => x"38798307",
         11846 => x"5a757726",
         11847 => x"9e387656",
         11848 => x"885b8b7e",
         11849 => x"822b81fc",
         11850 => x"06771857",
         11851 => x"5f5d7715",
         11852 => x"70228118",
         11853 => x"58565374",
         11854 => x"ff9538a0",
         11855 => x"1c335776",
         11856 => x"81e52e83",
         11857 => x"84387c88",
         11858 => x"2e82e338",
         11859 => x"7d8c0658",
         11860 => x"778c2e82",
         11861 => x"ed387d83",
         11862 => x"06557483",
         11863 => x"2e82e338",
         11864 => x"79812a81",
         11865 => x"0656759d",
         11866 => x"387d8106",
         11867 => x"5d7c802e",
         11868 => x"85387990",
         11869 => x"075a7d82",
         11870 => x"2a81065e",
         11871 => x"7d802e85",
         11872 => x"38798807",
         11873 => x"5a79ab1d",
         11874 => x"347b51e4",
         11875 => x"ec3f84bb",
         11876 => x"8408ab1d",
         11877 => x"33565484",
         11878 => x"bb840880",
         11879 => x"2e81ac38",
         11880 => x"84bb8408",
         11881 => x"842e0981",
         11882 => x"06fbf738",
         11883 => x"74852a81",
         11884 => x"065a7980",
         11885 => x"2e84f038",
         11886 => x"74822a81",
         11887 => x"06597882",
         11888 => x"98387b08",
         11889 => x"65555673",
         11890 => x"428c1608",
         11891 => x"588057f9",
         11892 => x"ce398116",
         11893 => x"70117911",
         11894 => x"70224040",
         11895 => x"56567ca0",
         11896 => x"2ef03875",
         11897 => x"802efd85",
         11898 => x"38798307",
         11899 => x"5afd8a39",
         11900 => x"82182256",
         11901 => x"75ae2e09",
         11902 => x"8106fcac",
         11903 => x"38772254",
         11904 => x"73ae2e09",
         11905 => x"8106fca0",
         11906 => x"38761018",
         11907 => x"5b807b23",
         11908 => x"800ba01d",
         11909 => x"5653ae54",
         11910 => x"76732683",
         11911 => x"38a05473",
         11912 => x"75708105",
         11913 => x"57348113",
         11914 => x"538a7327",
         11915 => x"e93879a0",
         11916 => x"075877ab",
         11917 => x"1d347b51",
         11918 => x"e3bf3f84",
         11919 => x"bb8408ab",
         11920 => x"1d335654",
         11921 => x"84bb8408",
         11922 => x"fed63874",
         11923 => x"822a8106",
         11924 => x"5877face",
         11925 => x"38861c33",
         11926 => x"70842a81",
         11927 => x"06565d74",
         11928 => x"802e83cd",
         11929 => x"38901c08",
         11930 => x"83ff0660",
         11931 => x"0580d311",
         11932 => x"3380d212",
         11933 => x"3371882b",
         11934 => x"07623341",
         11935 => x"5754547d",
         11936 => x"832e82d8",
         11937 => x"3874881d",
         11938 => x"0c7b0865",
         11939 => x"5556feb7",
         11940 => x"39772255",
         11941 => x"74ae2efe",
         11942 => x"f0387617",
         11943 => x"5976fb88",
         11944 => x"38fbab39",
         11945 => x"79830776",
         11946 => x"17565afd",
         11947 => x"81397d82",
         11948 => x"2b81fc06",
         11949 => x"708c0659",
         11950 => x"5e778c2e",
         11951 => x"098106fd",
         11952 => x"95387982",
         11953 => x"075afd98",
         11954 => x"39850ba0",
         11955 => x"1d347c88",
         11956 => x"2e098106",
         11957 => x"fcf638d6",
         11958 => x"39ff800b",
         11959 => x"ab1d3480",
         11960 => x"0b84bb84",
         11961 => x"0c933d0d",
         11962 => x"047480ff",
         11963 => x"269d3881",
         11964 => x"ff752780",
         11965 => x"c938ff1d",
         11966 => x"59787b26",
         11967 => x"81f73879",
         11968 => x"83077d77",
         11969 => x"18575c5a",
         11970 => x"fca43979",
         11971 => x"82075a83",
         11972 => x"b5527451",
         11973 => x"8185bd3f",
         11974 => x"84bb8408",
         11975 => x"83ffff06",
         11976 => x"70872a81",
         11977 => x"065a5578",
         11978 => x"802ec438",
         11979 => x"7480ff06",
         11980 => x"83e79411",
         11981 => x"33565474",
         11982 => x"81ff26ff",
         11983 => x"b9387480",
         11984 => x"2e818538",
         11985 => x"83e6ac0b",
         11986 => x"83e6ac33",
         11987 => x"7081ff06",
         11988 => x"56545973",
         11989 => x"802e80e0",
         11990 => x"3873752e",
         11991 => x"8f388119",
         11992 => x"70337081",
         11993 => x"ff065654",
         11994 => x"5973ee38",
         11995 => x"7281ff06",
         11996 => x"597880d4",
         11997 => x"38ffbf15",
         11998 => x"54739926",
         11999 => x"8a387d82",
         12000 => x"077081ff",
         12001 => x"065f53ff",
         12002 => x"9f155978",
         12003 => x"99269338",
         12004 => x"7d810770",
         12005 => x"81ff06e0",
         12006 => x"177083ff",
         12007 => x"ff065856",
         12008 => x"5f537b1b",
         12009 => x"a0055974",
         12010 => x"7934811b",
         12011 => x"5b751655",
         12012 => x"fafc3980",
         12013 => x"53fab339",
         12014 => x"83e6ac33",
         12015 => x"7081ff06",
         12016 => x"5a537880",
         12017 => x"2effae38",
         12018 => x"80df7a83",
         12019 => x"077d1da0",
         12020 => x"055b5b55",
         12021 => x"74793481",
         12022 => x"1b5bd239",
         12023 => x"80cd1433",
         12024 => x"80cc1533",
         12025 => x"71982b71",
         12026 => x"902b0777",
         12027 => x"07881f0c",
         12028 => x"5a57fd95",
         12029 => x"397b1ba0",
         12030 => x"0575882a",
         12031 => x"54547274",
         12032 => x"34811b7c",
         12033 => x"11a0055a",
         12034 => x"5b747934",
         12035 => x"811b5bff",
         12036 => x"9c397983",
         12037 => x"07a01d33",
         12038 => x"585a7681",
         12039 => x"e52e0981",
         12040 => x"06faa338",
         12041 => x"fda33974",
         12042 => x"822a8106",
         12043 => x"5c7bf6f2",
         12044 => x"38850b84",
         12045 => x"bb840c93",
         12046 => x"3d0d04eb",
         12047 => x"3d0d6769",
         12048 => x"02880580",
         12049 => x"e7053342",
         12050 => x"425e8061",
         12051 => x"0cff7e08",
         12052 => x"70595b42",
         12053 => x"79802e85",
         12054 => x"d7387970",
         12055 => x"81055b33",
         12056 => x"709f2656",
         12057 => x"5675ba2e",
         12058 => x"85d03874",
         12059 => x"ed3875ba",
         12060 => x"2e85c738",
         12061 => x"84e2e033",
         12062 => x"56807624",
         12063 => x"85b23875",
         12064 => x"101084e2",
         12065 => x"cc057008",
         12066 => x"585a8c58",
         12067 => x"76802e85",
         12068 => x"96387661",
         12069 => x"0c7f81fe",
         12070 => x"0677335d",
         12071 => x"597b802e",
         12072 => x"9b388117",
         12073 => x"3351ffbb",
         12074 => x"b03f84bb",
         12075 => x"840881ff",
         12076 => x"06708106",
         12077 => x"5e587c80",
         12078 => x"2e869638",
         12079 => x"80773475",
         12080 => x"165d84ba",
         12081 => x"f81d3381",
         12082 => x"18348152",
         12083 => x"81173351",
         12084 => x"ffbba43f",
         12085 => x"84bb8408",
         12086 => x"81ff0670",
         12087 => x"81064156",
         12088 => x"83587f84",
         12089 => x"c2387880",
         12090 => x"2e8d3875",
         12091 => x"822a8106",
         12092 => x"418a5860",
         12093 => x"84b13880",
         12094 => x"5b7a8318",
         12095 => x"34ff0bb4",
         12096 => x"180c7a7b",
         12097 => x"5a558154",
         12098 => x"7a53b817",
         12099 => x"70538118",
         12100 => x"335258ff",
         12101 => x"bb953f84",
         12102 => x"bb84087b",
         12103 => x"2e8538ff",
         12104 => x"55815974",
         12105 => x"b4180c84",
         12106 => x"56789938",
         12107 => x"84b71733",
         12108 => x"84b61833",
         12109 => x"71882b07",
         12110 => x"56568356",
         12111 => x"7482d4d5",
         12112 => x"2e85a538",
         12113 => x"7581268b",
         12114 => x"3884baf9",
         12115 => x"1d334261",
         12116 => x"85bf3881",
         12117 => x"5875842e",
         12118 => x"83cd388d",
         12119 => x"58758126",
         12120 => x"83c53880",
         12121 => x"c4173380",
         12122 => x"c3183371",
         12123 => x"882b075e",
         12124 => x"597c8480",
         12125 => x"2e098106",
         12126 => x"83ad3880",
         12127 => x"cf173380",
         12128 => x"ce183371",
         12129 => x"882b0757",
         12130 => x"5a75a438",
         12131 => x"80dc1783",
         12132 => x"11338212",
         12133 => x"3371902b",
         12134 => x"71882b07",
         12135 => x"81143370",
         12136 => x"7207882b",
         12137 => x"75337107",
         12138 => x"565a4543",
         12139 => x"5e5f5675",
         12140 => x"a0180c80",
         12141 => x"c8173382",
         12142 => x"183480c8",
         12143 => x"1733ff11",
         12144 => x"7081ff06",
         12145 => x"5f40598d",
         12146 => x"587c8126",
         12147 => x"82d93878",
         12148 => x"81ff0676",
         12149 => x"712980c5",
         12150 => x"19335a5f",
         12151 => x"5a778a18",
         12152 => x"23775977",
         12153 => x"802e87c4",
         12154 => x"38ff1878",
         12155 => x"06426187",
         12156 => x"bb3880ca",
         12157 => x"173380c9",
         12158 => x"18337188",
         12159 => x"2b075640",
         12160 => x"74881823",
         12161 => x"74758f06",
         12162 => x"5e5a8d58",
         12163 => x"7c829838",
         12164 => x"80cc1733",
         12165 => x"80cb1833",
         12166 => x"71882b07",
         12167 => x"565c74a4",
         12168 => x"3880d817",
         12169 => x"83113382",
         12170 => x"12337190",
         12171 => x"2b71882b",
         12172 => x"07811433",
         12173 => x"70720788",
         12174 => x"2b753371",
         12175 => x"0753445a",
         12176 => x"58424242",
         12177 => x"80c71733",
         12178 => x"80c61833",
         12179 => x"71882b07",
         12180 => x"5d588d58",
         12181 => x"7b802e81",
         12182 => x"ce387d1c",
         12183 => x"7a842a05",
         12184 => x"5a797526",
         12185 => x"81c13878",
         12186 => x"52747a31",
         12187 => x"51fdecb5",
         12188 => x"3f84bb84",
         12189 => x"085684bb",
         12190 => x"8408802e",
         12191 => x"81a93884",
         12192 => x"bb840880",
         12193 => x"fffffff5",
         12194 => x"26833883",
         12195 => x"5d7583ff",
         12196 => x"f5268338",
         12197 => x"825d759f",
         12198 => x"f52685eb",
         12199 => x"38815d82",
         12200 => x"16709c19",
         12201 => x"0c7ba419",
         12202 => x"0c7b1d70",
         12203 => x"a81a0c7b",
         12204 => x"1db01a0c",
         12205 => x"57597c83",
         12206 => x"2e8a8738",
         12207 => x"8817225c",
         12208 => x"8d587b80",
         12209 => x"2e80e038",
         12210 => x"7d16ac18",
         12211 => x"0c781955",
         12212 => x"7c822e8d",
         12213 => x"38781019",
         12214 => x"70812a7a",
         12215 => x"81060556",
         12216 => x"5a83ff15",
         12217 => x"892a598d",
         12218 => x"5878a018",
         12219 => x"0826b838",
         12220 => x"ff0b9418",
         12221 => x"0cff0b90",
         12222 => x"180cff80",
         12223 => x"0b841834",
         12224 => x"7c832e86",
         12225 => x"96387c77",
         12226 => x"3484e2dc",
         12227 => x"2281055d",
         12228 => x"7c84e2dc",
         12229 => x"237c8618",
         12230 => x"2384e2e4",
         12231 => x"0b8c180c",
         12232 => x"800b9818",
         12233 => x"0c805877",
         12234 => x"84bb840c",
         12235 => x"973d0d04",
         12236 => x"8b0b84bb",
         12237 => x"840c973d",
         12238 => x"0d047633",
         12239 => x"d0117081",
         12240 => x"ff065757",
         12241 => x"58748926",
         12242 => x"91388217",
         12243 => x"7881ff06",
         12244 => x"d0055d59",
         12245 => x"787a2e87",
         12246 => x"fe38807e",
         12247 => x"0883e6f4",
         12248 => x"5f405c7c",
         12249 => x"087f5a5b",
         12250 => x"7a708105",
         12251 => x"5c337970",
         12252 => x"81055b33",
         12253 => x"ff9f125a",
         12254 => x"58567799",
         12255 => x"268938e0",
         12256 => x"167081ff",
         12257 => x"065755ff",
         12258 => x"9f175877",
         12259 => x"99268938",
         12260 => x"e0177081",
         12261 => x"ff065855",
         12262 => x"7530709f",
         12263 => x"2a595575",
         12264 => x"772e0981",
         12265 => x"06853877",
         12266 => x"ffbe3878",
         12267 => x"7a327030",
         12268 => x"7072079f",
         12269 => x"2a7a075d",
         12270 => x"58557a80",
         12271 => x"2e879838",
         12272 => x"811c841e",
         12273 => x"5e5c837c",
         12274 => x"25ff9838",
         12275 => x"6156f9a9",
         12276 => x"3978802e",
         12277 => x"fecf3877",
         12278 => x"822a8106",
         12279 => x"5e8a587d",
         12280 => x"fec53880",
         12281 => x"58fec039",
         12282 => x"7a783357",
         12283 => x"597581e9",
         12284 => x"2e098106",
         12285 => x"83388159",
         12286 => x"7581eb32",
         12287 => x"70307080",
         12288 => x"257b075a",
         12289 => x"5b5c7783",
         12290 => x"ad387581",
         12291 => x"e82e83a6",
         12292 => x"38933d77",
         12293 => x"575a8359",
         12294 => x"83fa1633",
         12295 => x"70595b7a",
         12296 => x"802ea538",
         12297 => x"84811633",
         12298 => x"84801733",
         12299 => x"71902b71",
         12300 => x"882b0783",
         12301 => x"ff193370",
         12302 => x"7207882b",
         12303 => x"83fe1b33",
         12304 => x"71075259",
         12305 => x"5b404040",
         12306 => x"777a7084",
         12307 => x"055c0cff",
         12308 => x"19901757",
         12309 => x"59788025",
         12310 => x"ffbe3884",
         12311 => x"baf91d33",
         12312 => x"7030709f",
         12313 => x"2a727131",
         12314 => x"9b3d7110",
         12315 => x"1005f005",
         12316 => x"84b61c44",
         12317 => x"5d52435b",
         12318 => x"4278085b",
         12319 => x"83567a80",
         12320 => x"2e80fb38",
         12321 => x"800b8318",
         12322 => x"34ff0bb4",
         12323 => x"180c7a55",
         12324 => x"80567aff",
         12325 => x"2ea53881",
         12326 => x"547a53b8",
         12327 => x"17528117",
         12328 => x"3351ffb4",
         12329 => x"863f84bb",
         12330 => x"8408762e",
         12331 => x"8538ff55",
         12332 => x"815674b4",
         12333 => x"180c8458",
         12334 => x"75bf3881",
         12335 => x"1f337f33",
         12336 => x"71882b07",
         12337 => x"5d5e8358",
         12338 => x"7b82d4d5",
         12339 => x"2e098106",
         12340 => x"a838800b",
         12341 => x"b8183357",
         12342 => x"587581e9",
         12343 => x"2e82b738",
         12344 => x"7581eb32",
         12345 => x"70307080",
         12346 => x"257a0742",
         12347 => x"42427fbc",
         12348 => x"387581e8",
         12349 => x"2eb63882",
         12350 => x"587781ff",
         12351 => x"0656800b",
         12352 => x"84baf91e",
         12353 => x"335d587b",
         12354 => x"782e0981",
         12355 => x"06833881",
         12356 => x"58817627",
         12357 => x"f8bd3877",
         12358 => x"802ef8b7",
         12359 => x"38811a84",
         12360 => x"1a5a5a83",
         12361 => x"7a27fed1",
         12362 => x"38f8a839",
         12363 => x"830b80ee",
         12364 => x"1883e6b4",
         12365 => x"405d587b",
         12366 => x"7081055d",
         12367 => x"337e7081",
         12368 => x"05403371",
         12369 => x"7131ff1b",
         12370 => x"5b525656",
         12371 => x"77802e80",
         12372 => x"c5387580",
         12373 => x"2ee13885",
         12374 => x"0b818a18",
         12375 => x"83e6b840",
         12376 => x"5d587b70",
         12377 => x"81055d33",
         12378 => x"7e708105",
         12379 => x"40337171",
         12380 => x"31ff1b5b",
         12381 => x"58424077",
         12382 => x"802e858e",
         12383 => x"3875802e",
         12384 => x"e1388258",
         12385 => x"fef3398d",
         12386 => x"587cfa93",
         12387 => x"387784bb",
         12388 => x"840c973d",
         12389 => x"0d047558",
         12390 => x"75802efe",
         12391 => x"dc38850b",
         12392 => x"818a1883",
         12393 => x"e6b8405d",
         12394 => x"58ffb739",
         12395 => x"8d0b84bb",
         12396 => x"840c973d",
         12397 => x"0d04830b",
         12398 => x"80ee1883",
         12399 => x"e6b45c5a",
         12400 => x"58787081",
         12401 => x"055a337a",
         12402 => x"7081055c",
         12403 => x"33717131",
         12404 => x"ff1b5b57",
         12405 => x"5f5f7780",
         12406 => x"2e83d138",
         12407 => x"74802ee1",
         12408 => x"38850b81",
         12409 => x"8a1883e6",
         12410 => x"b85c5a58",
         12411 => x"78708105",
         12412 => x"5a337a70",
         12413 => x"81055c33",
         12414 => x"717131ff",
         12415 => x"1b5b5842",
         12416 => x"4077802e",
         12417 => x"84913875",
         12418 => x"802ee138",
         12419 => x"933d7757",
         12420 => x"5a8359fc",
         12421 => x"83398158",
         12422 => x"fdc63980",
         12423 => x"e9173380",
         12424 => x"e8183371",
         12425 => x"882b0757",
         12426 => x"5575812e",
         12427 => x"098106f9",
         12428 => x"d538811b",
         12429 => x"58805ab4",
         12430 => x"1708782e",
         12431 => x"b1388317",
         12432 => x"335b7a7a",
         12433 => x"2e098106",
         12434 => x"829b3881",
         12435 => x"547753b8",
         12436 => x"17528117",
         12437 => x"3351ffb0",
         12438 => x"d23f84bb",
         12439 => x"8408802e",
         12440 => x"8538ff58",
         12441 => x"815a77b4",
         12442 => x"180c79f9",
         12443 => x"99387984",
         12444 => x"183484b7",
         12445 => x"173384b6",
         12446 => x"18337188",
         12447 => x"2b07575e",
         12448 => x"7582d4d5",
         12449 => x"2e098106",
         12450 => x"f8fc38b8",
         12451 => x"17831133",
         12452 => x"82123371",
         12453 => x"902b7188",
         12454 => x"2b078114",
         12455 => x"33707207",
         12456 => x"882b7533",
         12457 => x"71075e41",
         12458 => x"5945425c",
         12459 => x"5977848b",
         12460 => x"85a4d22e",
         12461 => x"098106f8",
         12462 => x"cd38849c",
         12463 => x"17831133",
         12464 => x"82123371",
         12465 => x"902b7188",
         12466 => x"2b078114",
         12467 => x"33707207",
         12468 => x"882b7533",
         12469 => x"71074744",
         12470 => x"405b5c5a",
         12471 => x"5e60868a",
         12472 => x"85e4f22e",
         12473 => x"098106f8",
         12474 => x"9d3884a0",
         12475 => x"17831133",
         12476 => x"82123371",
         12477 => x"902b7188",
         12478 => x"2b078114",
         12479 => x"33707207",
         12480 => x"882b7533",
         12481 => x"7107941e",
         12482 => x"0c5d84a4",
         12483 => x"1c831133",
         12484 => x"82123371",
         12485 => x"902b7188",
         12486 => x"2b078114",
         12487 => x"33707207",
         12488 => x"882b7533",
         12489 => x"71076290",
         12490 => x"050c5944",
         12491 => x"49465c45",
         12492 => x"40455b56",
         12493 => x"5a7c7734",
         12494 => x"84e2dc22",
         12495 => x"81055d7c",
         12496 => x"84e2dc23",
         12497 => x"7c861823",
         12498 => x"84e2e40b",
         12499 => x"8c180c80",
         12500 => x"0b98180c",
         12501 => x"f7cf397b",
         12502 => x"8324f8f0",
         12503 => x"387b7a7f",
         12504 => x"0c56f295",
         12505 => x"397554b4",
         12506 => x"170853b8",
         12507 => x"17705381",
         12508 => x"18335259",
         12509 => x"ffafb33f",
         12510 => x"84bb8408",
         12511 => x"7a2e0981",
         12512 => x"0681a438",
         12513 => x"84bb8408",
         12514 => x"831834b4",
         12515 => x"1708a818",
         12516 => x"0831407f",
         12517 => x"a0180827",
         12518 => x"8b388217",
         12519 => x"33416082",
         12520 => x"2e818d38",
         12521 => x"84bb8408",
         12522 => x"5afda039",
         12523 => x"74567480",
         12524 => x"2ef39138",
         12525 => x"850b818a",
         12526 => x"1883e6b8",
         12527 => x"5c5a58fc",
         12528 => x"ab3980e3",
         12529 => x"173380e2",
         12530 => x"18337188",
         12531 => x"2b075f5a",
         12532 => x"8d587df6",
         12533 => x"d2388817",
         12534 => x"224261f6",
         12535 => x"ca3880e4",
         12536 => x"17831133",
         12537 => x"82123371",
         12538 => x"902b7188",
         12539 => x"2b078114",
         12540 => x"33707207",
         12541 => x"882b7533",
         12542 => x"7107ac1e",
         12543 => x"0c5a7d82",
         12544 => x"2b5a4344",
         12545 => x"405940f5",
         12546 => x"d8397558",
         12547 => x"75802ef9",
         12548 => x"e8388258",
         12549 => x"f9e33975",
         12550 => x"802ef2a8",
         12551 => x"38933d77",
         12552 => x"575a8359",
         12553 => x"f7f23975",
         12554 => x"5a79f5da",
         12555 => x"38fcbf39",
         12556 => x"7554b417",
         12557 => x"08a01808",
         12558 => x"05537852",
         12559 => x"81173351",
         12560 => x"ffade73f",
         12561 => x"fc8539f0",
         12562 => x"3d0d0280",
         12563 => x"d3053364",
         12564 => x"7043933d",
         12565 => x"41575dff",
         12566 => x"765a4075",
         12567 => x"802e80e9",
         12568 => x"38787081",
         12569 => x"055a3370",
         12570 => x"9f265555",
         12571 => x"74ba2e80",
         12572 => x"e23873ed",
         12573 => x"3874ba2e",
         12574 => x"80d93884",
         12575 => x"e2e03354",
         12576 => x"80742480",
         12577 => x"c4387310",
         12578 => x"1084e2cc",
         12579 => x"05700855",
         12580 => x"5573802e",
         12581 => x"84388074",
         12582 => x"34625473",
         12583 => x"802e8638",
         12584 => x"80743462",
         12585 => x"5473750c",
         12586 => x"7c547c80",
         12587 => x"2e923880",
         12588 => x"53933d70",
         12589 => x"53840551",
         12590 => x"ef813f84",
         12591 => x"bb840854",
         12592 => x"7384bb84",
         12593 => x"0c923d0d",
         12594 => x"048b0b84",
         12595 => x"bb840c92",
         12596 => x"3d0d0475",
         12597 => x"33d01170",
         12598 => x"81ff0656",
         12599 => x"56577389",
         12600 => x"26913882",
         12601 => x"167781ff",
         12602 => x"06d0055c",
         12603 => x"5877792e",
         12604 => x"80f73880",
         12605 => x"7f0883e6",
         12606 => x"f45e5f5b",
         12607 => x"7b087e59",
         12608 => x"5a797081",
         12609 => x"055b3378",
         12610 => x"7081055a",
         12611 => x"33ff9f12",
         12612 => x"59575576",
         12613 => x"99268938",
         12614 => x"e0157081",
         12615 => x"ff065654",
         12616 => x"ff9f1657",
         12617 => x"76992689",
         12618 => x"38e01670",
         12619 => x"81ff0657",
         12620 => x"54743070",
         12621 => x"9f2a5854",
         12622 => x"74762e09",
         12623 => x"81068538",
         12624 => x"76ffbe38",
         12625 => x"77793270",
         12626 => x"30707207",
         12627 => x"9f2a7907",
         12628 => x"5c575479",
         12629 => x"802e9238",
         12630 => x"811b841d",
         12631 => x"5d5b837b",
         12632 => x"25ff9938",
         12633 => x"7f54fe98",
         12634 => x"397a8324",
         12635 => x"f7387a79",
         12636 => x"600c54fe",
         12637 => x"8b39e63d",
         12638 => x"0d6c0284",
         12639 => x"0580fb05",
         12640 => x"33565a89",
         12641 => x"5679802e",
         12642 => x"a63874bf",
         12643 => x"0670549d",
         12644 => x"3dcc0553",
         12645 => x"9e3d8405",
         12646 => x"5259ed9f",
         12647 => x"3f84bb84",
         12648 => x"085784bb",
         12649 => x"8408802e",
         12650 => x"8f38807a",
         12651 => x"0c765675",
         12652 => x"84bb840c",
         12653 => x"9c3d0d04",
         12654 => x"7e406d52",
         12655 => x"903d7052",
         12656 => x"5ce19a3f",
         12657 => x"84bb8408",
         12658 => x"5784bb84",
         12659 => x"08802e81",
         12660 => x"ba38789c",
         12661 => x"065d7c80",
         12662 => x"2e81ca38",
         12663 => x"76802e83",
         12664 => x"e0387684",
         12665 => x"2e84f238",
         12666 => x"78880759",
         12667 => x"76ffbb38",
         12668 => x"78832a81",
         12669 => x"06587780",
         12670 => x"2e81d138",
         12671 => x"669b1133",
         12672 => x"9a123371",
         12673 => x"882b0761",
         12674 => x"70334258",
         12675 => x"5d5e567d",
         12676 => x"832e8697",
         12677 => x"38800b8e",
         12678 => x"1734800b",
         12679 => x"8f1734a1",
         12680 => x"0b901734",
         12681 => x"80cc0b91",
         12682 => x"17346656",
         12683 => x"a00b8b17",
         12684 => x"347e6757",
         12685 => x"5e800b9a",
         12686 => x"1734800b",
         12687 => x"9b17347d",
         12688 => x"335d7c83",
         12689 => x"2e85d738",
         12690 => x"6658800b",
         12691 => x"9c193480",
         12692 => x"0b9d1934",
         12693 => x"800b9e19",
         12694 => x"34800b9f",
         12695 => x"19347e55",
         12696 => x"810b8316",
         12697 => x"347a802e",
         12698 => x"80e2387e",
         12699 => x"b411087c",
         12700 => x"7e085957",
         12701 => x"5f57817b",
         12702 => x"2789389c",
         12703 => x"16087b26",
         12704 => x"83ec3882",
         12705 => x"57807a0c",
         12706 => x"fea33902",
         12707 => x"80e70533",
         12708 => x"70982b5c",
         12709 => x"587a8025",
         12710 => x"feb83886",
         12711 => x"799c065e",
         12712 => x"577cfeb8",
         12713 => x"3876fe82",
         12714 => x"380280c2",
         12715 => x"05337084",
         12716 => x"2a81065d",
         12717 => x"567b82b0",
         12718 => x"3878812a",
         12719 => x"81065d7c",
         12720 => x"802e8938",
         12721 => x"75810658",
         12722 => x"77829538",
         12723 => x"78832a81",
         12724 => x"06567580",
         12725 => x"2e863878",
         12726 => x"80c00759",
         12727 => x"7eb41108",
         12728 => x"a01c0c67",
         12729 => x"a41c0c67",
         12730 => x"9b11339a",
         12731 => x"12337188",
         12732 => x"2b077333",
         12733 => x"405b4057",
         12734 => x"5b7b832e",
         12735 => x"81fb3877",
         12736 => x"881b0c9c",
         12737 => x"16831133",
         12738 => x"82123371",
         12739 => x"902b7188",
         12740 => x"2b078114",
         12741 => x"33707207",
         12742 => x"882b7533",
         12743 => x"7107608c",
         12744 => x"050c437f",
         12745 => x"7f0c4158",
         12746 => x"5e595686",
         12747 => x"1b22841b",
         12748 => x"2378901b",
         12749 => x"34800b91",
         12750 => x"1b34800b",
         12751 => x"9c1b0c80",
         12752 => x"0b941b0c",
         12753 => x"a81a5c84",
         12754 => x"807c5755",
         12755 => x"80767081",
         12756 => x"055834ff",
         12757 => x"155574f4",
         12758 => x"3878852a",
         12759 => x"81065978",
         12760 => x"802efcc9",
         12761 => x"388c1a08",
         12762 => x"5574802e",
         12763 => x"fcbf3874",
         12764 => x"941b0c8a",
         12765 => x"1b227089",
         12766 => x"2b881c08",
         12767 => x"77595a5a",
         12768 => x"5b763070",
         12769 => x"78078025",
         12770 => x"51557876",
         12771 => x"2783e738",
         12772 => x"81707606",
         12773 => x"5e5b7c80",
         12774 => x"2e83db38",
         12775 => x"77527951",
         12776 => x"ffacbb3f",
         12777 => x"84bb8408",
         12778 => x"5884bb84",
         12779 => x"08812683",
         12780 => x"38825784",
         12781 => x"bb8408ff",
         12782 => x"2eb63875",
         12783 => x"793156c1",
         12784 => x"390280c2",
         12785 => x"05339106",
         12786 => x"5e7d9538",
         12787 => x"78822a81",
         12788 => x"06557480",
         12789 => x"2efc9938",
         12790 => x"8857807a",
         12791 => x"0cfbce39",
         12792 => x"8757807a",
         12793 => x"0cfbc639",
         12794 => x"8457807a",
         12795 => x"0cfbbe39",
         12796 => x"7a767a31",
         12797 => x"5757ff89",
         12798 => x"39951633",
         12799 => x"94173371",
         12800 => x"982b7190",
         12801 => x"2b077a07",
         12802 => x"881d0c9c",
         12803 => x"18831133",
         12804 => x"82123371",
         12805 => x"902b7188",
         12806 => x"2b078114",
         12807 => x"33707207",
         12808 => x"882b7533",
         12809 => x"7107628c",
         12810 => x"050c4561",
         12811 => x"610c555a",
         12812 => x"545b585e",
         12813 => x"5c861b22",
         12814 => x"841b2378",
         12815 => x"901b3480",
         12816 => x"0b911b34",
         12817 => x"800b9c1b",
         12818 => x"0c800b94",
         12819 => x"1b0ca81a",
         12820 => x"5c84807c",
         12821 => x"5755fdf4",
         12822 => x"397b51cc",
         12823 => x"c23f84bb",
         12824 => x"84087988",
         12825 => x"075a5776",
         12826 => x"fac038fb",
         12827 => x"83397452",
         12828 => x"7b51ffaa",
         12829 => x"e93f84bb",
         12830 => x"84085d84",
         12831 => x"bb840880",
         12832 => x"2e80cb38",
         12833 => x"84bb8408",
         12834 => x"812efbf7",
         12835 => x"3884bb84",
         12836 => x"08ff2e82",
         12837 => x"b7388053",
         12838 => x"74527551",
         12839 => x"ffb1a03f",
         12840 => x"84bb8408",
         12841 => x"838f389c",
         12842 => x"1608fe11",
         12843 => x"94180859",
         12844 => x"56587675",
         12845 => x"27903881",
         12846 => x"1794170c",
         12847 => x"84163381",
         12848 => x"07557484",
         12849 => x"17347c55",
         12850 => x"777d26ff",
         12851 => x"a138807f",
         12852 => x"7f725f59",
         12853 => x"575db416",
         12854 => x"087e2eaf",
         12855 => x"38831633",
         12856 => x"58777d2e",
         12857 => x"09810681",
         12858 => x"eb388154",
         12859 => x"7d53b816",
         12860 => x"52811633",
         12861 => x"51ffa3b3",
         12862 => x"3f84bb84",
         12863 => x"08802e85",
         12864 => x"38ff5781",
         12865 => x"5c76b417",
         12866 => x"0c7e567b",
         12867 => x"ff1c9018",
         12868 => x"0c577b80",
         12869 => x"2efbb538",
         12870 => x"807a0cf9",
         12871 => x"9039800b",
         12872 => x"94173480",
         12873 => x"0b951734",
         12874 => x"fa9e3995",
         12875 => x"16339417",
         12876 => x"3371982b",
         12877 => x"71902b07",
         12878 => x"7d075d56",
         12879 => x"58800b8e",
         12880 => x"1734800b",
         12881 => x"8f1734a1",
         12882 => x"0b901734",
         12883 => x"80cc0b91",
         12884 => x"17346656",
         12885 => x"a00b8b17",
         12886 => x"347e6757",
         12887 => x"5e800b9a",
         12888 => x"1734800b",
         12889 => x"9b17347d",
         12890 => x"335d7c83",
         12891 => x"2e098106",
         12892 => x"f9d638ff",
         12893 => x"a9397798",
         12894 => x"1b0c76f8",
         12895 => x"ad387583",
         12896 => x"ff065978",
         12897 => x"802ef8a5",
         12898 => x"387efe19",
         12899 => x"9c1208fe",
         12900 => x"05405959",
         12901 => x"777e27f9",
         12902 => x"ea388a19",
         12903 => x"22787129",
         12904 => x"b01b0805",
         12905 => x"565b7480",
         12906 => x"2ef9d838",
         12907 => x"75892a15",
         12908 => x"709c1c0c",
         12909 => x"58815477",
         12910 => x"537b5281",
         12911 => x"193351ff",
         12912 => x"a1e93f84",
         12913 => x"bb840880",
         12914 => x"2ef7e238",
         12915 => x"8157807a",
         12916 => x"0cf7da39",
         12917 => x"8154b416",
         12918 => x"0853b816",
         12919 => x"70538117",
         12920 => x"335258ff",
         12921 => x"a2c43f84",
         12922 => x"bb84087d",
         12923 => x"2e098106",
         12924 => x"80ce3884",
         12925 => x"bb840883",
         12926 => x"1734b416",
         12927 => x"08a81708",
         12928 => x"3184bb84",
         12929 => x"085d5574",
         12930 => x"a0170827",
         12931 => x"fddc3882",
         12932 => x"16335574",
         12933 => x"822e0981",
         12934 => x"06fdcf38",
         12935 => x"8154b416",
         12936 => x"08a01708",
         12937 => x"05537752",
         12938 => x"81163351",
         12939 => x"ffa1fb3f",
         12940 => x"7c5cfdb6",
         12941 => x"3984bb84",
         12942 => x"0857807a",
         12943 => x"0cf6ee39",
         12944 => x"815cfdc5",
         12945 => x"39f23d0d",
         12946 => x"60636564",
         12947 => x"40405b59",
         12948 => x"807e0c89",
         12949 => x"5778802e",
         12950 => x"9f387808",
         12951 => x"5675802e",
         12952 => x"97387533",
         12953 => x"5574802e",
         12954 => x"8f388616",
         12955 => x"22841a22",
         12956 => x"595b7a78",
         12957 => x"2e83b438",
         12958 => x"8055745f",
         12959 => x"76557681",
         12960 => x"e7389119",
         12961 => x"33557481",
         12962 => x"df389019",
         12963 => x"33810657",
         12964 => x"87567680",
         12965 => x"2e81c838",
         12966 => x"9419088c",
         12967 => x"1a087131",
         12968 => x"56567975",
         12969 => x"2681ca38",
         12970 => x"79802e81",
         12971 => x"b0387583",
         12972 => x"ff065c7b",
         12973 => x"8299387e",
         12974 => x"8a1122ff",
         12975 => x"0577892a",
         12976 => x"065d587b",
         12977 => x"9b387582",
         12978 => x"d0388819",
         12979 => x"08558175",
         12980 => x"2783c338",
         12981 => x"74ff2e83",
         12982 => x"ae387498",
         12983 => x"1a0c7e58",
         12984 => x"981908fe",
         12985 => x"059c1908",
         12986 => x"fe055c57",
         12987 => x"767b2783",
         12988 => x"a5388a18",
         12989 => x"22707829",
         12990 => x"b01a0805",
         12991 => x"56567480",
         12992 => x"2e839338",
         12993 => x"7b157a89",
         12994 => x"2a5c577a",
         12995 => x"802e80e6",
         12996 => x"387a1c55",
         12997 => x"75752785",
         12998 => x"38757c31",
         12999 => x"5b7a5476",
         13000 => x"537c5281",
         13001 => x"183351ff",
         13002 => x"9f813f84",
         13003 => x"bb840882",
         13004 => x"d6389019",
         13005 => x"3370982b",
         13006 => x"59568078",
         13007 => x"24828738",
         13008 => x"7a892b57",
         13009 => x"7977317e",
         13010 => x"08187f0c",
         13011 => x"771e941b",
         13012 => x"08197059",
         13013 => x"941c0c5e",
         13014 => x"5a79fed2",
         13015 => x"38805675",
         13016 => x"84bb840c",
         13017 => x"903d0d04",
         13018 => x"7484bb84",
         13019 => x"0c903d0d",
         13020 => x"04745afe",
         13021 => x"b3399c19",
         13022 => x"08567577",
         13023 => x"2e80c838",
         13024 => x"90193370",
         13025 => x"982ba81b",
         13026 => x"525d5b7b",
         13027 => x"8025a338",
         13028 => x"81547553",
         13029 => x"7a528118",
         13030 => x"3351ff9f",
         13031 => x"8d3f84bb",
         13032 => x"840881e3",
         13033 => x"38901933",
         13034 => x"80ff0655",
         13035 => x"74901a34",
         13036 => x"7e588154",
         13037 => x"76537a52",
         13038 => x"81183351",
         13039 => x"ff9dec3f",
         13040 => x"84bb8408",
         13041 => x"81c13876",
         13042 => x"9c1a0c94",
         13043 => x"19085675",
         13044 => x"83ff0684",
         13045 => x"80713158",
         13046 => x"55797727",
         13047 => x"83387957",
         13048 => x"767d7a17",
         13049 => x"a8055759",
         13050 => x"5676802e",
         13051 => x"fed63874",
         13052 => x"70810556",
         13053 => x"33787081",
         13054 => x"055a34ff",
         13055 => x"16567580",
         13056 => x"2efec138",
         13057 => x"74708105",
         13058 => x"56337870",
         13059 => x"81055a34",
         13060 => x"ff165675",
         13061 => x"da38feac",
         13062 => x"39981908",
         13063 => x"527851ff",
         13064 => x"a3bc3f84",
         13065 => x"bb840855",
         13066 => x"fda43981",
         13067 => x"163351ff",
         13068 => x"9ca73f84",
         13069 => x"bb840881",
         13070 => x"065574fc",
         13071 => x"bb387479",
         13072 => x"085657fc",
         13073 => x"b5399c19",
         13074 => x"08773156",
         13075 => x"757b27fd",
         13076 => x"ef388480",
         13077 => x"7671291e",
         13078 => x"a81b5858",
         13079 => x"55757081",
         13080 => x"05573377",
         13081 => x"70810559",
         13082 => x"34ff1555",
         13083 => x"74802efd",
         13084 => x"cf387570",
         13085 => x"81055733",
         13086 => x"77708105",
         13087 => x"5934ff15",
         13088 => x"5574da38",
         13089 => x"fdba3981",
         13090 => x"0b911a34",
         13091 => x"810b84bb",
         13092 => x"840c903d",
         13093 => x"0d04820b",
         13094 => x"911a3482",
         13095 => x"0b84bb84",
         13096 => x"0c903d0d",
         13097 => x"04f13d0d",
         13098 => x"61646665",
         13099 => x"41415c59",
         13100 => x"807f0c89",
         13101 => x"5778802e",
         13102 => x"9f387808",
         13103 => x"5675802e",
         13104 => x"97387533",
         13105 => x"5574802e",
         13106 => x"8f388616",
         13107 => x"22841a22",
         13108 => x"595a7978",
         13109 => x"2e84a838",
         13110 => x"80557440",
         13111 => x"76557682",
         13112 => x"cc389119",
         13113 => x"33557482",
         13114 => x"c4389019",
         13115 => x"3370812a",
         13116 => x"81065858",
         13117 => x"87567680",
         13118 => x"2e82a938",
         13119 => x"9419087b",
         13120 => x"115d577b",
         13121 => x"77278438",
         13122 => x"76095b7a",
         13123 => x"802e8289",
         13124 => x"387683ff",
         13125 => x"065d7c82",
         13126 => x"cd387f8a",
         13127 => x"1122ff05",
         13128 => x"78892a06",
         13129 => x"5e587caa",
         13130 => x"387682f9",
         13131 => x"38881908",
         13132 => x"5574802e",
         13133 => x"838c3874",
         13134 => x"812e83ed",
         13135 => x"3874ff2e",
         13136 => x"83d83874",
         13137 => x"981a0c88",
         13138 => x"19088538",
         13139 => x"74881a0c",
         13140 => x"7f589019",
         13141 => x"3370982b",
         13142 => x"5b57807a",
         13143 => x"2482f938",
         13144 => x"981908fe",
         13145 => x"059c1908",
         13146 => x"fe055d57",
         13147 => x"767c2783",
         13148 => x"b8388a18",
         13149 => x"22707829",
         13150 => x"b01a0805",
         13151 => x"56567480",
         13152 => x"2e83a638",
         13153 => x"7c157b89",
         13154 => x"2a5b5c79",
         13155 => x"802e81a6",
         13156 => x"38791d55",
         13157 => x"75752785",
         13158 => x"38757d31",
         13159 => x"5a79547b",
         13160 => x"537d5281",
         13161 => x"183351ff",
         13162 => x"9b803f84",
         13163 => x"bb840882",
         13164 => x"e9389c19",
         13165 => x"087c3156",
         13166 => x"757a27ab",
         13167 => x"3884800b",
         13168 => x"a81a7772",
         13169 => x"29600558",
         13170 => x"58557570",
         13171 => x"81055733",
         13172 => x"77708105",
         13173 => x"5934ff15",
         13174 => x"5574ef38",
         13175 => x"90193380",
         13176 => x"ff065d7c",
         13177 => x"901a3479",
         13178 => x"892b587a",
         13179 => x"78317f08",
         13180 => x"19600c78",
         13181 => x"1f941b08",
         13182 => x"1a707194",
         13183 => x"1e0c8c1d",
         13184 => x"08595a58",
         13185 => x"5f5b7476",
         13186 => x"27833875",
         13187 => x"55748c1a",
         13188 => x"0c7afdfd",
         13189 => x"38901933",
         13190 => x"587780c0",
         13191 => x"075b7a90",
         13192 => x"1a348056",
         13193 => x"7584bb84",
         13194 => x"0c913d0d",
         13195 => x"047484bb",
         13196 => x"840c913d",
         13197 => x"0d049c19",
         13198 => x"087c2ea2",
         13199 => x"38941908",
         13200 => x"57768c1a",
         13201 => x"08279b38",
         13202 => x"81547b53",
         13203 => x"a8195281",
         13204 => x"183351ff",
         13205 => x"98d53f84",
         13206 => x"bb840881",
         13207 => x"bd389419",
         13208 => x"08577b9c",
         13209 => x"1a0c7683",
         13210 => x"ff068480",
         13211 => x"71315955",
         13212 => x"7a782783",
         13213 => x"387a5877",
         13214 => x"7916a805",
         13215 => x"7f595656",
         13216 => x"77802e93",
         13217 => x"38767081",
         13218 => x"05583375",
         13219 => x"70810557",
         13220 => x"34ff1656",
         13221 => x"75ef3890",
         13222 => x"1933ff80",
         13223 => x"075a7990",
         13224 => x"1a34fec7",
         13225 => x"39981908",
         13226 => x"527851ff",
         13227 => x"acef3f84",
         13228 => x"bb840855",
         13229 => x"84bb8408",
         13230 => x"fcfd3890",
         13231 => x"193358fe",
         13232 => x"d8397652",
         13233 => x"7851ffac",
         13234 => x"d43f84bb",
         13235 => x"84085584",
         13236 => x"bb8408fc",
         13237 => x"e238e439",
         13238 => x"81549c19",
         13239 => x"0853a819",
         13240 => x"52811833",
         13241 => x"51ff98c2",
         13242 => x"3f84bb84",
         13243 => x"08ac3890",
         13244 => x"193380ff",
         13245 => x"06567590",
         13246 => x"1a347f58",
         13247 => x"fce23981",
         13248 => x"163351ff",
         13249 => x"96d33f84",
         13250 => x"bb840881",
         13251 => x"065574fb",
         13252 => x"c7387479",
         13253 => x"085657fb",
         13254 => x"c139810b",
         13255 => x"911a3481",
         13256 => x"0b84bb84",
         13257 => x"0c913d0d",
         13258 => x"04820b91",
         13259 => x"1a34820b",
         13260 => x"84bb840c",
         13261 => x"913d0d04",
         13262 => x"f53d0d7d",
         13263 => x"58895777",
         13264 => x"802e9f38",
         13265 => x"77085675",
         13266 => x"802e9738",
         13267 => x"75335574",
         13268 => x"802e8f38",
         13269 => x"86162284",
         13270 => x"19225a5a",
         13271 => x"79792e83",
         13272 => x"d2388055",
         13273 => x"745c7656",
         13274 => x"7681ee38",
         13275 => x"90183370",
         13276 => x"862a8106",
         13277 => x"5c577a80",
         13278 => x"2e81de38",
         13279 => x"76982b56",
         13280 => x"80762483",
         13281 => x"c9387ba0",
         13282 => x"19085856",
         13283 => x"b4160877",
         13284 => x"2eb83880",
         13285 => x"0b831733",
         13286 => x"715b5c5a",
         13287 => x"7a7a2e09",
         13288 => x"810681c0",
         13289 => x"38815476",
         13290 => x"53b81652",
         13291 => x"81163351",
         13292 => x"ff95f83f",
         13293 => x"84bb8408",
         13294 => x"802e8538",
         13295 => x"ff578159",
         13296 => x"76b4170c",
         13297 => x"78567881",
         13298 => x"9038a418",
         13299 => x"088b1133",
         13300 => x"a0075657",
         13301 => x"748b1834",
         13302 => x"77088819",
         13303 => x"087083ff",
         13304 => x"ff065d5a",
         13305 => x"567a9a18",
         13306 => x"347a882a",
         13307 => x"5a799b18",
         13308 => x"349c1776",
         13309 => x"3396195c",
         13310 => x"565b7483",
         13311 => x"2e81c838",
         13312 => x"8c180855",
         13313 => x"747b3474",
         13314 => x"882a5b7a",
         13315 => x"9d183474",
         13316 => x"902a5675",
         13317 => x"9e183474",
         13318 => x"982a5978",
         13319 => x"9f183480",
         13320 => x"7a34800b",
         13321 => x"971834a1",
         13322 => x"0b981834",
         13323 => x"80cc0b99",
         13324 => x"1834800b",
         13325 => x"92183480",
         13326 => x"0b931834",
         13327 => x"7b5b810b",
         13328 => x"831c347b",
         13329 => x"51ff9895",
         13330 => x"3f84bb84",
         13331 => x"08901933",
         13332 => x"81bf065b",
         13333 => x"56799019",
         13334 => x"34755574",
         13335 => x"84bb840c",
         13336 => x"8d3d0d04",
         13337 => x"8154b416",
         13338 => x"0853b816",
         13339 => x"70538117",
         13340 => x"33525bff",
         13341 => x"95b43f81",
         13342 => x"5984bb84",
         13343 => x"087a2e09",
         13344 => x"8106fec0",
         13345 => x"3884bb84",
         13346 => x"08831734",
         13347 => x"b41608a8",
         13348 => x"17083184",
         13349 => x"bb84085a",
         13350 => x"5574a017",
         13351 => x"0827fe85",
         13352 => x"38821633",
         13353 => x"5574822e",
         13354 => x"098106fd",
         13355 => x"f8388154",
         13356 => x"b41608a0",
         13357 => x"17080553",
         13358 => x"7a528116",
         13359 => x"3351ff94",
         13360 => x"e93f7959",
         13361 => x"fddf3978",
         13362 => x"902a5574",
         13363 => x"94183474",
         13364 => x"882a5675",
         13365 => x"9518348c",
         13366 => x"18085574",
         13367 => x"7b347488",
         13368 => x"2a5b7a9d",
         13369 => x"18347490",
         13370 => x"2a56759e",
         13371 => x"18347498",
         13372 => x"2a59789f",
         13373 => x"1834807a",
         13374 => x"34800b97",
         13375 => x"1834a10b",
         13376 => x"98183480",
         13377 => x"cc0b9918",
         13378 => x"34800b92",
         13379 => x"1834800b",
         13380 => x"9318347b",
         13381 => x"5b810b83",
         13382 => x"1c347b51",
         13383 => x"ff96be3f",
         13384 => x"84bb8408",
         13385 => x"90193381",
         13386 => x"bf065b56",
         13387 => x"79901934",
         13388 => x"fea73981",
         13389 => x"163351ff",
         13390 => x"929f3f84",
         13391 => x"bb840881",
         13392 => x"065574fc",
         13393 => x"9d387478",
         13394 => x"085657fc",
         13395 => x"97398154",
         13396 => x"9c180853",
         13397 => x"a818527b",
         13398 => x"81113352",
         13399 => x"57ff93ca",
         13400 => x"3f815584",
         13401 => x"bb8408fd",
         13402 => x"f2389018",
         13403 => x"3380ff06",
         13404 => x"59789019",
         13405 => x"347ba019",
         13406 => x"085856b4",
         13407 => x"1608772e",
         13408 => x"098106fc",
         13409 => x"8e38fcc2",
         13410 => x"39f93d0d",
         13411 => x"79705255",
         13412 => x"fba63f84",
         13413 => x"bb840854",
         13414 => x"84bb8408",
         13415 => x"b1388956",
         13416 => x"74802e9e",
         13417 => x"38740853",
         13418 => x"72802e96",
         13419 => x"38723352",
         13420 => x"71802e8e",
         13421 => x"38861322",
         13422 => x"84162258",
         13423 => x"5271772e",
         13424 => x"96388052",
         13425 => x"71587554",
         13426 => x"75843875",
         13427 => x"750c7384",
         13428 => x"bb840c89",
         13429 => x"3d0d0481",
         13430 => x"133351ff",
         13431 => x"90fb3f84",
         13432 => x"bb840881",
         13433 => x"065372da",
         13434 => x"38737508",
         13435 => x"5356d539",
         13436 => x"f63d0dff",
         13437 => x"7d705b57",
         13438 => x"5b75802e",
         13439 => x"b2387570",
         13440 => x"81055733",
         13441 => x"709f2652",
         13442 => x"5271ba2e",
         13443 => x"ac3870ee",
         13444 => x"3871ba2e",
         13445 => x"a43884e2",
         13446 => x"e0335180",
         13447 => x"71249038",
         13448 => x"7084e2e0",
         13449 => x"34800b84",
         13450 => x"bb840c8c",
         13451 => x"3d0d048b",
         13452 => x"0b84bb84",
         13453 => x"0c8c3d0d",
         13454 => x"047833d0",
         13455 => x"117081ff",
         13456 => x"06535353",
         13457 => x"70892691",
         13458 => x"38821973",
         13459 => x"81ff06d0",
         13460 => x"05595473",
         13461 => x"762e80f5",
         13462 => x"38800b83",
         13463 => x"e6f45b58",
         13464 => x"79087956",
         13465 => x"57767081",
         13466 => x"05583375",
         13467 => x"70810557",
         13468 => x"33ff9f12",
         13469 => x"53545270",
         13470 => x"99268938",
         13471 => x"e0127081",
         13472 => x"ff065354",
         13473 => x"ff9f1351",
         13474 => x"70992689",
         13475 => x"38e01370",
         13476 => x"81ff0654",
         13477 => x"54713070",
         13478 => x"9f2a5551",
         13479 => x"71732e09",
         13480 => x"81068538",
         13481 => x"73ffbe38",
         13482 => x"74763270",
         13483 => x"30707207",
         13484 => x"9f2a7607",
         13485 => x"59525276",
         13486 => x"802e9238",
         13487 => x"8118841b",
         13488 => x"5b588378",
         13489 => x"25ff9938",
         13490 => x"7a51fecf",
         13491 => x"39778324",
         13492 => x"f7387776",
         13493 => x"5e51fec3",
         13494 => x"39ea3d0d",
         13495 => x"8053983d",
         13496 => x"cc055299",
         13497 => x"3d51d2d3",
         13498 => x"3f84bb84",
         13499 => x"085584bb",
         13500 => x"8408802e",
         13501 => x"8a387484",
         13502 => x"bb840c98",
         13503 => x"3d0d047a",
         13504 => x"5c685298",
         13505 => x"3dd00551",
         13506 => x"c6d33f84",
         13507 => x"bb840855",
         13508 => x"84bb8408",
         13509 => x"80c63802",
         13510 => x"80d70533",
         13511 => x"70982b58",
         13512 => x"5a807724",
         13513 => x"80e23802",
         13514 => x"b2053370",
         13515 => x"842a8106",
         13516 => x"57597580",
         13517 => x"2eb2387a",
         13518 => x"639b1133",
         13519 => x"9a123371",
         13520 => x"882b0773",
         13521 => x"335e5a5b",
         13522 => x"57587983",
         13523 => x"2ea43876",
         13524 => x"98190c74",
         13525 => x"84bb840c",
         13526 => x"983d0d04",
         13527 => x"84bb8408",
         13528 => x"842e0981",
         13529 => x"06ff8f38",
         13530 => x"850b84bb",
         13531 => x"840c983d",
         13532 => x"0d049516",
         13533 => x"33941733",
         13534 => x"71982b71",
         13535 => x"902b0779",
         13536 => x"07981b0c",
         13537 => x"5b54cc39",
         13538 => x"7a7e9812",
         13539 => x"0c587484",
         13540 => x"bb840c98",
         13541 => x"3d0d04ff",
         13542 => x"9e3d0d80",
         13543 => x"e63d0880",
         13544 => x"e63d085d",
         13545 => x"40807c34",
         13546 => x"805380e4",
         13547 => x"3dfdb405",
         13548 => x"5280e53d",
         13549 => x"51d1843f",
         13550 => x"84bb8408",
         13551 => x"5984bb84",
         13552 => x"0883c838",
         13553 => x"6080d93d",
         13554 => x"0c7f6198",
         13555 => x"110880dd",
         13556 => x"3d0c5880",
         13557 => x"db3d085b",
         13558 => x"5879802e",
         13559 => x"82cc3880",
         13560 => x"d83d983d",
         13561 => x"405ba052",
         13562 => x"7a51ffa5",
         13563 => x"e93f84bb",
         13564 => x"84085984",
         13565 => x"bb840883",
         13566 => x"92386080",
         13567 => x"df3d0858",
         13568 => x"56b41608",
         13569 => x"772eb138",
         13570 => x"84bb8408",
         13571 => x"8317335f",
         13572 => x"5d7d83c7",
         13573 => x"38815476",
         13574 => x"53b81652",
         13575 => x"81163351",
         13576 => x"ff8d883f",
         13577 => x"84bb8408",
         13578 => x"802e8538",
         13579 => x"ff578159",
         13580 => x"76b4170c",
         13581 => x"7882d438",
         13582 => x"80df3d08",
         13583 => x"9b11339a",
         13584 => x"12337188",
         13585 => x"2b076370",
         13586 => x"335d4059",
         13587 => x"56567883",
         13588 => x"2e82da38",
         13589 => x"7680db3d",
         13590 => x"0c80527a",
         13591 => x"51ffa4f6",
         13592 => x"3f84bb84",
         13593 => x"085984bb",
         13594 => x"8408829f",
         13595 => x"3880527a",
         13596 => x"51ffaab4",
         13597 => x"3f84bb84",
         13598 => x"085984bb",
         13599 => x"8408bb38",
         13600 => x"80df3d08",
         13601 => x"9b11339a",
         13602 => x"12337188",
         13603 => x"2b076370",
         13604 => x"33425859",
         13605 => x"5e567d83",
         13606 => x"2e81fd38",
         13607 => x"767a2ea4",
         13608 => x"3884bb84",
         13609 => x"08527a51",
         13610 => x"ffa6a13f",
         13611 => x"84bb8408",
         13612 => x"5984bb84",
         13613 => x"08802eff",
         13614 => x"b4387884",
         13615 => x"2e83d838",
         13616 => x"7881c838",
         13617 => x"80e43dfd",
         13618 => x"b805527a",
         13619 => x"51ffbec8",
         13620 => x"3f787f82",
         13621 => x"05335b57",
         13622 => x"79802e90",
         13623 => x"38821f56",
         13624 => x"81178117",
         13625 => x"70335f57",
         13626 => x"577cf538",
         13627 => x"81175675",
         13628 => x"78268195",
         13629 => x"3876802e",
         13630 => x"9c387e17",
         13631 => x"820556ff",
         13632 => x"1880e63d",
         13633 => x"0811ff19",
         13634 => x"ff195959",
         13635 => x"56587533",
         13636 => x"753476eb",
         13637 => x"38ff1880",
         13638 => x"e63d0811",
         13639 => x"5f58af7e",
         13640 => x"3480da3d",
         13641 => x"085a79fd",
         13642 => x"bd387760",
         13643 => x"2e828a38",
         13644 => x"800b84e2",
         13645 => x"e0337010",
         13646 => x"1083e6f4",
         13647 => x"05700870",
         13648 => x"33435959",
         13649 => x"5e5a7e7a",
         13650 => x"2e8d3881",
         13651 => x"1a701770",
         13652 => x"33575f5a",
         13653 => x"74f53882",
         13654 => x"1a5b7a78",
         13655 => x"26ab3880",
         13656 => x"57767a27",
         13657 => x"94387616",
         13658 => x"5f7e337c",
         13659 => x"7081055e",
         13660 => x"34811757",
         13661 => x"797726ee",
         13662 => x"38ba7c70",
         13663 => x"81055e34",
         13664 => x"76ff2e09",
         13665 => x"810681df",
         13666 => x"38915980",
         13667 => x"7c347884",
         13668 => x"bb840c80",
         13669 => x"e43d0d04",
         13670 => x"95163394",
         13671 => x"17337198",
         13672 => x"2b71902b",
         13673 => x"07790759",
         13674 => x"565efdf0",
         13675 => x"39951633",
         13676 => x"94173371",
         13677 => x"982b7190",
         13678 => x"2b077907",
         13679 => x"80dd3d0c",
         13680 => x"5a5d8052",
         13681 => x"7a51ffa2",
         13682 => x"8d3f84bb",
         13683 => x"84085984",
         13684 => x"bb840880",
         13685 => x"2efd9638",
         13686 => x"ffb13981",
         13687 => x"54b41608",
         13688 => x"53b81670",
         13689 => x"53811733",
         13690 => x"525eff8a",
         13691 => x"bd3f8159",
         13692 => x"84bb8408",
         13693 => x"fcbe3884",
         13694 => x"bb840883",
         13695 => x"1734b416",
         13696 => x"08a81708",
         13697 => x"3184bb84",
         13698 => x"085a5574",
         13699 => x"a0170827",
         13700 => x"fc833882",
         13701 => x"16335574",
         13702 => x"822e0981",
         13703 => x"06fbf638",
         13704 => x"8154b416",
         13705 => x"08a01708",
         13706 => x"05537d52",
         13707 => x"81163351",
         13708 => x"ff89f73f",
         13709 => x"7c59fbdd",
         13710 => x"39ff1880",
         13711 => x"e63d0811",
         13712 => x"5c58af7b",
         13713 => x"34800b84",
         13714 => x"e2e03370",
         13715 => x"101083e6",
         13716 => x"f4057008",
         13717 => x"70334359",
         13718 => x"595e5a7e",
         13719 => x"7a2e0981",
         13720 => x"06fde838",
         13721 => x"fdf13980",
         13722 => x"e53d0818",
         13723 => x"8119595a",
         13724 => x"79337c70",
         13725 => x"81055e34",
         13726 => x"776027fe",
         13727 => x"8e3880e5",
         13728 => x"3d081881",
         13729 => x"19595a79",
         13730 => x"337c7081",
         13731 => x"055e347f",
         13732 => x"7826d438",
         13733 => x"fdf53982",
         13734 => x"59807c34",
         13735 => x"7884bb84",
         13736 => x"0c80e43d",
         13737 => x"0d04f53d",
         13738 => x"0d7d7f5a",
         13739 => x"57895876",
         13740 => x"802e9f38",
         13741 => x"76085675",
         13742 => x"802e9738",
         13743 => x"75335574",
         13744 => x"802e8f38",
         13745 => x"86162284",
         13746 => x"18225b5b",
         13747 => x"7a7a2e83",
         13748 => x"ee388055",
         13749 => x"745c7755",
         13750 => x"7782fb38",
         13751 => x"91173355",
         13752 => x"7482f338",
         13753 => x"8c170858",
         13754 => x"78782682",
         13755 => x"f2389417",
         13756 => x"0856805a",
         13757 => x"787a2e83",
         13758 => x"85387b8a",
         13759 => x"11227089",
         13760 => x"2b525c58",
         13761 => x"757a2e82",
         13762 => x"fc387752",
         13763 => x"ff1951fd",
         13764 => x"bb933f84",
         13765 => x"bb8408ff",
         13766 => x"17795470",
         13767 => x"535755fd",
         13768 => x"bb833f84",
         13769 => x"bb840875",
         13770 => x"2682da38",
         13771 => x"77307606",
         13772 => x"7094190c",
         13773 => x"79713198",
         13774 => x"1908585a",
         13775 => x"5b75802e",
         13776 => x"81923877",
         13777 => x"792780d3",
         13778 => x"38787831",
         13779 => x"94180819",
         13780 => x"94190c90",
         13781 => x"18337081",
         13782 => x"2a810651",
         13783 => x"5c597a80",
         13784 => x"2e82cc38",
         13785 => x"75527651",
         13786 => x"ff9bb23f",
         13787 => x"84bb8408",
         13788 => x"5684bb84",
         13789 => x"08802e9e",
         13790 => x"3875ff2e",
         13791 => x"81d13881",
         13792 => x"76278382",
         13793 => x"387b5575",
         13794 => x"9c160827",
         13795 => x"82f83875",
         13796 => x"98180cff",
         13797 => x"ae3984bb",
         13798 => x"84085994",
         13799 => x"17081994",
         13800 => x"180c7883",
         13801 => x"ff065877",
         13802 => x"802ea938",
         13803 => x"7bfe179c",
         13804 => x"1208fe05",
         13805 => x"5c575875",
         13806 => x"7a2782ca",
         13807 => x"388a1822",
         13808 => x"767129b0",
         13809 => x"1a08057a",
         13810 => x"892a115c",
         13811 => x"5c557a80",
         13812 => x"2e82b338",
         13813 => x"8c170858",
         13814 => x"94170856",
         13815 => x"77762790",
         13816 => x"38758c18",
         13817 => x"0c901733",
         13818 => x"80c00759",
         13819 => x"78901834",
         13820 => x"7583ff06",
         13821 => x"5b7a802e",
         13822 => x"81ab389c",
         13823 => x"17085675",
         13824 => x"7a2e81a1",
         13825 => x"38901733",
         13826 => x"70982ba8",
         13827 => x"195a5659",
         13828 => x"748025a2",
         13829 => x"38815475",
         13830 => x"5377527b",
         13831 => x"81113352",
         13832 => x"56ff8686",
         13833 => x"3f84bb84",
         13834 => x"08a53890",
         13835 => x"173380ff",
         13836 => x"06557490",
         13837 => x"18348154",
         13838 => x"79537752",
         13839 => x"7b811133",
         13840 => x"5258ff84",
         13841 => x"e63f84bb",
         13842 => x"8408802e",
         13843 => x"80d33881",
         13844 => x"0b911834",
         13845 => x"81557484",
         13846 => x"bb840c8d",
         13847 => x"3d0d0490",
         13848 => x"17337081",
         13849 => x"2a810657",
         13850 => x"5a75fd82",
         13851 => x"38779418",
         13852 => x"08575980",
         13853 => x"5a787a2e",
         13854 => x"098106fc",
         13855 => x"fd387994",
         13856 => x"180cfed4",
         13857 => x"39800b94",
         13858 => x"180c8817",
         13859 => x"08567580",
         13860 => x"2e80c738",
         13861 => x"7598180c",
         13862 => x"75802efe",
         13863 => x"b738fda3",
         13864 => x"39799c18",
         13865 => x"0c800b84",
         13866 => x"bb840c8d",
         13867 => x"3d0d0475",
         13868 => x"527651ff",
         13869 => x"8aa83f84",
         13870 => x"bb840856",
         13871 => x"fdbb3981",
         13872 => x"163351ff",
         13873 => x"83933f84",
         13874 => x"bb840881",
         13875 => x"065574fc",
         13876 => x"81387477",
         13877 => x"085658fb",
         13878 => x"fb397552",
         13879 => x"7651ff98",
         13880 => x"bc3f84bb",
         13881 => x"84085684",
         13882 => x"bb840881",
         13883 => x"2e983884",
         13884 => x"bb8408ff",
         13885 => x"2efed838",
         13886 => x"84bb8408",
         13887 => x"88180c75",
         13888 => x"98180cff",
         13889 => x"9339820b",
         13890 => x"91183482",
         13891 => x"0b84bb84",
         13892 => x"0c8d3d0d",
         13893 => x"04f63d0d",
         13894 => x"7c568954",
         13895 => x"75802ea2",
         13896 => x"3880538c",
         13897 => x"3dfc0552",
         13898 => x"8d3d8405",
         13899 => x"51c68c3f",
         13900 => x"84bb8408",
         13901 => x"5584bb84",
         13902 => x"08802e8f",
         13903 => x"3880760c",
         13904 => x"74547384",
         13905 => x"bb840c8c",
         13906 => x"3d0d047a",
         13907 => x"760c7d52",
         13908 => x"7551ffba",
         13909 => x"883f84bb",
         13910 => x"84085584",
         13911 => x"bb840880",
         13912 => x"d138ab16",
         13913 => x"3370982b",
         13914 => x"59598078",
         13915 => x"24af3886",
         13916 => x"16337084",
         13917 => x"2a81065b",
         13918 => x"5479802e",
         13919 => x"80c5389c",
         13920 => x"16089b11",
         13921 => x"339a1233",
         13922 => x"71882b07",
         13923 => x"7d70335d",
         13924 => x"5d5a5557",
         13925 => x"78832eb3",
         13926 => x"38778817",
         13927 => x"0c7a5886",
         13928 => x"18228417",
         13929 => x"23745275",
         13930 => x"51ff9aaa",
         13931 => x"3f84bb84",
         13932 => x"08557484",
         13933 => x"2e8d3874",
         13934 => x"802eff84",
         13935 => x"3880760c",
         13936 => x"fefe3985",
         13937 => x"5580760c",
         13938 => x"fef63995",
         13939 => x"17339418",
         13940 => x"3371982b",
         13941 => x"71902b07",
         13942 => x"7a078819",
         13943 => x"0c5a5aff",
         13944 => x"bc39fa3d",
         13945 => x"0d785589",
         13946 => x"5474802e",
         13947 => x"9e387408",
         13948 => x"5372802e",
         13949 => x"96387233",
         13950 => x"5271802e",
         13951 => x"8e388613",
         13952 => x"22841622",
         13953 => x"57527176",
         13954 => x"2e943880",
         13955 => x"52715773",
         13956 => x"84387375",
         13957 => x"0c7384bb",
         13958 => x"840c883d",
         13959 => x"0d048113",
         13960 => x"3351ff80",
         13961 => x"b43f84bb",
         13962 => x"84088106",
         13963 => x"5271dc38",
         13964 => x"71750853",
         13965 => x"54d739f8",
         13966 => x"3d0d7a7c",
         13967 => x"58558956",
         13968 => x"74802e9f",
         13969 => x"38740854",
         13970 => x"73802e97",
         13971 => x"38733353",
         13972 => x"72802e8f",
         13973 => x"38861422",
         13974 => x"84162259",
         13975 => x"5372782e",
         13976 => x"81973880",
         13977 => x"53725975",
         13978 => x"537580c7",
         13979 => x"3876802e",
         13980 => x"80f33875",
         13981 => x"527451ff",
         13982 => x"9eae3f84",
         13983 => x"bb840853",
         13984 => x"84bb8408",
         13985 => x"842eb538",
         13986 => x"84bb8408",
         13987 => x"a6387652",
         13988 => x"7451ffb3",
         13989 => x"833f7252",
         13990 => x"7451ff9a",
         13991 => x"af3f84bb",
         13992 => x"84088432",
         13993 => x"70307072",
         13994 => x"079f2c84",
         13995 => x"bb840806",
         13996 => x"55575472",
         13997 => x"84bb840c",
         13998 => x"8a3d0d04",
         13999 => x"75775375",
         14000 => x"5253ffb2",
         14001 => x"d33f7252",
         14002 => x"7451ff99",
         14003 => x"ff3f84bb",
         14004 => x"84088432",
         14005 => x"70307072",
         14006 => x"079f2c84",
         14007 => x"bb840806",
         14008 => x"555754cf",
         14009 => x"39755274",
         14010 => x"51ff97ea",
         14011 => x"3f84bb84",
         14012 => x"0884bb84",
         14013 => x"0c8a3d0d",
         14014 => x"04811433",
         14015 => x"51fefed9",
         14016 => x"3f84bb84",
         14017 => x"08810653",
         14018 => x"72fed838",
         14019 => x"72750854",
         14020 => x"56fed239",
         14021 => x"ed3d0d66",
         14022 => x"57805389",
         14023 => x"3d705397",
         14024 => x"3d5256c2",
         14025 => x"963f84bb",
         14026 => x"84085584",
         14027 => x"bb840880",
         14028 => x"2e8a3874",
         14029 => x"84bb840c",
         14030 => x"953d0d04",
         14031 => x"65527551",
         14032 => x"ffb69a3f",
         14033 => x"84bb8408",
         14034 => x"5584bb84",
         14035 => x"08e53802",
         14036 => x"80cb0533",
         14037 => x"70982b55",
         14038 => x"58807424",
         14039 => x"97387680",
         14040 => x"2ed13876",
         14041 => x"527551ff",
         14042 => x"b1ae3f74",
         14043 => x"84bb840c",
         14044 => x"953d0d04",
         14045 => x"860b84bb",
         14046 => x"840c953d",
         14047 => x"0d04ed3d",
         14048 => x"0d666856",
         14049 => x"5f805395",
         14050 => x"3dec0552",
         14051 => x"963d51c1",
         14052 => x"aa3f84bb",
         14053 => x"84085a84",
         14054 => x"bb84089a",
         14055 => x"387f750c",
         14056 => x"74089c11",
         14057 => x"08fe1194",
         14058 => x"13085957",
         14059 => x"59577575",
         14060 => x"268d3875",
         14061 => x"7f0c7984",
         14062 => x"bb840c95",
         14063 => x"3d0d0484",
         14064 => x"bb840877",
         14065 => x"335a5b78",
         14066 => x"812e8293",
         14067 => x"3877a818",
         14068 => x"0884bb84",
         14069 => x"085a5d59",
         14070 => x"7780c138",
         14071 => x"7b811d71",
         14072 => x"5c5d56b4",
         14073 => x"1708762e",
         14074 => x"82ef3883",
         14075 => x"1733785f",
         14076 => x"5d7c818d",
         14077 => x"38815475",
         14078 => x"53b81752",
         14079 => x"81173351",
         14080 => x"fefda83f",
         14081 => x"84bb8408",
         14082 => x"802e8538",
         14083 => x"ff5a815e",
         14084 => x"79b4180c",
         14085 => x"7f7e5b57",
         14086 => x"7d80cc38",
         14087 => x"76335e7d",
         14088 => x"822e828d",
         14089 => x"387717b8",
         14090 => x"05831133",
         14091 => x"82123371",
         14092 => x"902b7188",
         14093 => x"2b078114",
         14094 => x"33707207",
         14095 => x"882b7533",
         14096 => x"7180ffff",
         14097 => x"fe800607",
         14098 => x"70307080",
         14099 => x"25630560",
         14100 => x"840583ff",
         14101 => x"0662ff05",
         14102 => x"43414353",
         14103 => x"54525358",
         14104 => x"405e5678",
         14105 => x"fef2387a",
         14106 => x"7f0c7a94",
         14107 => x"180c8417",
         14108 => x"33810758",
         14109 => x"77841834",
         14110 => x"7984bb84",
         14111 => x"0c953d0d",
         14112 => x"048154b4",
         14113 => x"170853b8",
         14114 => x"17705381",
         14115 => x"1833525d",
         14116 => x"fefd973f",
         14117 => x"815e84bb",
         14118 => x"8408fef8",
         14119 => x"3884bb84",
         14120 => x"08831834",
         14121 => x"b41708a8",
         14122 => x"18083184",
         14123 => x"bb84085f",
         14124 => x"5574a018",
         14125 => x"0827febd",
         14126 => x"38821733",
         14127 => x"5574822e",
         14128 => x"098106fe",
         14129 => x"b0388154",
         14130 => x"b41708a0",
         14131 => x"18080553",
         14132 => x"7c528117",
         14133 => x"3351fefc",
         14134 => x"d13f775e",
         14135 => x"fe973982",
         14136 => x"7742923d",
         14137 => x"59567552",
         14138 => x"7751ff81",
         14139 => x"f13f84bb",
         14140 => x"8408ff2e",
         14141 => x"80e83884",
         14142 => x"bb840881",
         14143 => x"2e80f738",
         14144 => x"84bb8408",
         14145 => x"307084bb",
         14146 => x"84080780",
         14147 => x"257c0581",
         14148 => x"18625a58",
         14149 => x"5c5c9c17",
         14150 => x"087626ca",
         14151 => x"387a7f0c",
         14152 => x"7a94180c",
         14153 => x"84173381",
         14154 => x"07587784",
         14155 => x"1834fec8",
         14156 => x"397717b8",
         14157 => x"05811133",
         14158 => x"71337188",
         14159 => x"2b077030",
         14160 => x"7080251f",
         14161 => x"821d83ff",
         14162 => x"06ff1f5f",
         14163 => x"5d5f595f",
         14164 => x"5f5578fd",
         14165 => x"8338fe8f",
         14166 => x"39775afd",
         14167 => x"bf398160",
         14168 => x"585a7a7f",
         14169 => x"0c7a9418",
         14170 => x"0c841733",
         14171 => x"81075877",
         14172 => x"841834fe",
         14173 => x"83398260",
         14174 => x"585ae739",
         14175 => x"f63d0d7c",
         14176 => x"58895777",
         14177 => x"802e9f38",
         14178 => x"77085675",
         14179 => x"802e9738",
         14180 => x"75335574",
         14181 => x"802e8f38",
         14182 => x"86162284",
         14183 => x"19225a5a",
         14184 => x"79792e82",
         14185 => x"81388055",
         14186 => x"745b7681",
         14187 => x"83389118",
         14188 => x"33577680",
         14189 => x"fb389018",
         14190 => x"3370812a",
         14191 => x"81065659",
         14192 => x"87567480",
         14193 => x"2e80eb38",
         14194 => x"94180855",
         14195 => x"748c1908",
         14196 => x"2780dd38",
         14197 => x"7481fb38",
         14198 => x"88180878",
         14199 => x"08585581",
         14200 => x"75278938",
         14201 => x"9c170875",
         14202 => x"2680d838",
         14203 => x"8257800b",
         14204 => x"88190c94",
         14205 => x"18088c19",
         14206 => x"0c7880c0",
         14207 => x"07557490",
         14208 => x"193476a8",
         14209 => x"3874982b",
         14210 => x"5a798025",
         14211 => x"a3388154",
         14212 => x"9c180853",
         14213 => x"a818527a",
         14214 => x"81113352",
         14215 => x"59fefa8a",
         14216 => x"3f84bb84",
         14217 => x"08802e83",
         14218 => x"90388157",
         14219 => x"76911934",
         14220 => x"76567584",
         14221 => x"bb840c8c",
         14222 => x"3d0d0479",
         14223 => x"55797927",
         14224 => x"80ff3874",
         14225 => x"527751fe",
         14226 => x"ff943f84",
         14227 => x"bb84085a",
         14228 => x"84bb8408",
         14229 => x"802e80e9",
         14230 => x"3884bb84",
         14231 => x"08812e82",
         14232 => x"e83884bb",
         14233 => x"8408ff2e",
         14234 => x"82f53880",
         14235 => x"53745276",
         14236 => x"51ff85cb",
         14237 => x"3f84bb84",
         14238 => x"0882d838",
         14239 => x"9c1708fe",
         14240 => x"11941908",
         14241 => x"58565975",
         14242 => x"7527ffaf",
         14243 => x"38811694",
         14244 => x"180c8417",
         14245 => x"33810755",
         14246 => x"74841834",
         14247 => x"7955787a",
         14248 => x"26ffa038",
         14249 => x"9c398116",
         14250 => x"3351fef7",
         14251 => x"ac3f84bb",
         14252 => x"84088106",
         14253 => x"5574fdee",
         14254 => x"38747808",
         14255 => x"5657fde8",
         14256 => x"39800b90",
         14257 => x"19335a55",
         14258 => x"7457800b",
         14259 => x"88190cfe",
         14260 => x"a2399818",
         14261 => x"08527751",
         14262 => x"fefe833f",
         14263 => x"84bb8408",
         14264 => x"ff2e81c2",
         14265 => x"3884bb84",
         14266 => x"08812e81",
         14267 => x"be387681",
         14268 => x"ae387a59",
         14269 => x"84bb8408",
         14270 => x"9c1a0827",
         14271 => x"81a13884",
         14272 => x"bb840898",
         14273 => x"19087908",
         14274 => x"59575581",
         14275 => x"0b84bb84",
         14276 => x"082781a1",
         14277 => x"3884bb84",
         14278 => x"089c1808",
         14279 => x"27819638",
         14280 => x"75802e97",
         14281 => x"38ff5375",
         14282 => x"527651ff",
         14283 => x"84913f84",
         14284 => x"bb840856",
         14285 => x"84bb8408",
         14286 => x"80e33874",
         14287 => x"527751fe",
         14288 => x"fd9c3f84",
         14289 => x"bb84085a",
         14290 => x"84bb8408",
         14291 => x"802e80cb",
         14292 => x"3884bb84",
         14293 => x"08812e80",
         14294 => x"dc3884bb",
         14295 => x"8408ff2e",
         14296 => x"818f3880",
         14297 => x"53745276",
         14298 => x"51ff83d3",
         14299 => x"3f84bb84",
         14300 => x"0880f638",
         14301 => x"9c1708fe",
         14302 => x"11941908",
         14303 => x"58565975",
         14304 => x"75279038",
         14305 => x"81169418",
         14306 => x"0c841733",
         14307 => x"81075574",
         14308 => x"84183479",
         14309 => x"55787a26",
         14310 => x"ffa13880",
         14311 => x"56755790",
         14312 => x"183359fc",
         14313 => x"ce398157",
         14314 => x"febb3982",
         14315 => x"0b901933",
         14316 => x"5a57fcbf",
         14317 => x"398257e7",
         14318 => x"39901833",
         14319 => x"80ff0655",
         14320 => x"74901934",
         14321 => x"7656fcea",
         14322 => x"39820b90",
         14323 => x"19335a55",
         14324 => x"fdf63984",
         14325 => x"bb840890",
         14326 => x"19335a55",
         14327 => x"fdea3981",
         14328 => x"0b901933",
         14329 => x"5a55fde0",
         14330 => x"3984bb84",
         14331 => x"0857ffaf",
         14332 => x"398157ff",
         14333 => x"aa39db3d",
         14334 => x"0d8253a7",
         14335 => x"3dff9c05",
         14336 => x"52a83d51",
         14337 => x"ffb8b43f",
         14338 => x"84bb8408",
         14339 => x"5684bb84",
         14340 => x"08802e8a",
         14341 => x"387584bb",
         14342 => x"840ca73d",
         14343 => x"0d047d4b",
         14344 => x"a83d0852",
         14345 => x"9b3d7052",
         14346 => x"59ffacb1",
         14347 => x"3f84bb84",
         14348 => x"085684bb",
         14349 => x"8408de38",
         14350 => x"02819305",
         14351 => x"3370852a",
         14352 => x"81065957",
         14353 => x"865677cd",
         14354 => x"3876982b",
         14355 => x"5b807b24",
         14356 => x"c4380280",
         14357 => x"ee053370",
         14358 => x"81065d57",
         14359 => x"87567bff",
         14360 => x"b4387da3",
         14361 => x"3d089b11",
         14362 => x"339a1233",
         14363 => x"71882b07",
         14364 => x"7333415e",
         14365 => x"5c57587c",
         14366 => x"832e80d5",
         14367 => x"3876842a",
         14368 => x"81065776",
         14369 => x"802e80ed",
         14370 => x"38875698",
         14371 => x"18087b2e",
         14372 => x"ff833877",
         14373 => x"5f7a4184",
         14374 => x"bb840852",
         14375 => x"8f3d7052",
         14376 => x"55ff8cb2",
         14377 => x"3f84bb84",
         14378 => x"085684bb",
         14379 => x"8408fee5",
         14380 => x"3884bb84",
         14381 => x"08527451",
         14382 => x"ff91ed3f",
         14383 => x"84bb8408",
         14384 => x"5684bb84",
         14385 => x"08a03887",
         14386 => x"0b84bb84",
         14387 => x"0ca73d0d",
         14388 => x"04951633",
         14389 => x"94173371",
         14390 => x"982b7190",
         14391 => x"2b077d07",
         14392 => x"5d5d5dff",
         14393 => x"983984bb",
         14394 => x"8408842e",
         14395 => x"883884bb",
         14396 => x"8408fea1",
         14397 => x"3878086f",
         14398 => x"a83d0857",
         14399 => x"5d5774ff",
         14400 => x"2e80d338",
         14401 => x"74527851",
         14402 => x"ff8bcb3f",
         14403 => x"84bb8408",
         14404 => x"5684bb84",
         14405 => x"08802ebe",
         14406 => x"38753070",
         14407 => x"77078025",
         14408 => x"565a7a80",
         14409 => x"2e9a3874",
         14410 => x"802e9538",
         14411 => x"7a790858",
         14412 => x"55817b27",
         14413 => x"89389c17",
         14414 => x"087b2681",
         14415 => x"fd388256",
         14416 => x"75fdd238",
         14417 => x"7d51fef6",
         14418 => x"943f84bb",
         14419 => x"840884bb",
         14420 => x"840ca73d",
         14421 => x"0d04b817",
         14422 => x"5d981908",
         14423 => x"56805ab4",
         14424 => x"1708762e",
         14425 => x"82b93883",
         14426 => x"17337a59",
         14427 => x"55747a2e",
         14428 => x"09810680",
         14429 => x"dd388154",
         14430 => x"7553b817",
         14431 => x"52811733",
         14432 => x"51fef2a7",
         14433 => x"3f84bb84",
         14434 => x"08802e85",
         14435 => x"38ff5681",
         14436 => x"5875b418",
         14437 => x"0c775677",
         14438 => x"ab389c19",
         14439 => x"0858e578",
         14440 => x"34810b83",
         14441 => x"18349019",
         14442 => x"087c27fe",
         14443 => x"ec388052",
         14444 => x"7851ff8c",
         14445 => x"973f84bb",
         14446 => x"84085684",
         14447 => x"bb840880",
         14448 => x"2eff9638",
         14449 => x"75842e09",
         14450 => x"8106fecd",
         14451 => x"388256fe",
         14452 => x"c8398154",
         14453 => x"b4170853",
         14454 => x"7c528117",
         14455 => x"3351fef2",
         14456 => x"c93f8158",
         14457 => x"84bb8408",
         14458 => x"7a2e0981",
         14459 => x"06ffa638",
         14460 => x"84bb8408",
         14461 => x"831834b4",
         14462 => x"1708a818",
         14463 => x"083184bb",
         14464 => x"84085955",
         14465 => x"74a01808",
         14466 => x"27feeb38",
         14467 => x"82173355",
         14468 => x"74822e09",
         14469 => x"8106fede",
         14470 => x"388154b4",
         14471 => x"1708a018",
         14472 => x"0805537c",
         14473 => x"52811733",
         14474 => x"51fef1fe",
         14475 => x"3f7958fe",
         14476 => x"c5397955",
         14477 => x"79782780",
         14478 => x"e1387452",
         14479 => x"7851fef7",
         14480 => x"9d3f84bb",
         14481 => x"84085a84",
         14482 => x"bb840880",
         14483 => x"2e80cb38",
         14484 => x"84bb8408",
         14485 => x"812efde6",
         14486 => x"3884bb84",
         14487 => x"08ff2e80",
         14488 => x"cb388053",
         14489 => x"74527651",
         14490 => x"fefdd43f",
         14491 => x"84bb8408",
         14492 => x"b3389c17",
         14493 => x"08fe1194",
         14494 => x"1908585c",
         14495 => x"58757b27",
         14496 => x"ffb03881",
         14497 => x"1694180c",
         14498 => x"84173381",
         14499 => x"075c7b84",
         14500 => x"18347955",
         14501 => x"777a26ff",
         14502 => x"a1388056",
         14503 => x"fda23979",
         14504 => x"56fdf739",
         14505 => x"84bb8408",
         14506 => x"56fd9539",
         14507 => x"8156fd90",
         14508 => x"39e33d0d",
         14509 => x"82539f3d",
         14510 => x"ffbc0552",
         14511 => x"a03d51ff",
         14512 => x"b2f93f84",
         14513 => x"bb840856",
         14514 => x"84bb8408",
         14515 => x"802e8a38",
         14516 => x"7584bb84",
         14517 => x"0c9f3d0d",
         14518 => x"047d436f",
         14519 => x"52933d70",
         14520 => x"525affa6",
         14521 => x"f83f84bb",
         14522 => x"84085684",
         14523 => x"bb84088b",
         14524 => x"38880b84",
         14525 => x"bb840c9f",
         14526 => x"3d0d0484",
         14527 => x"bb840884",
         14528 => x"2e098106",
         14529 => x"cb380280",
         14530 => x"f3053370",
         14531 => x"852a8106",
         14532 => x"56588656",
         14533 => x"74ffb938",
         14534 => x"7d5f7452",
         14535 => x"8f3d7052",
         14536 => x"5dff83f9",
         14537 => x"3f84bb84",
         14538 => x"0875575c",
         14539 => x"84bb8408",
         14540 => x"83388756",
         14541 => x"84bb8408",
         14542 => x"812e80f9",
         14543 => x"3884bb84",
         14544 => x"08ff2e81",
         14545 => x"cb387581",
         14546 => x"c9387d84",
         14547 => x"bb840883",
         14548 => x"12335d5a",
         14549 => x"577a80e2",
         14550 => x"38fe199c",
         14551 => x"1808fe05",
         14552 => x"5a56805b",
         14553 => x"7579278d",
         14554 => x"388a1722",
         14555 => x"767129b0",
         14556 => x"1908055c",
         14557 => x"587ab418",
         14558 => x"0cb81759",
         14559 => x"84807957",
         14560 => x"55807670",
         14561 => x"81055834",
         14562 => x"ff155574",
         14563 => x"f4387458",
         14564 => x"8a172255",
         14565 => x"77752781",
         14566 => x"f9388154",
         14567 => x"771b5378",
         14568 => x"52811733",
         14569 => x"51feef82",
         14570 => x"3f84bb84",
         14571 => x"0881df38",
         14572 => x"811858dc",
         14573 => x"398256ff",
         14574 => x"84398154",
         14575 => x"b4170853",
         14576 => x"b8177053",
         14577 => x"81183352",
         14578 => x"58feeede",
         14579 => x"3f815684",
         14580 => x"bb8408be",
         14581 => x"3884bb84",
         14582 => x"08831834",
         14583 => x"b41708a8",
         14584 => x"18083155",
         14585 => x"74a01808",
         14586 => x"27feee38",
         14587 => x"8217335b",
         14588 => x"7a822e09",
         14589 => x"8106fee1",
         14590 => x"387554b4",
         14591 => x"1708a018",
         14592 => x"08055377",
         14593 => x"52811733",
         14594 => x"51feee9e",
         14595 => x"3ffeca39",
         14596 => x"81567b7d",
         14597 => x"08585581",
         14598 => x"7c27fdb4",
         14599 => x"387b9c18",
         14600 => x"0827fdac",
         14601 => x"3874527c",
         14602 => x"51fef3b2",
         14603 => x"3f84bb84",
         14604 => x"085a84bb",
         14605 => x"8408802e",
         14606 => x"fd963884",
         14607 => x"bb840881",
         14608 => x"2efd8d38",
         14609 => x"84bb8408",
         14610 => x"ff2efd84",
         14611 => x"38805374",
         14612 => x"527651fe",
         14613 => x"f9e93f84",
         14614 => x"bb8408fc",
         14615 => x"f3389c17",
         14616 => x"08fe1194",
         14617 => x"19085a5c",
         14618 => x"59777b27",
         14619 => x"90388118",
         14620 => x"94180c84",
         14621 => x"17338107",
         14622 => x"5c7b8418",
         14623 => x"34795578",
         14624 => x"7a26ffa1",
         14625 => x"387584bb",
         14626 => x"840c9f3d",
         14627 => x"0d048a17",
         14628 => x"22557483",
         14629 => x"ffff0657",
         14630 => x"81567678",
         14631 => x"2e098106",
         14632 => x"fef0388b",
         14633 => x"0bb81f56",
         14634 => x"56a07570",
         14635 => x"81055734",
         14636 => x"ff165675",
         14637 => x"f4387d57",
         14638 => x"ae0bb818",
         14639 => x"347d5890",
         14640 => x"0b80c319",
         14641 => x"347d5975",
         14642 => x"80ce1a34",
         14643 => x"7580cf1a",
         14644 => x"34a10b80",
         14645 => x"d01a3480",
         14646 => x"cc0b80d1",
         14647 => x"1a347d7c",
         14648 => x"83ffff06",
         14649 => x"59567780",
         14650 => x"d2173477",
         14651 => x"882a5b7a",
         14652 => x"80d31734",
         14653 => x"75335574",
         14654 => x"832e81cc",
         14655 => x"387d59a0",
         14656 => x"0b80d81a",
         14657 => x"b81b5758",
         14658 => x"56747081",
         14659 => x"05563377",
         14660 => x"70810559",
         14661 => x"34ff1656",
         14662 => x"75ef387d",
         14663 => x"56ae0b80",
         14664 => x"d9173464",
         14665 => x"7e7183ff",
         14666 => x"ff065b57",
         14667 => x"577880f2",
         14668 => x"17347888",
         14669 => x"2a5b7a80",
         14670 => x"f3173475",
         14671 => x"33557483",
         14672 => x"2e80f038",
         14673 => x"7d5b810b",
         14674 => x"831c3479",
         14675 => x"51ff92cf",
         14676 => x"3f84bb84",
         14677 => x"085684bb",
         14678 => x"8408fdb6",
         14679 => x"38695684",
         14680 => x"bb840896",
         14681 => x"173484bb",
         14682 => x"84089717",
         14683 => x"34a10b98",
         14684 => x"173480cc",
         14685 => x"0b991734",
         14686 => x"7d6a585d",
         14687 => x"779a1834",
         14688 => x"77882a59",
         14689 => x"789b1834",
         14690 => x"7c335a79",
         14691 => x"832e80d9",
         14692 => x"38695590",
         14693 => x"0b8b1634",
         14694 => x"7d57810b",
         14695 => x"8318347d",
         14696 => x"51feedb9",
         14697 => x"3f84bb84",
         14698 => x"08567584",
         14699 => x"bb840c9f",
         14700 => x"3d0d0476",
         14701 => x"902a5574",
         14702 => x"80ec1734",
         14703 => x"74882a57",
         14704 => x"7680ed17",
         14705 => x"34fefd39",
         14706 => x"7b902a5b",
         14707 => x"7a80cc17",
         14708 => x"347a882a",
         14709 => x"557480cd",
         14710 => x"17347d59",
         14711 => x"a00b80d8",
         14712 => x"1ab81b57",
         14713 => x"5856fea1",
         14714 => x"397b902a",
         14715 => x"58779418",
         14716 => x"3477882a",
         14717 => x"5c7b9518",
         14718 => x"34695590",
         14719 => x"0b8b1634",
         14720 => x"7d57810b",
         14721 => x"8318347d",
         14722 => x"51feecd1",
         14723 => x"3f84bb84",
         14724 => x"0856ff96",
         14725 => x"39d13d0d",
         14726 => x"b33db43d",
         14727 => x"0870595b",
         14728 => x"5f79802e",
         14729 => x"9b387970",
         14730 => x"81055b33",
         14731 => x"709f2656",
         14732 => x"5675ba2e",
         14733 => x"81b83874",
         14734 => x"ed3875ba",
         14735 => x"2e81af38",
         14736 => x"8253b13d",
         14737 => x"fefc0552",
         14738 => x"b23d51ff",
         14739 => x"abed3f84",
         14740 => x"bb840856",
         14741 => x"84bb8408",
         14742 => x"802e8a38",
         14743 => x"7584bb84",
         14744 => x"0cb13d0d",
         14745 => x"047fa63d",
         14746 => x"0cb23d08",
         14747 => x"52a53d70",
         14748 => x"5259ff9f",
         14749 => x"e83f84bb",
         14750 => x"84085684",
         14751 => x"bb8408dc",
         14752 => x"380281bb",
         14753 => x"053381a0",
         14754 => x"065d8656",
         14755 => x"7cce38a0",
         14756 => x"0b923dae",
         14757 => x"3d085858",
         14758 => x"55757081",
         14759 => x"05573377",
         14760 => x"70810559",
         14761 => x"34ff1555",
         14762 => x"74ef3899",
         14763 => x"3d58b078",
         14764 => x"7a585855",
         14765 => x"75708105",
         14766 => x"57337770",
         14767 => x"81055934",
         14768 => x"ff155574",
         14769 => x"ef38b33d",
         14770 => x"08527751",
         14771 => x"ff9f8e3f",
         14772 => x"84bb8408",
         14773 => x"5684bb84",
         14774 => x"0885d838",
         14775 => x"6aa83d08",
         14776 => x"2e81cb38",
         14777 => x"880b84bb",
         14778 => x"840cb13d",
         14779 => x"0d047633",
         14780 => x"d0117081",
         14781 => x"ff065757",
         14782 => x"58748926",
         14783 => x"91388217",
         14784 => x"7881ff06",
         14785 => x"d0055d59",
         14786 => x"787a2e80",
         14787 => x"fa38807f",
         14788 => x"0883e6f4",
         14789 => x"7008725d",
         14790 => x"5e5f5f5c",
         14791 => x"7a708105",
         14792 => x"5c337970",
         14793 => x"81055b33",
         14794 => x"ff9f125a",
         14795 => x"58567799",
         14796 => x"268938e0",
         14797 => x"167081ff",
         14798 => x"065755ff",
         14799 => x"9f175877",
         14800 => x"99268938",
         14801 => x"e0177081",
         14802 => x"ff065855",
         14803 => x"7530709f",
         14804 => x"2a595575",
         14805 => x"772e0981",
         14806 => x"06853877",
         14807 => x"ffbe3878",
         14808 => x"7a327030",
         14809 => x"7072079f",
         14810 => x"2a7a075d",
         14811 => x"58557a80",
         14812 => x"2e953881",
         14813 => x"1c841e5e",
         14814 => x"5c7b8324",
         14815 => x"fdc2387c",
         14816 => x"087e5a5b",
         14817 => x"ff96397b",
         14818 => x"8324fdb4",
         14819 => x"38797f0c",
         14820 => x"8253b13d",
         14821 => x"fefc0552",
         14822 => x"b23d51ff",
         14823 => x"a99d3f84",
         14824 => x"bb840856",
         14825 => x"84bb8408",
         14826 => x"fdb238fd",
         14827 => x"b8396caa",
         14828 => x"3d082e09",
         14829 => x"8106feac",
         14830 => x"387751ff",
         14831 => x"8de13f84",
         14832 => x"bb840856",
         14833 => x"84bb8408",
         14834 => x"fd92386f",
         14835 => x"58930b8d",
         14836 => x"19028805",
         14837 => x"80cd0558",
         14838 => x"565a7570",
         14839 => x"81055733",
         14840 => x"75708105",
         14841 => x"5734ff1a",
         14842 => x"5a79ef38",
         14843 => x"0280cb05",
         14844 => x"338b1934",
         14845 => x"8b183370",
         14846 => x"842a8106",
         14847 => x"40567e89",
         14848 => x"3875a007",
         14849 => x"57768b19",
         14850 => x"347f5d81",
         14851 => x"0b831e34",
         14852 => x"8b183370",
         14853 => x"842a8106",
         14854 => x"575c7580",
         14855 => x"2e81c538",
         14856 => x"a73d086b",
         14857 => x"2e81bd38",
         14858 => x"7f9b1933",
         14859 => x"9a1a3371",
         14860 => x"882b0772",
         14861 => x"3341585c",
         14862 => x"577d832e",
         14863 => x"82e038fe",
         14864 => x"169c1808",
         14865 => x"fe055e56",
         14866 => x"757d2782",
         14867 => x"c7388a17",
         14868 => x"22767129",
         14869 => x"b0190805",
         14870 => x"575e7580",
         14871 => x"2e82b538",
         14872 => x"757a5d58",
         14873 => x"b4170876",
         14874 => x"2eaa3883",
         14875 => x"17335f7e",
         14876 => x"83bc3881",
         14877 => x"547553b8",
         14878 => x"17528117",
         14879 => x"3351fee4",
         14880 => x"aa3f84bb",
         14881 => x"8408802e",
         14882 => x"8538ff58",
         14883 => x"815c77b4",
         14884 => x"180c7f57",
         14885 => x"7b80d818",
         14886 => x"56567bfb",
         14887 => x"bf388115",
         14888 => x"335a79ae",
         14889 => x"2e098106",
         14890 => x"bb386a70",
         14891 => x"83ffff06",
         14892 => x"5d567b80",
         14893 => x"f218347b",
         14894 => x"882a5877",
         14895 => x"80f31834",
         14896 => x"76335b7a",
         14897 => x"832e0981",
         14898 => x"06933875",
         14899 => x"902a5e7d",
         14900 => x"80ec1834",
         14901 => x"7d882a56",
         14902 => x"7580ed18",
         14903 => x"347f5781",
         14904 => x"0b831834",
         14905 => x"7808aa3d",
         14906 => x"08b23d08",
         14907 => x"575c5674",
         14908 => x"ff2e9538",
         14909 => x"74527851",
         14910 => x"fefbdb3f",
         14911 => x"84bb8408",
         14912 => x"5584bb84",
         14913 => x"0880f538",
         14914 => x"b8165c98",
         14915 => x"19085780",
         14916 => x"5ab41608",
         14917 => x"772eb438",
         14918 => x"8316337a",
         14919 => x"595f7e7a",
         14920 => x"2e098106",
         14921 => x"81a83881",
         14922 => x"547653b8",
         14923 => x"16528116",
         14924 => x"3351fee2",
         14925 => x"f63f84bb",
         14926 => x"8408802e",
         14927 => x"8538ff57",
         14928 => x"815876b4",
         14929 => x"170c7755",
         14930 => x"77aa389c",
         14931 => x"19085ae5",
         14932 => x"7a34810b",
         14933 => x"83173490",
         14934 => x"19087b27",
         14935 => x"a5388052",
         14936 => x"7851fefc",
         14937 => x"e73f84bb",
         14938 => x"84085584",
         14939 => x"bb840880",
         14940 => x"2eff9838",
         14941 => x"82567484",
         14942 => x"2ef9e138",
         14943 => x"745674f9",
         14944 => x"db387f51",
         14945 => x"fee5d63f",
         14946 => x"84bb8408",
         14947 => x"84bb840c",
         14948 => x"b13d0d04",
         14949 => x"820b84bb",
         14950 => x"840cb13d",
         14951 => x"0d049518",
         14952 => x"33941933",
         14953 => x"71982b71",
         14954 => x"902b0778",
         14955 => x"0758565c",
         14956 => x"fd8d3984",
         14957 => x"bb840884",
         14958 => x"2efbfe38",
         14959 => x"84bb8408",
         14960 => x"802efea0",
         14961 => x"387584bb",
         14962 => x"840cb13d",
         14963 => x"0d048154",
         14964 => x"b4160853",
         14965 => x"7b528116",
         14966 => x"3351fee2",
         14967 => x"cd3f8158",
         14968 => x"84bb8408",
         14969 => x"7a2e0981",
         14970 => x"06fedb38",
         14971 => x"84bb8408",
         14972 => x"831734b4",
         14973 => x"1608a817",
         14974 => x"083184bb",
         14975 => x"84085955",
         14976 => x"74a01708",
         14977 => x"27fea038",
         14978 => x"8216335d",
         14979 => x"7c822e09",
         14980 => x"8106fe93",
         14981 => x"388154b4",
         14982 => x"1608a017",
         14983 => x"0805537b",
         14984 => x"52811633",
         14985 => x"51fee282",
         14986 => x"3f7958fd",
         14987 => x"fa398154",
         14988 => x"b4170853",
         14989 => x"b8177053",
         14990 => x"81183352",
         14991 => x"5bfee1ea",
         14992 => x"3f815c84",
         14993 => x"bb8408fc",
         14994 => x"c93884bb",
         14995 => x"84088318",
         14996 => x"34b41708",
         14997 => x"a8180831",
         14998 => x"84bb8408",
         14999 => x"5d5574a0",
         15000 => x"180827fc",
         15001 => x"8e388217",
         15002 => x"335d7c82",
         15003 => x"2e098106",
         15004 => x"fc813881",
         15005 => x"54b41708",
         15006 => x"a0180805",
         15007 => x"537a5281",
         15008 => x"173351fe",
         15009 => x"e1a43f79",
         15010 => x"5cfbe839",
         15011 => x"ec3d0d02",
         15012 => x"80df0533",
         15013 => x"02840580",
         15014 => x"e3053356",
         15015 => x"57825396",
         15016 => x"3dcc0552",
         15017 => x"973d51ff",
         15018 => x"a3913f84",
         15019 => x"bb840856",
         15020 => x"84bb8408",
         15021 => x"802e8a38",
         15022 => x"7584bb84",
         15023 => x"0c963d0d",
         15024 => x"04785a66",
         15025 => x"52963dd0",
         15026 => x"0551ff97",
         15027 => x"903f84bb",
         15028 => x"84085684",
         15029 => x"bb8408e0",
         15030 => x"380280cf",
         15031 => x"053381a0",
         15032 => x"06548656",
         15033 => x"73d23874",
         15034 => x"a7066171",
         15035 => x"098b1233",
         15036 => x"71067a74",
         15037 => x"06075156",
         15038 => x"5755738b",
         15039 => x"17347855",
         15040 => x"810b8316",
         15041 => x"347851fe",
         15042 => x"e2d33f84",
         15043 => x"bb840884",
         15044 => x"bb840c96",
         15045 => x"3d0d04ec",
         15046 => x"3d0d6757",
         15047 => x"8253963d",
         15048 => x"cc055297",
         15049 => x"3d51ffa2",
         15050 => x"923f84bb",
         15051 => x"84085584",
         15052 => x"bb840880",
         15053 => x"2e8a3874",
         15054 => x"84bb840c",
         15055 => x"963d0d04",
         15056 => x"785a6652",
         15057 => x"963dd005",
         15058 => x"51ff9691",
         15059 => x"3f84bb84",
         15060 => x"085584bb",
         15061 => x"8408e038",
         15062 => x"0280cf05",
         15063 => x"3381a006",
         15064 => x"56865575",
         15065 => x"d2386084",
         15066 => x"18228619",
         15067 => x"2271902b",
         15068 => x"07595956",
         15069 => x"76961734",
         15070 => x"76882a55",
         15071 => x"74971734",
         15072 => x"76902a58",
         15073 => x"77981734",
         15074 => x"76982a54",
         15075 => x"73991734",
         15076 => x"7857810b",
         15077 => x"83183478",
         15078 => x"51fee1c1",
         15079 => x"3f84bb84",
         15080 => x"0884bb84",
         15081 => x"0c963d0d",
         15082 => x"04e83d0d",
         15083 => x"6b6d5d5b",
         15084 => x"80539a3d",
         15085 => x"cc05529b",
         15086 => x"3d51ffa0",
         15087 => x"fe3f84bb",
         15088 => x"840884bb",
         15089 => x"84083070",
         15090 => x"84bb8408",
         15091 => x"07802551",
         15092 => x"56577a80",
         15093 => x"2e8b3881",
         15094 => x"7076065a",
         15095 => x"567881a4",
         15096 => x"38763070",
         15097 => x"78078025",
         15098 => x"565b7b80",
         15099 => x"2e818c38",
         15100 => x"81707606",
         15101 => x"5a587880",
         15102 => x"2e818038",
         15103 => x"7ca41108",
         15104 => x"5856805a",
         15105 => x"b4160877",
         15106 => x"2e82f638",
         15107 => x"8316337a",
         15108 => x"5a55747a",
         15109 => x"2e098106",
         15110 => x"81983881",
         15111 => x"547653b8",
         15112 => x"16528116",
         15113 => x"3351fedd",
         15114 => x"823f84bb",
         15115 => x"8408802e",
         15116 => x"8538ff57",
         15117 => x"815976b4",
         15118 => x"170c7857",
         15119 => x"78bd387c",
         15120 => x"70335658",
         15121 => x"80c35674",
         15122 => x"832e8b38",
         15123 => x"80e45674",
         15124 => x"842e8338",
         15125 => x"a7567518",
         15126 => x"b8058311",
         15127 => x"33821233",
         15128 => x"71902b71",
         15129 => x"882b0781",
         15130 => x"14337072",
         15131 => x"07882b75",
         15132 => x"33710762",
         15133 => x"0c5f5d5e",
         15134 => x"57595676",
         15135 => x"84bb840c",
         15136 => x"9a3d0d04",
         15137 => x"7c5e8040",
         15138 => x"80528e3d",
         15139 => x"705255fe",
         15140 => x"f4c43f84",
         15141 => x"bb840857",
         15142 => x"84bb8408",
         15143 => x"802e818d",
         15144 => x"3876842e",
         15145 => x"098106fe",
         15146 => x"b838807b",
         15147 => x"348057fe",
         15148 => x"b0397754",
         15149 => x"b4160853",
         15150 => x"b8167053",
         15151 => x"81173352",
         15152 => x"5bfedce6",
         15153 => x"3f775984",
         15154 => x"bb84087a",
         15155 => x"2e098106",
         15156 => x"fee83884",
         15157 => x"bb840883",
         15158 => x"1734b416",
         15159 => x"08a81708",
         15160 => x"3184bb84",
         15161 => x"085a5574",
         15162 => x"a0170827",
         15163 => x"fead3882",
         15164 => x"16335574",
         15165 => x"822e0981",
         15166 => x"06fea038",
         15167 => x"7754b416",
         15168 => x"08a01708",
         15169 => x"05537a52",
         15170 => x"81163351",
         15171 => x"fedc9b3f",
         15172 => x"79598154",
         15173 => x"7653b816",
         15174 => x"52811633",
         15175 => x"51fedb8b",
         15176 => x"3f84bb84",
         15177 => x"08802efe",
         15178 => x"8d38fe86",
         15179 => x"39755274",
         15180 => x"51fef8f4",
         15181 => x"3f84bb84",
         15182 => x"085784bb",
         15183 => x"8408fee1",
         15184 => x"3884bb84",
         15185 => x"0884bb84",
         15186 => x"08665c59",
         15187 => x"59791881",
         15188 => x"197c1b57",
         15189 => x"59567533",
         15190 => x"75348119",
         15191 => x"598a7827",
         15192 => x"ec388b70",
         15193 => x"1c575880",
         15194 => x"76347780",
         15195 => x"2efcf238",
         15196 => x"ff187b11",
         15197 => x"70335c57",
         15198 => x"5879a02e",
         15199 => x"ea38fce1",
         15200 => x"397957fd",
         15201 => x"ba39e13d",
         15202 => x"0d8253a1",
         15203 => x"3dffb405",
         15204 => x"52a23d51",
         15205 => x"ff9da43f",
         15206 => x"84bb8408",
         15207 => x"5684bb84",
         15208 => x"0882a638",
         15209 => x"8f3d5d8b",
         15210 => x"7d5755a0",
         15211 => x"76708105",
         15212 => x"5834ff15",
         15213 => x"5574f438",
         15214 => x"74a33d08",
         15215 => x"70337081",
         15216 => x"ff065b58",
         15217 => x"585a9f78",
         15218 => x"2781b738",
         15219 => x"a23d903d",
         15220 => x"5c5c7581",
         15221 => x"ff068118",
         15222 => x"57557481",
         15223 => x"f538757c",
         15224 => x"0c7483ff",
         15225 => x"ff2681ff",
         15226 => x"387451a1",
         15227 => x"953f83b5",
         15228 => x"5284bb84",
         15229 => x"08519fdc",
         15230 => x"3f84bb84",
         15231 => x"0883ffff",
         15232 => x"06577680",
         15233 => x"2e81e038",
         15234 => x"83e8940b",
         15235 => x"83e89433",
         15236 => x"7081ff06",
         15237 => x"5b565878",
         15238 => x"802e81d6",
         15239 => x"38745678",
         15240 => x"772e9938",
         15241 => x"81187033",
         15242 => x"7081ff06",
         15243 => x"57575874",
         15244 => x"802e8938",
         15245 => x"74772e09",
         15246 => x"8106e938",
         15247 => x"7581ff06",
         15248 => x"597881a3",
         15249 => x"3881ff77",
         15250 => x"2781f838",
         15251 => x"79892681",
         15252 => x"963881ff",
         15253 => x"77278f38",
         15254 => x"76882a55",
         15255 => x"747b7081",
         15256 => x"055d3481",
         15257 => x"1a5a767b",
         15258 => x"7081055d",
         15259 => x"34811aa3",
         15260 => x"3d087033",
         15261 => x"7081ff06",
         15262 => x"5b58585a",
         15263 => x"779f26fe",
         15264 => x"d1388f3d",
         15265 => x"33578656",
         15266 => x"7681e52e",
         15267 => x"bc387980",
         15268 => x"2e993802",
         15269 => x"b7055679",
         15270 => x"1670335c",
         15271 => x"5c7aa02e",
         15272 => x"09810687",
         15273 => x"38ff1a5a",
         15274 => x"79ed387d",
         15275 => x"45804780",
         15276 => x"52953d70",
         15277 => x"5256fef0",
         15278 => x"9d3f84bb",
         15279 => x"84085584",
         15280 => x"bb840880",
         15281 => x"2eb43874",
         15282 => x"567584bb",
         15283 => x"840ca13d",
         15284 => x"0d0483b5",
         15285 => x"5274519e",
         15286 => x"e73f84bb",
         15287 => x"840883ff",
         15288 => x"ff065574",
         15289 => x"fdf83886",
         15290 => x"567584bb",
         15291 => x"840ca13d",
         15292 => x"0d0483e8",
         15293 => x"943356fe",
         15294 => x"c3398152",
         15295 => x"7551fef5",
         15296 => x"a73f84bb",
         15297 => x"84085584",
         15298 => x"bb840880",
         15299 => x"c1387980",
         15300 => x"2e82c438",
         15301 => x"8b6c7e59",
         15302 => x"57557670",
         15303 => x"81055833",
         15304 => x"76708105",
         15305 => x"5834ff15",
         15306 => x"5574ef38",
         15307 => x"7d5d810b",
         15308 => x"831e347d",
         15309 => x"51fedaa5",
         15310 => x"3f84bb84",
         15311 => x"08557456",
         15312 => x"ff87398a",
         15313 => x"7a27fe8a",
         15314 => x"388656ff",
         15315 => x"9c3984bb",
         15316 => x"8408842e",
         15317 => x"098106fe",
         15318 => x"ee388055",
         15319 => x"79752efe",
         15320 => x"e6387508",
         15321 => x"75537652",
         15322 => x"58feeeea",
         15323 => x"3f84bb84",
         15324 => x"085784bb",
         15325 => x"8408752e",
         15326 => x"09810681",
         15327 => x"843884bb",
         15328 => x"8408b819",
         15329 => x"5c5a9816",
         15330 => x"08578059",
         15331 => x"b4180877",
         15332 => x"2eb23883",
         15333 => x"18335574",
         15334 => x"792e0981",
         15335 => x"0681d738",
         15336 => x"81547653",
         15337 => x"b8185281",
         15338 => x"183351fe",
         15339 => x"d5fd3f84",
         15340 => x"bb840880",
         15341 => x"2e8538ff",
         15342 => x"57815976",
         15343 => x"b4190c78",
         15344 => x"5778be38",
         15345 => x"789c1708",
         15346 => x"7033575a",
         15347 => x"577481e5",
         15348 => x"2e819e38",
         15349 => x"74307080",
         15350 => x"25780756",
         15351 => x"5c74802e",
         15352 => x"81d73881",
         15353 => x"1a5a7981",
         15354 => x"2ea53881",
         15355 => x"527551fe",
         15356 => x"efda3f84",
         15357 => x"bb840857",
         15358 => x"84bb8408",
         15359 => x"802eff86",
         15360 => x"38875576",
         15361 => x"842efdbf",
         15362 => x"38765576",
         15363 => x"fdb938a0",
         15364 => x"6c575580",
         15365 => x"76708105",
         15366 => x"5834ff15",
         15367 => x"5574f438",
         15368 => x"6b56880b",
         15369 => x"8b17348b",
         15370 => x"6c7e5957",
         15371 => x"55767081",
         15372 => x"05583376",
         15373 => x"70810558",
         15374 => x"34ff1555",
         15375 => x"74802efd",
         15376 => x"eb387670",
         15377 => x"81055833",
         15378 => x"76708105",
         15379 => x"5834ff15",
         15380 => x"5574da38",
         15381 => x"fdd6396b",
         15382 => x"5ae57a34",
         15383 => x"7d5d810b",
         15384 => x"831e347d",
         15385 => x"51fed7f5",
         15386 => x"3f84bb84",
         15387 => x"0855fdce",
         15388 => x"398157fe",
         15389 => x"df398154",
         15390 => x"b4180853",
         15391 => x"7a528118",
         15392 => x"3351fed5",
         15393 => x"a53f84bb",
         15394 => x"8408792e",
         15395 => x"09810680",
         15396 => x"c33884bb",
         15397 => x"84088319",
         15398 => x"34b41808",
         15399 => x"a8190831",
         15400 => x"5c7ba019",
         15401 => x"08278a38",
         15402 => x"82183355",
         15403 => x"74822eb1",
         15404 => x"3884bb84",
         15405 => x"0859fde8",
         15406 => x"39745a81",
         15407 => x"527551fe",
         15408 => x"ee8a3f84",
         15409 => x"bb840857",
         15410 => x"84bb8408",
         15411 => x"802efdb6",
         15412 => x"38feae39",
         15413 => x"81705859",
         15414 => x"78802efd",
         15415 => x"e738fea1",
         15416 => x"398154b4",
         15417 => x"1808a019",
         15418 => x"0805537a",
         15419 => x"52811833",
         15420 => x"51fed4b6",
         15421 => x"3ffda939",
         15422 => x"f23d0d60",
         15423 => x"62028805",
         15424 => x"80cb0533",
         15425 => x"5e5b5789",
         15426 => x"5676802e",
         15427 => x"9f387608",
         15428 => x"5574802e",
         15429 => x"97387433",
         15430 => x"5473802e",
         15431 => x"8f388615",
         15432 => x"22841822",
         15433 => x"59597878",
         15434 => x"2e81c238",
         15435 => x"8054735f",
         15436 => x"7581a538",
         15437 => x"91173356",
         15438 => x"75819d38",
         15439 => x"79802e81",
         15440 => x"a2388c17",
         15441 => x"08819c38",
         15442 => x"90173370",
         15443 => x"812a8106",
         15444 => x"565d7480",
         15445 => x"2e818c38",
         15446 => x"7e8a1122",
         15447 => x"70892b70",
         15448 => x"557c5457",
         15449 => x"5c59fd86",
         15450 => x"bc3fff15",
         15451 => x"7a067030",
         15452 => x"7072079f",
         15453 => x"2a84bb84",
         15454 => x"0805901c",
         15455 => x"08794253",
         15456 => x"5f555881",
         15457 => x"78278838",
         15458 => x"9c190878",
         15459 => x"26833882",
         15460 => x"58777856",
         15461 => x"5b805974",
         15462 => x"527651fe",
         15463 => x"d8c03f81",
         15464 => x"157f5555",
         15465 => x"9c140875",
         15466 => x"26833882",
         15467 => x"5584bb84",
         15468 => x"08812e81",
         15469 => x"dc3884bb",
         15470 => x"8408ff2e",
         15471 => x"81d83884",
         15472 => x"bb840881",
         15473 => x"c5388119",
         15474 => x"59787d2e",
         15475 => x"bb387478",
         15476 => x"2e098106",
         15477 => x"c2388756",
         15478 => x"75547384",
         15479 => x"bb840c90",
         15480 => x"3d0d0487",
         15481 => x"0b84bb84",
         15482 => x"0c903d0d",
         15483 => x"04811533",
         15484 => x"51fed0e5",
         15485 => x"3f84bb84",
         15486 => x"08810654",
         15487 => x"73fead38",
         15488 => x"73770855",
         15489 => x"56fea739",
         15490 => x"7b802e81",
         15491 => x"8e387a7d",
         15492 => x"56587c80",
         15493 => x"2eab3881",
         15494 => x"18547481",
         15495 => x"2e80e638",
         15496 => x"73537752",
         15497 => x"7e51fede",
         15498 => x"963f84bb",
         15499 => x"84085684",
         15500 => x"bb8408ff",
         15501 => x"a3387781",
         15502 => x"19ff1757",
         15503 => x"595e74d7",
         15504 => x"387e7e90",
         15505 => x"120c557b",
         15506 => x"802eff8c",
         15507 => x"387a8818",
         15508 => x"0c798c18",
         15509 => x"0c901733",
         15510 => x"80c0075c",
         15511 => x"7b901834",
         15512 => x"9c1508fe",
         15513 => x"05941608",
         15514 => x"585a767a",
         15515 => x"26fee938",
         15516 => x"767d3194",
         15517 => x"160c8415",
         15518 => x"3381075d",
         15519 => x"7c841634",
         15520 => x"7554fed6",
         15521 => x"39ff54ff",
         15522 => x"9739745b",
         15523 => x"8059febe",
         15524 => x"398254fe",
         15525 => x"c5398154",
         15526 => x"fec039ff",
         15527 => x"1b5effa1",
         15528 => x"3984bb90",
         15529 => x"08e33d0d",
         15530 => x"a33d08a5",
         15531 => x"3d080288",
         15532 => x"05818705",
         15533 => x"3344425f",
         15534 => x"ff0ba23d",
         15535 => x"08705f5b",
         15536 => x"4079802e",
         15537 => x"858a3879",
         15538 => x"7081055b",
         15539 => x"33709f26",
         15540 => x"565675ba",
         15541 => x"2e859b38",
         15542 => x"74ed3875",
         15543 => x"ba2e8592",
         15544 => x"3884e2e0",
         15545 => x"33568076",
         15546 => x"2484e538",
         15547 => x"75101084",
         15548 => x"e2cc0570",
         15549 => x"08565a74",
         15550 => x"802e8438",
         15551 => x"80753475",
         15552 => x"1684baf8",
         15553 => x"113384ba",
         15554 => x"f9123340",
         15555 => x"5b5d8152",
         15556 => x"7951fece",
         15557 => x"e23f84bb",
         15558 => x"840881ff",
         15559 => x"06708106",
         15560 => x"5d568357",
         15561 => x"7b84ab38",
         15562 => x"75822a81",
         15563 => x"06408a57",
         15564 => x"7f849f38",
         15565 => x"9f3dfc05",
         15566 => x"53835279",
         15567 => x"51fed0e9",
         15568 => x"3f84bb84",
         15569 => x"08849838",
         15570 => x"6d557480",
         15571 => x"2e849038",
         15572 => x"74828080",
         15573 => x"26848838",
         15574 => x"ff157506",
         15575 => x"557483ff",
         15576 => x"387e802e",
         15577 => x"88388480",
         15578 => x"7f2683f8",
         15579 => x"387e8180",
         15580 => x"0a2683f0",
         15581 => x"38ff1f7f",
         15582 => x"06557483",
         15583 => x"e7387e89",
         15584 => x"2aa63d08",
         15585 => x"892a7089",
         15586 => x"2b77594c",
         15587 => x"475b6080",
         15588 => x"2e85ab38",
         15589 => x"65307080",
         15590 => x"25770756",
         15591 => x"5f915774",
         15592 => x"83b0387d",
         15593 => x"802e84df",
         15594 => x"38815474",
         15595 => x"53605279",
         15596 => x"51fecdf7",
         15597 => x"3f815784",
         15598 => x"bb840883",
         15599 => x"95386083",
         15600 => x"ff053361",
         15601 => x"83fe0533",
         15602 => x"71882b07",
         15603 => x"59568e57",
         15604 => x"7782d4d5",
         15605 => x"2e098106",
         15606 => x"82f8387d",
         15607 => x"90296105",
         15608 => x"83b21133",
         15609 => x"44586280",
         15610 => x"2e82e738",
         15611 => x"83b61883",
         15612 => x"11338212",
         15613 => x"3371902b",
         15614 => x"71882b07",
         15615 => x"81143370",
         15616 => x"7207882b",
         15617 => x"75337107",
         15618 => x"83ba1f83",
         15619 => x"11338212",
         15620 => x"3371902b",
         15621 => x"71882b07",
         15622 => x"81143370",
         15623 => x"7207882b",
         15624 => x"75337107",
         15625 => x"5ca23d0c",
         15626 => x"42a33d0c",
         15627 => x"a33d0c44",
         15628 => x"4e544559",
         15629 => x"4f415a4b",
         15630 => x"784d8e57",
         15631 => x"80ff7927",
         15632 => x"82903893",
         15633 => x"577a8180",
         15634 => x"26828738",
         15635 => x"61812a70",
         15636 => x"81064549",
         15637 => x"63802e83",
         15638 => x"f9386187",
         15639 => x"06456482",
         15640 => x"2e893861",
         15641 => x"81064766",
         15642 => x"83f43883",
         15643 => x"6e70304a",
         15644 => x"46437a58",
         15645 => x"62832e8a",
         15646 => x"c2387aae",
         15647 => x"38788c2a",
         15648 => x"57810b83",
         15649 => x"e8a82256",
         15650 => x"5874802e",
         15651 => x"9d387477",
         15652 => x"26983883",
         15653 => x"e8a85677",
         15654 => x"10821770",
         15655 => x"22575758",
         15656 => x"74802e86",
         15657 => x"38767527",
         15658 => x"ee387752",
         15659 => x"7851fcff",
         15660 => x"f43f84bb",
         15661 => x"84081084",
         15662 => x"055584bb",
         15663 => x"84089ff5",
         15664 => x"26963881",
         15665 => x"0b84bb84",
         15666 => x"081084bb",
         15667 => x"84080571",
         15668 => x"11722a83",
         15669 => x"05574c43",
         15670 => x"83ff1589",
         15671 => x"2a5d815c",
         15672 => x"a0477b1f",
         15673 => x"7d116805",
         15674 => x"6611ff05",
         15675 => x"706b0672",
         15676 => x"31584e57",
         15677 => x"4462832e",
         15678 => x"89b83874",
         15679 => x"1d5d7790",
         15680 => x"29167060",
         15681 => x"31565774",
         15682 => x"792682f2",
         15683 => x"38787c31",
         15684 => x"7d317853",
         15685 => x"70683152",
         15686 => x"56fcff89",
         15687 => x"3f84bb84",
         15688 => x"08406283",
         15689 => x"2e89f638",
         15690 => x"62822e09",
         15691 => x"810682dd",
         15692 => x"3883fff5",
         15693 => x"0b84bb84",
         15694 => x"082782ac",
         15695 => x"387a89f9",
         15696 => x"38771855",
         15697 => x"7480c026",
         15698 => x"89ef3874",
         15699 => x"5bfea339",
         15700 => x"8b577684",
         15701 => x"bb840c9f",
         15702 => x"3d0d84bb",
         15703 => x"900c0481",
         15704 => x"4efbfe39",
         15705 => x"930b84bb",
         15706 => x"840c9f3d",
         15707 => x"0d84bb90",
         15708 => x"0c047c33",
         15709 => x"d0117081",
         15710 => x"ff065757",
         15711 => x"57748926",
         15712 => x"9138821d",
         15713 => x"7781ff06",
         15714 => x"d0055d58",
         15715 => x"777a2e81",
         15716 => x"b238800b",
         15717 => x"83e6f45f",
         15718 => x"5c7d087d",
         15719 => x"575b7a70",
         15720 => x"81055c33",
         15721 => x"76708105",
         15722 => x"5833ff9f",
         15723 => x"12455957",
         15724 => x"62992689",
         15725 => x"38e01770",
         15726 => x"81ff0658",
         15727 => x"44ff9f18",
         15728 => x"45649926",
         15729 => x"8938e018",
         15730 => x"7081ff06",
         15731 => x"59467630",
         15732 => x"709f2a5a",
         15733 => x"4776782e",
         15734 => x"09810685",
         15735 => x"3878ffbe",
         15736 => x"38757a32",
         15737 => x"70307072",
         15738 => x"079f2a7b",
         15739 => x"075d4a4a",
         15740 => x"7a802e80",
         15741 => x"ce38811c",
         15742 => x"841f5f5c",
         15743 => x"837c25ff",
         15744 => x"98387f56",
         15745 => x"f9e0399f",
         15746 => x"3df80553",
         15747 => x"81527951",
         15748 => x"fecb963f",
         15749 => x"815784bb",
         15750 => x"8408feb6",
         15751 => x"3861832a",
         15752 => x"770684bb",
         15753 => x"84084056",
         15754 => x"758338bf",
         15755 => x"5f6c558e",
         15756 => x"577e7526",
         15757 => x"fe9c3874",
         15758 => x"7f3159fb",
         15759 => x"fb398156",
         15760 => x"fad2397b",
         15761 => x"8324ffba",
         15762 => x"387b7aa3",
         15763 => x"3d0c56f9",
         15764 => x"95396181",
         15765 => x"06489357",
         15766 => x"67802efd",
         15767 => x"f538826e",
         15768 => x"70304a46",
         15769 => x"43fc8b39",
         15770 => x"84bb8408",
         15771 => x"9ff5269d",
         15772 => x"387a8b38",
         15773 => x"77185b81",
         15774 => x"807b27fb",
         15775 => x"f5388e57",
         15776 => x"7684bb84",
         15777 => x"0c9f3d0d",
         15778 => x"84bb900c",
         15779 => x"04805562",
         15780 => x"812e8699",
         15781 => x"389ff560",
         15782 => x"278b3874",
         15783 => x"81065b8e",
         15784 => x"577afdae",
         15785 => x"38848061",
         15786 => x"57558076",
         15787 => x"70810558",
         15788 => x"34ff1555",
         15789 => x"74f4388b",
         15790 => x"6183e6c0",
         15791 => x"59575576",
         15792 => x"70810558",
         15793 => x"33767081",
         15794 => x"055834ff",
         15795 => x"155574ef",
         15796 => x"38608b05",
         15797 => x"45746534",
         15798 => x"82618c05",
         15799 => x"3477618d",
         15800 => x"05347b83",
         15801 => x"ffff064b",
         15802 => x"6a618e05",
         15803 => x"346a882a",
         15804 => x"5c7b618f",
         15805 => x"05348161",
         15806 => x"90053462",
         15807 => x"83327030",
         15808 => x"5a488061",
         15809 => x"91053478",
         15810 => x"9e2a8206",
         15811 => x"49686192",
         15812 => x"05346c56",
         15813 => x"7583ffff",
         15814 => x"2686ad38",
         15815 => x"7583ffff",
         15816 => x"06557461",
         15817 => x"93053474",
         15818 => x"882a4c6b",
         15819 => x"61940534",
         15820 => x"f8619505",
         15821 => x"34bf6198",
         15822 => x"05348061",
         15823 => x"990534ff",
         15824 => x"619a0534",
         15825 => x"80619b05",
         15826 => x"347e619c",
         15827 => x"05347e88",
         15828 => x"2a486761",
         15829 => x"9d05347e",
         15830 => x"902a4c6b",
         15831 => x"619e0534",
         15832 => x"7e982a84",
         15833 => x"bb900c84",
         15834 => x"bb900861",
         15835 => x"9f053462",
         15836 => x"832e85f7",
         15837 => x"388061a7",
         15838 => x"05348061",
         15839 => x"a80534a1",
         15840 => x"61a90534",
         15841 => x"80cc61aa",
         15842 => x"05347c83",
         15843 => x"ffff0655",
         15844 => x"74619605",
         15845 => x"3474882a",
         15846 => x"4b6a6197",
         15847 => x"0534ff80",
         15848 => x"61a40534",
         15849 => x"a961a605",
         15850 => x"349361ab",
         15851 => x"0583e6cc",
         15852 => x"59575576",
         15853 => x"70810558",
         15854 => x"33767081",
         15855 => x"055834ff",
         15856 => x"155574ef",
         15857 => x"386083fe",
         15858 => x"054980d5",
         15859 => x"69346083",
         15860 => x"ff054bff",
         15861 => x"aa6b3481",
         15862 => x"547e5360",
         15863 => x"527951fe",
         15864 => x"c6c83f81",
         15865 => x"5784bb84",
         15866 => x"08fae738",
         15867 => x"60175c62",
         15868 => x"832e879c",
         15869 => x"38696157",
         15870 => x"55807670",
         15871 => x"81055834",
         15872 => x"ff155574",
         15873 => x"f4386375",
         15874 => x"415b6283",
         15875 => x"2e86c038",
         15876 => x"87fffff8",
         15877 => x"5762812e",
         15878 => x"8338f857",
         15879 => x"76613476",
         15880 => x"882a7c45",
         15881 => x"55746470",
         15882 => x"81054634",
         15883 => x"76902a59",
         15884 => x"78647081",
         15885 => x"05463476",
         15886 => x"982a5675",
         15887 => x"64347c57",
         15888 => x"65597666",
         15889 => x"26833876",
         15890 => x"5978547a",
         15891 => x"53605279",
         15892 => x"51fec5d6",
         15893 => x"3f84bb84",
         15894 => x"0885e638",
         15895 => x"84806157",
         15896 => x"55807670",
         15897 => x"81055834",
         15898 => x"ff155574",
         15899 => x"f438781b",
         15900 => x"777a3158",
         15901 => x"5b76c938",
         15902 => x"7f810540",
         15903 => x"7f802eff",
         15904 => x"89387756",
         15905 => x"62832e83",
         15906 => x"38665665",
         15907 => x"55756626",
         15908 => x"83387555",
         15909 => x"74547a53",
         15910 => x"60527951",
         15911 => x"fec58b3f",
         15912 => x"84bb8408",
         15913 => x"859b3874",
         15914 => x"1b767631",
         15915 => x"575b75db",
         15916 => x"388c5862",
         15917 => x"832e9338",
         15918 => x"86586c83",
         15919 => x"ffff268a",
         15920 => x"38845862",
         15921 => x"822e8338",
         15922 => x"81587d84",
         15923 => x"c1386183",
         15924 => x"2a81065e",
         15925 => x"7d81b338",
         15926 => x"84806156",
         15927 => x"59807570",
         15928 => x"81055734",
         15929 => x"ff195978",
         15930 => x"f43880d5",
         15931 => x"6934ffaa",
         15932 => x"6b346083",
         15933 => x"be054778",
         15934 => x"67348167",
         15935 => x"81053481",
         15936 => x"67820534",
         15937 => x"78678305",
         15938 => x"34776784",
         15939 => x"05346c43",
         15940 => x"80fdc152",
         15941 => x"621f51fc",
         15942 => x"f78b3ffe",
         15943 => x"67850534",
         15944 => x"84bb8408",
         15945 => x"822abf07",
         15946 => x"57766786",
         15947 => x"053484bb",
         15948 => x"84086787",
         15949 => x"05347e61",
         15950 => x"83c60534",
         15951 => x"676183c7",
         15952 => x"05346b61",
         15953 => x"83c80534",
         15954 => x"84bb9008",
         15955 => x"6183c905",
         15956 => x"34626183",
         15957 => x"ca053462",
         15958 => x"882a4564",
         15959 => x"6183cb05",
         15960 => x"3462902a",
         15961 => x"58776183",
         15962 => x"cc053462",
         15963 => x"982a5f7e",
         15964 => x"6183cd05",
         15965 => x"34815478",
         15966 => x"53605279",
         15967 => x"51fec3aa",
         15968 => x"3f815784",
         15969 => x"bb8408f7",
         15970 => x"c9388053",
         15971 => x"80527951",
         15972 => x"fec4963f",
         15973 => x"815784bb",
         15974 => x"8408f7b6",
         15975 => x"3884bb84",
         15976 => x"0884bb84",
         15977 => x"0c9f3d0d",
         15978 => x"84bb900c",
         15979 => x"046255f9",
         15980 => x"e439741c",
         15981 => x"6416455c",
         15982 => x"f6c4397a",
         15983 => x"ae387891",
         15984 => x"2a57810b",
         15985 => x"83e8b822",
         15986 => x"56587480",
         15987 => x"2e9d3874",
         15988 => x"77269838",
         15989 => x"83e8b856",
         15990 => x"77108217",
         15991 => x"70225757",
         15992 => x"5874802e",
         15993 => x"86387675",
         15994 => x"27ee3877",
         15995 => x"527851fc",
         15996 => x"f5b33f84",
         15997 => x"bb840810",
         15998 => x"10848705",
         15999 => x"70892a5e",
         16000 => x"5ca05c80",
         16001 => x"0b84bb84",
         16002 => x"08fc808a",
         16003 => x"055847fd",
         16004 => x"fff00a77",
         16005 => x"27f5cb38",
         16006 => x"8e57f8e4",
         16007 => x"3984bb84",
         16008 => x"0883fff5",
         16009 => x"26f8e638",
         16010 => x"7af8d338",
         16011 => x"77812a5b",
         16012 => x"7af4bf38",
         16013 => x"8e57f8c8",
         16014 => x"39688106",
         16015 => x"4463802e",
         16016 => x"f8af3883",
         16017 => x"43f4ab39",
         16018 => x"7561a005",
         16019 => x"3475882a",
         16020 => x"496861a1",
         16021 => x"05347590",
         16022 => x"2a5b7a61",
         16023 => x"a2053475",
         16024 => x"982a5776",
         16025 => x"61a30534",
         16026 => x"f9c63980",
         16027 => x"6180c305",
         16028 => x"34806180",
         16029 => x"c40534a1",
         16030 => x"6180c505",
         16031 => x"3480cc61",
         16032 => x"80c60534",
         16033 => x"7c61a405",
         16034 => x"347c882a",
         16035 => x"5c7b61a5",
         16036 => x"05347c90",
         16037 => x"2a597861",
         16038 => x"a605347c",
         16039 => x"982a5675",
         16040 => x"61a70534",
         16041 => x"8261ac05",
         16042 => x"348061ad",
         16043 => x"05348061",
         16044 => x"ae053480",
         16045 => x"61af0534",
         16046 => x"8161b005",
         16047 => x"348061b1",
         16048 => x"05348661",
         16049 => x"b2053480",
         16050 => x"61b30534",
         16051 => x"ff806180",
         16052 => x"c00534a9",
         16053 => x"6180c205",
         16054 => x"34936180",
         16055 => x"c70583e6",
         16056 => x"e0595755",
         16057 => x"76708105",
         16058 => x"58337670",
         16059 => x"81055834",
         16060 => x"ff155574",
         16061 => x"802ef9cd",
         16062 => x"38767081",
         16063 => x"05583376",
         16064 => x"70810558",
         16065 => x"34ff1555",
         16066 => x"74da38f9",
         16067 => x"b8398154",
         16068 => x"80536052",
         16069 => x"7951febf",
         16070 => x"923f8157",
         16071 => x"84bb8408",
         16072 => x"f4b0387d",
         16073 => x"90296105",
         16074 => x"42776283",
         16075 => x"b2053476",
         16076 => x"5484bb84",
         16077 => x"08536052",
         16078 => x"7951febf",
         16079 => x"ed3ffcc3",
         16080 => x"39810b84",
         16081 => x"bb840c9f",
         16082 => x"3d0d84bb",
         16083 => x"900c04f8",
         16084 => x"61347b4a",
         16085 => x"ff6a7081",
         16086 => x"054c34ff",
         16087 => x"6a708105",
         16088 => x"4c34ff6a",
         16089 => x"34ff6184",
         16090 => x"0534ff61",
         16091 => x"850534ff",
         16092 => x"61860534",
         16093 => x"ff618705",
         16094 => x"34ff6188",
         16095 => x"0534ff61",
         16096 => x"890534ff",
         16097 => x"618a0534",
         16098 => x"8f65347c",
         16099 => x"57f9b139",
         16100 => x"7654861f",
         16101 => x"53605279",
         16102 => x"51febf8e",
         16103 => x"3f848061",
         16104 => x"56578075",
         16105 => x"70810557",
         16106 => x"34ff1757",
         16107 => x"76f43860",
         16108 => x"5c80d27c",
         16109 => x"7081055e",
         16110 => x"347b5580",
         16111 => x"d2757081",
         16112 => x"05573480",
         16113 => x"e1757081",
         16114 => x"05573480",
         16115 => x"c1753480",
         16116 => x"f26183e4",
         16117 => x"053480f2",
         16118 => x"6183e505",
         16119 => x"3480c161",
         16120 => x"83e60534",
         16121 => x"80e16183",
         16122 => x"e705347f",
         16123 => x"ff055b7a",
         16124 => x"6183e805",
         16125 => x"347a882a",
         16126 => x"59786183",
         16127 => x"e905347a",
         16128 => x"902a5675",
         16129 => x"6183ea05",
         16130 => x"347a982a",
         16131 => x"407f6183",
         16132 => x"eb053482",
         16133 => x"6183ec05",
         16134 => x"34766183",
         16135 => x"ed053476",
         16136 => x"6183ee05",
         16137 => x"34766183",
         16138 => x"ef053480",
         16139 => x"d56934ff",
         16140 => x"aa6b3481",
         16141 => x"54871f53",
         16142 => x"60527951",
         16143 => x"febdeb3f",
         16144 => x"8154811f",
         16145 => x"53605279",
         16146 => x"51febdde",
         16147 => x"3f696157",
         16148 => x"55f7a639",
         16149 => x"f43d0d7e",
         16150 => x"615b5b80",
         16151 => x"7b61ff05",
         16152 => x"5a575776",
         16153 => x"7825b838",
         16154 => x"8d3d598e",
         16155 => x"3df80554",
         16156 => x"81537852",
         16157 => x"7951ff9b",
         16158 => x"cc3f7b81",
         16159 => x"2e098106",
         16160 => x"9e388d3d",
         16161 => x"3355748d",
         16162 => x"2e903874",
         16163 => x"76708105",
         16164 => x"58348117",
         16165 => x"57748a2e",
         16166 => x"86387777",
         16167 => x"24cd3880",
         16168 => x"76347a55",
         16169 => x"76833876",
         16170 => x"557484bb",
         16171 => x"840c8e3d",
         16172 => x"0d04f73d",
         16173 => x"0d7b0284",
         16174 => x"05b30533",
         16175 => x"5957778a",
         16176 => x"2e80d538",
         16177 => x"84170856",
         16178 => x"8076249e",
         16179 => x"38881708",
         16180 => x"77178c05",
         16181 => x"56597775",
         16182 => x"34811655",
         16183 => x"74bb248e",
         16184 => x"38748418",
         16185 => x"0c811988",
         16186 => x"180c8b3d",
         16187 => x"0d048b3d",
         16188 => x"fc055474",
         16189 => x"538c1752",
         16190 => x"760851ff",
         16191 => x"9fa73f74",
         16192 => x"7a327030",
         16193 => x"7072079f",
         16194 => x"2a703084",
         16195 => x"1b0c811c",
         16196 => x"881b0c5a",
         16197 => x"5656d339",
         16198 => x"8d527651",
         16199 => x"ff943fff",
         16200 => x"a339e33d",
         16201 => x"0d0280ff",
         16202 => x"05338d3d",
         16203 => x"585880cc",
         16204 => x"77575580",
         16205 => x"76708105",
         16206 => x"5834ff15",
         16207 => x"5574f438",
         16208 => x"a13d0877",
         16209 => x"0c778a2e",
         16210 => x"80f7387c",
         16211 => x"56807624",
         16212 => x"80c0387d",
         16213 => x"77178c05",
         16214 => x"56597775",
         16215 => x"34811655",
         16216 => x"74bb24b8",
         16217 => x"38748418",
         16218 => x"0c811988",
         16219 => x"180c7c55",
         16220 => x"8075249e",
         16221 => x"389f3dff",
         16222 => x"ac115575",
         16223 => x"54c00552",
         16224 => x"760851ff",
         16225 => x"9e9f3f84",
         16226 => x"bb840886",
         16227 => x"387c7a2e",
         16228 => x"ba38ff0b",
         16229 => x"84bb840c",
         16230 => x"9f3d0d04",
         16231 => x"9f3dffb0",
         16232 => x"11557554",
         16233 => x"c0055276",
         16234 => x"0851ff9d",
         16235 => x"f83f747b",
         16236 => x"32703070",
         16237 => x"72079f2a",
         16238 => x"7030525a",
         16239 => x"5656ffa5",
         16240 => x"398d5276",
         16241 => x"51fdeb3f",
         16242 => x"ff81397d",
         16243 => x"84bb840c",
         16244 => x"9f3d0d04",
         16245 => x"fd3d0d75",
         16246 => x"0284059a",
         16247 => x"05225253",
         16248 => x"80527280",
         16249 => x"ff269038",
         16250 => x"7283ffff",
         16251 => x"06527184",
         16252 => x"bb840c85",
         16253 => x"3d0d0483",
         16254 => x"ffff7327",
         16255 => x"547083b5",
         16256 => x"2e098106",
         16257 => x"e9387380",
         16258 => x"2ee43883",
         16259 => x"e8c82251",
         16260 => x"72712e9c",
         16261 => x"38811270",
         16262 => x"83ffff06",
         16263 => x"53547180",
         16264 => x"ff268d38",
         16265 => x"711083e8",
         16266 => x"c8057022",
         16267 => x"5151e139",
         16268 => x"81801270",
         16269 => x"81ff0684",
         16270 => x"bb840c53",
         16271 => x"853d0d04",
         16272 => x"fe3d0d02",
         16273 => x"92052202",
         16274 => x"84059605",
         16275 => x"22535180",
         16276 => x"537080ff",
         16277 => x"268c3870",
         16278 => x"537284bb",
         16279 => x"840c843d",
         16280 => x"0d047183",
         16281 => x"b52e0981",
         16282 => x"06ef3870",
         16283 => x"81ff26e9",
         16284 => x"38701083",
         16285 => x"e6c80570",
         16286 => x"2284bb84",
         16287 => x"0c51843d",
         16288 => x"0d04fb3d",
         16289 => x"0d775170",
         16290 => x"83ffff26",
         16291 => x"80e13870",
         16292 => x"83ffff06",
         16293 => x"83eac856",
         16294 => x"56759fff",
         16295 => x"2680d938",
         16296 => x"74708205",
         16297 => x"56227571",
         16298 => x"30708025",
         16299 => x"737a2607",
         16300 => x"54565353",
         16301 => x"70b73871",
         16302 => x"70820553",
         16303 => x"22727188",
         16304 => x"2a545681",
         16305 => x"ff067014",
         16306 => x"52547076",
         16307 => x"24b13871",
         16308 => x"cf387310",
         16309 => x"15707082",
         16310 => x"05522254",
         16311 => x"73307080",
         16312 => x"25757926",
         16313 => x"07535552",
         16314 => x"70802ecb",
         16315 => x"38755170",
         16316 => x"84bb840c",
         16317 => x"873d0d04",
         16318 => x"83eebc55",
         16319 => x"ffa23971",
         16320 => x"8826ea38",
         16321 => x"71101083",
         16322 => x"caf00554",
         16323 => x"730804c7",
         16324 => x"a0167083",
         16325 => x"ffff0657",
         16326 => x"517551d3",
         16327 => x"39ffb016",
         16328 => x"7083ffff",
         16329 => x"065751f1",
         16330 => x"39881670",
         16331 => x"83ffff06",
         16332 => x"5751e639",
         16333 => x"e6167083",
         16334 => x"ffff0657",
         16335 => x"51db39d0",
         16336 => x"167083ff",
         16337 => x"ff065751",
         16338 => x"d039e016",
         16339 => x"7083ffff",
         16340 => x"065751c5",
         16341 => x"39f01670",
         16342 => x"83ffff06",
         16343 => x"5751ffb9",
         16344 => x"39757331",
         16345 => x"81067671",
         16346 => x"317083ff",
         16347 => x"ff065852",
         16348 => x"55ffa639",
         16349 => x"75733110",
         16350 => x"75057022",
         16351 => x"5252feef",
         16352 => x"39000000",
         16353 => x"00ffffff",
         16354 => x"ff00ffff",
         16355 => x"ffff00ff",
         16356 => x"ffffff00",
         16357 => x"0000198b",
         16358 => x"00001980",
         16359 => x"00001975",
         16360 => x"0000196a",
         16361 => x"0000195f",
         16362 => x"00001954",
         16363 => x"00001949",
         16364 => x"0000193e",
         16365 => x"00001933",
         16366 => x"00001928",
         16367 => x"0000191d",
         16368 => x"00001912",
         16369 => x"00001907",
         16370 => x"000018fc",
         16371 => x"000018f1",
         16372 => x"000018e6",
         16373 => x"000018db",
         16374 => x"000018d0",
         16375 => x"000018c5",
         16376 => x"000018ba",
         16377 => x"00001eca",
         16378 => x"00001f64",
         16379 => x"00001f64",
         16380 => x"00001f64",
         16381 => x"00001f64",
         16382 => x"00001f64",
         16383 => x"00001f64",
         16384 => x"00001f64",
         16385 => x"00001f64",
         16386 => x"00001f64",
         16387 => x"00001f64",
         16388 => x"00001f64",
         16389 => x"00001f64",
         16390 => x"00001f64",
         16391 => x"00001f64",
         16392 => x"00001f64",
         16393 => x"00001f64",
         16394 => x"00001f64",
         16395 => x"00001f64",
         16396 => x"00001f64",
         16397 => x"00001f64",
         16398 => x"00001f64",
         16399 => x"00001f64",
         16400 => x"00001f64",
         16401 => x"00001f64",
         16402 => x"00001f64",
         16403 => x"00001f64",
         16404 => x"00001f64",
         16405 => x"00001f64",
         16406 => x"00001f64",
         16407 => x"00001f64",
         16408 => x"00001f64",
         16409 => x"00001f64",
         16410 => x"00001f64",
         16411 => x"00001f64",
         16412 => x"00001f64",
         16413 => x"00001f64",
         16414 => x"00001f64",
         16415 => x"00001f64",
         16416 => x"00001f64",
         16417 => x"00001f64",
         16418 => x"00001f64",
         16419 => x"00001f64",
         16420 => x"00002481",
         16421 => x"00001f64",
         16422 => x"00001f64",
         16423 => x"00001f64",
         16424 => x"00001f64",
         16425 => x"00001f64",
         16426 => x"00001f64",
         16427 => x"00001f64",
         16428 => x"00001f64",
         16429 => x"00001f64",
         16430 => x"00001f64",
         16431 => x"00001f64",
         16432 => x"00001f64",
         16433 => x"00001f64",
         16434 => x"00001f64",
         16435 => x"00001f64",
         16436 => x"00001f64",
         16437 => x"00002417",
         16438 => x"00002316",
         16439 => x"00001f64",
         16440 => x"0000229a",
         16441 => x"000024b8",
         16442 => x"00002377",
         16443 => x"0000223c",
         16444 => x"000021de",
         16445 => x"00001f64",
         16446 => x"00001f64",
         16447 => x"00001f64",
         16448 => x"00001f64",
         16449 => x"00001f64",
         16450 => x"00001f64",
         16451 => x"00001f64",
         16452 => x"00001f64",
         16453 => x"00001f64",
         16454 => x"00001f64",
         16455 => x"00001f64",
         16456 => x"00001f64",
         16457 => x"00001f64",
         16458 => x"00001f64",
         16459 => x"00001f64",
         16460 => x"00001f64",
         16461 => x"00001f64",
         16462 => x"00001f64",
         16463 => x"00001f64",
         16464 => x"00001f64",
         16465 => x"00001f64",
         16466 => x"00001f64",
         16467 => x"00001f64",
         16468 => x"00001f64",
         16469 => x"00001f64",
         16470 => x"00001f64",
         16471 => x"00001f64",
         16472 => x"00001f64",
         16473 => x"00001f64",
         16474 => x"00001f64",
         16475 => x"00001f64",
         16476 => x"00001f64",
         16477 => x"00001f64",
         16478 => x"00001f64",
         16479 => x"00001f64",
         16480 => x"00001f64",
         16481 => x"00001f64",
         16482 => x"00001f64",
         16483 => x"00001f64",
         16484 => x"00001f64",
         16485 => x"00001f64",
         16486 => x"00001f64",
         16487 => x"00001f64",
         16488 => x"00001f64",
         16489 => x"00001f64",
         16490 => x"00001f64",
         16491 => x"00001f64",
         16492 => x"00001f64",
         16493 => x"00001f64",
         16494 => x"00001f64",
         16495 => x"00001f64",
         16496 => x"00001f64",
         16497 => x"000021bb",
         16498 => x"00002180",
         16499 => x"00001f64",
         16500 => x"00001f64",
         16501 => x"00001f64",
         16502 => x"00001f64",
         16503 => x"00001f64",
         16504 => x"00001f64",
         16505 => x"00001f64",
         16506 => x"00001f64",
         16507 => x"00002173",
         16508 => x"00002168",
         16509 => x"00001f64",
         16510 => x"00002150",
         16511 => x"00001f64",
         16512 => x"00002161",
         16513 => x"00002156",
         16514 => x"00002149",
         16515 => x"00003233",
         16516 => x"0000324b",
         16517 => x"00003257",
         16518 => x"00003263",
         16519 => x"0000326f",
         16520 => x"0000323f",
         16521 => x"00003c10",
         16522 => x"00003a9a",
         16523 => x"00003962",
         16524 => x"00003690",
         16525 => x"00003bac",
         16526 => x"000034fd",
         16527 => x"000037fc",
         16528 => x"000036b5",
         16529 => x"00003a44",
         16530 => x"000036e4",
         16531 => x"00003759",
         16532 => x"0000398b",
         16533 => x"000034fd",
         16534 => x"00003962",
         16535 => x"0000386c",
         16536 => x"000037fc",
         16537 => x"000034fd",
         16538 => x"000034fd",
         16539 => x"00003759",
         16540 => x"000036e4",
         16541 => x"000036b5",
         16542 => x"00003690",
         16543 => x"00004744",
         16544 => x"0000475d",
         16545 => x"00004782",
         16546 => x"000047a3",
         16547 => x"00004704",
         16548 => x"000047c8",
         16549 => x"0000471d",
         16550 => x"0000486d",
         16551 => x"0000482a",
         16552 => x"0000482a",
         16553 => x"0000482a",
         16554 => x"0000482a",
         16555 => x"0000482a",
         16556 => x"0000482a",
         16557 => x"00004803",
         16558 => x"0000482a",
         16559 => x"0000482a",
         16560 => x"0000482a",
         16561 => x"0000482a",
         16562 => x"0000482a",
         16563 => x"0000482a",
         16564 => x"0000482a",
         16565 => x"0000482a",
         16566 => x"0000482a",
         16567 => x"0000482a",
         16568 => x"0000482a",
         16569 => x"0000482a",
         16570 => x"0000482a",
         16571 => x"0000482a",
         16572 => x"0000482a",
         16573 => x"0000482a",
         16574 => x"0000482a",
         16575 => x"0000482a",
         16576 => x"0000482a",
         16577 => x"0000482a",
         16578 => x"0000482a",
         16579 => x"0000482a",
         16580 => x"00004942",
         16581 => x"00004930",
         16582 => x"0000491d",
         16583 => x"0000490a",
         16584 => x"00004834",
         16585 => x"000048f8",
         16586 => x"000048e5",
         16587 => x"0000484d",
         16588 => x"0000482a",
         16589 => x"0000484d",
         16590 => x"000048d5",
         16591 => x"00004952",
         16592 => x"0000487e",
         16593 => x"0000485c",
         16594 => x"000048c3",
         16595 => x"000048b1",
         16596 => x"0000489f",
         16597 => x"00004890",
         16598 => x"0000482a",
         16599 => x"00004834",
         16600 => x"000054d0",
         16601 => x"0000563f",
         16602 => x"00005611",
         16603 => x"00005568",
         16604 => x"00005545",
         16605 => x"00005524",
         16606 => x"000054fa",
         16607 => x"000056ca",
         16608 => x"00005351",
         16609 => x"000056a4",
         16610 => x"00005893",
         16611 => x"00005351",
         16612 => x"00005351",
         16613 => x"00005351",
         16614 => x"00005351",
         16615 => x"00005351",
         16616 => x"00005351",
         16617 => x"0000566d",
         16618 => x"0000587b",
         16619 => x"00005732",
         16620 => x"00005351",
         16621 => x"00005351",
         16622 => x"00005351",
         16623 => x"00005351",
         16624 => x"00005351",
         16625 => x"00005351",
         16626 => x"00005351",
         16627 => x"00005351",
         16628 => x"00005351",
         16629 => x"00005351",
         16630 => x"00005351",
         16631 => x"00005351",
         16632 => x"00005351",
         16633 => x"00005351",
         16634 => x"00005351",
         16635 => x"00005351",
         16636 => x"00005351",
         16637 => x"00005351",
         16638 => x"00005351",
         16639 => x"000055ef",
         16640 => x"00005351",
         16641 => x"00005351",
         16642 => x"00005351",
         16643 => x"00005592",
         16644 => x"000054a1",
         16645 => x"00005443",
         16646 => x"00005351",
         16647 => x"00005351",
         16648 => x"00005351",
         16649 => x"00005351",
         16650 => x"00005428",
         16651 => x"00005351",
         16652 => x"0000540b",
         16653 => x"00005a74",
         16654 => x"000059e9",
         16655 => x"000059e9",
         16656 => x"000059e9",
         16657 => x"000059e9",
         16658 => x"000059e9",
         16659 => x"000059e9",
         16660 => x"000059c4",
         16661 => x"000059e9",
         16662 => x"000059e9",
         16663 => x"000059e9",
         16664 => x"000059e9",
         16665 => x"000059e9",
         16666 => x"000059e9",
         16667 => x"000059e9",
         16668 => x"000059e9",
         16669 => x"000059e9",
         16670 => x"000059e9",
         16671 => x"000059e9",
         16672 => x"000059e9",
         16673 => x"000059e9",
         16674 => x"000059e9",
         16675 => x"000059e9",
         16676 => x"000059e9",
         16677 => x"000059e9",
         16678 => x"000059e9",
         16679 => x"000059e9",
         16680 => x"000059e9",
         16681 => x"000059e9",
         16682 => x"000059e9",
         16683 => x"00005a86",
         16684 => x"00005ace",
         16685 => x"00005abb",
         16686 => x"00005aa8",
         16687 => x"00005a96",
         16688 => x"00005b59",
         16689 => x"00005b46",
         16690 => x"00005b36",
         16691 => x"000059e9",
         16692 => x"00005b26",
         16693 => x"00005b16",
         16694 => x"00005b04",
         16695 => x"00005af2",
         16696 => x"00005ae0",
         16697 => x"00005a51",
         16698 => x"00005a40",
         16699 => x"00005a2f",
         16700 => x"00005a18",
         16701 => x"000059e9",
         16702 => x"00005a62",
         16703 => x"00006443",
         16704 => x"0000629f",
         16705 => x"0000629f",
         16706 => x"0000629f",
         16707 => x"0000629f",
         16708 => x"0000629f",
         16709 => x"0000629f",
         16710 => x"0000629f",
         16711 => x"0000629f",
         16712 => x"0000629f",
         16713 => x"0000629f",
         16714 => x"0000629f",
         16715 => x"0000629f",
         16716 => x"0000629f",
         16717 => x"00005fc1",
         16718 => x"0000629f",
         16719 => x"0000629f",
         16720 => x"0000629f",
         16721 => x"0000629f",
         16722 => x"0000629f",
         16723 => x"0000629f",
         16724 => x"0000648d",
         16725 => x"0000629f",
         16726 => x"0000629f",
         16727 => x"00006418",
         16728 => x"0000629f",
         16729 => x"0000642f",
         16730 => x"00005fa0",
         16731 => x"00006401",
         16732 => x"0000df74",
         16733 => x"0000df61",
         16734 => x"0000df55",
         16735 => x"0000df4a",
         16736 => x"0000df3f",
         16737 => x"0000df34",
         16738 => x"0000df29",
         16739 => x"0000df1d",
         16740 => x"0000df0f",
         16741 => x"00000e01",
         16742 => x"00000bfd",
         16743 => x"00000bfd",
         16744 => x"00000f49",
         16745 => x"00000bfd",
         16746 => x"00000bfd",
         16747 => x"00000bfd",
         16748 => x"00000bfd",
         16749 => x"00000bfd",
         16750 => x"00000bfd",
         16751 => x"00000bfd",
         16752 => x"00000dfd",
         16753 => x"00000bfd",
         16754 => x"00000f7f",
         16755 => x"00000f0d",
         16756 => x"00000bfd",
         16757 => x"00000bfd",
         16758 => x"00000bfd",
         16759 => x"00000bfd",
         16760 => x"00000bfd",
         16761 => x"00000bfd",
         16762 => x"00000bfd",
         16763 => x"00000bfd",
         16764 => x"00000bfd",
         16765 => x"00000bfd",
         16766 => x"00000bfd",
         16767 => x"00000bfd",
         16768 => x"00000bfd",
         16769 => x"00000bfd",
         16770 => x"00000bfd",
         16771 => x"00000bfd",
         16772 => x"00000bfd",
         16773 => x"00000bfd",
         16774 => x"00000bfd",
         16775 => x"00000bfd",
         16776 => x"00000bfd",
         16777 => x"00000bfd",
         16778 => x"00000bfd",
         16779 => x"00000bfd",
         16780 => x"00000bfd",
         16781 => x"00000bfd",
         16782 => x"00000bfd",
         16783 => x"00000bfd",
         16784 => x"00000bfd",
         16785 => x"00000bfd",
         16786 => x"00000bfd",
         16787 => x"00000bfd",
         16788 => x"00000bfd",
         16789 => x"00000bfd",
         16790 => x"00000bfd",
         16791 => x"00000bfd",
         16792 => x"00000f1d",
         16793 => x"00000bfd",
         16794 => x"00000bfd",
         16795 => x"00000bfd",
         16796 => x"00000bfd",
         16797 => x"00000e17",
         16798 => x"00000bfd",
         16799 => x"00000bfd",
         16800 => x"00000bfd",
         16801 => x"00000bfd",
         16802 => x"00000bfd",
         16803 => x"00000bfd",
         16804 => x"00000bfd",
         16805 => x"00000bfd",
         16806 => x"00000bfd",
         16807 => x"00000bfd",
         16808 => x"00000e2b",
         16809 => x"00000ee1",
         16810 => x"00000eb8",
         16811 => x"00000eb8",
         16812 => x"00000eb8",
         16813 => x"00000bfd",
         16814 => x"00000ee1",
         16815 => x"00000bfd",
         16816 => x"00000bfd",
         16817 => x"00000eff",
         16818 => x"00000bfd",
         16819 => x"00000bfd",
         16820 => x"00000c16",
         16821 => x"00000e0f",
         16822 => x"00000bfd",
         16823 => x"00000bfd",
         16824 => x"00000f58",
         16825 => x"00000bfd",
         16826 => x"00000c18",
         16827 => x"00000bfd",
         16828 => x"00000bfd",
         16829 => x"00000e17",
         16830 => x"64696e69",
         16831 => x"74000000",
         16832 => x"64696f63",
         16833 => x"746c0000",
         16834 => x"66696e69",
         16835 => x"74000000",
         16836 => x"666c6f61",
         16837 => x"64000000",
         16838 => x"66657865",
         16839 => x"63000000",
         16840 => x"6d636c65",
         16841 => x"61720000",
         16842 => x"6d636f70",
         16843 => x"79000000",
         16844 => x"6d646966",
         16845 => x"66000000",
         16846 => x"6d64756d",
         16847 => x"70000000",
         16848 => x"6d656200",
         16849 => x"6d656800",
         16850 => x"6d657700",
         16851 => x"68696400",
         16852 => x"68696500",
         16853 => x"68666400",
         16854 => x"68666500",
         16855 => x"63616c6c",
         16856 => x"00000000",
         16857 => x"6a6d7000",
         16858 => x"72657374",
         16859 => x"61727400",
         16860 => x"72657365",
         16861 => x"74000000",
         16862 => x"696e666f",
         16863 => x"00000000",
         16864 => x"74657374",
         16865 => x"00000000",
         16866 => x"636c7300",
         16867 => x"7a383000",
         16868 => x"74626173",
         16869 => x"69630000",
         16870 => x"6d626173",
         16871 => x"69630000",
         16872 => x"6b696c6f",
         16873 => x"00000000",
         16874 => x"65640000",
         16875 => x"556e6b6e",
         16876 => x"6f776e20",
         16877 => x"6572726f",
         16878 => x"722e0000",
         16879 => x"50617261",
         16880 => x"6d657465",
         16881 => x"72732069",
         16882 => x"6e636f72",
         16883 => x"72656374",
         16884 => x"2e000000",
         16885 => x"546f6f20",
         16886 => x"6d616e79",
         16887 => x"206f7065",
         16888 => x"6e206669",
         16889 => x"6c65732e",
         16890 => x"00000000",
         16891 => x"496e7375",
         16892 => x"66666963",
         16893 => x"69656e74",
         16894 => x"206d656d",
         16895 => x"6f72792e",
         16896 => x"00000000",
         16897 => x"46696c65",
         16898 => x"20697320",
         16899 => x"6c6f636b",
         16900 => x"65642e00",
         16901 => x"54696d65",
         16902 => x"6f75742c",
         16903 => x"206f7065",
         16904 => x"72617469",
         16905 => x"6f6e2063",
         16906 => x"616e6365",
         16907 => x"6c6c6564",
         16908 => x"2e000000",
         16909 => x"466f726d",
         16910 => x"61742061",
         16911 => x"626f7274",
         16912 => x"65642e00",
         16913 => x"4e6f2063",
         16914 => x"6f6d7061",
         16915 => x"7469626c",
         16916 => x"65206669",
         16917 => x"6c657379",
         16918 => x"7374656d",
         16919 => x"20666f75",
         16920 => x"6e64206f",
         16921 => x"6e206469",
         16922 => x"736b2e00",
         16923 => x"4469736b",
         16924 => x"206e6f74",
         16925 => x"20656e61",
         16926 => x"626c6564",
         16927 => x"2e000000",
         16928 => x"44726976",
         16929 => x"65206e75",
         16930 => x"6d626572",
         16931 => x"20697320",
         16932 => x"696e7661",
         16933 => x"6c69642e",
         16934 => x"00000000",
         16935 => x"53442069",
         16936 => x"73207772",
         16937 => x"69746520",
         16938 => x"70726f74",
         16939 => x"65637465",
         16940 => x"642e0000",
         16941 => x"46696c65",
         16942 => x"2068616e",
         16943 => x"646c6520",
         16944 => x"696e7661",
         16945 => x"6c69642e",
         16946 => x"00000000",
         16947 => x"46696c65",
         16948 => x"20616c72",
         16949 => x"65616479",
         16950 => x"20657869",
         16951 => x"7374732e",
         16952 => x"00000000",
         16953 => x"41636365",
         16954 => x"73732064",
         16955 => x"656e6965",
         16956 => x"642e0000",
         16957 => x"496e7661",
         16958 => x"6c696420",
         16959 => x"66696c65",
         16960 => x"6e616d65",
         16961 => x"2e000000",
         16962 => x"4e6f2070",
         16963 => x"61746820",
         16964 => x"666f756e",
         16965 => x"642e0000",
         16966 => x"4e6f2066",
         16967 => x"696c6520",
         16968 => x"666f756e",
         16969 => x"642e0000",
         16970 => x"4469736b",
         16971 => x"206e6f74",
         16972 => x"20726561",
         16973 => x"64792e00",
         16974 => x"496e7465",
         16975 => x"726e616c",
         16976 => x"20657272",
         16977 => x"6f722e00",
         16978 => x"4469736b",
         16979 => x"20457272",
         16980 => x"6f720000",
         16981 => x"53756363",
         16982 => x"6573732e",
         16983 => x"00000000",
         16984 => x"0a256c75",
         16985 => x"20627974",
         16986 => x"65732025",
         16987 => x"73206174",
         16988 => x"20256c75",
         16989 => x"20627974",
         16990 => x"65732f73",
         16991 => x"65632e0a",
         16992 => x"00000000",
         16993 => x"72656164",
         16994 => x"00000000",
         16995 => x"2530386c",
         16996 => x"58000000",
         16997 => x"3a202000",
         16998 => x"25303258",
         16999 => x"00000000",
         17000 => x"207c0000",
         17001 => x"7c000000",
         17002 => x"20200000",
         17003 => x"25303458",
         17004 => x"00000000",
         17005 => x"20202020",
         17006 => x"20202020",
         17007 => x"00000000",
         17008 => x"7a4f5300",
         17009 => x"2a2a2025",
         17010 => x"73202800",
         17011 => x"32352f30",
         17012 => x"372f3230",
         17013 => x"32310000",
         17014 => x"76312e33",
         17015 => x"32000000",
         17016 => x"205a5055",
         17017 => x"2c207265",
         17018 => x"76202530",
         17019 => x"32782920",
         17020 => x"25732025",
         17021 => x"73202a2a",
         17022 => x"0a0a0000",
         17023 => x"4f533a00",
         17024 => x"20202020",
         17025 => x"42617365",
         17026 => x"20416464",
         17027 => x"72657373",
         17028 => x"20202020",
         17029 => x"20202020",
         17030 => x"20202020",
         17031 => x"203d2025",
         17032 => x"30386c78",
         17033 => x"0a000000",
         17034 => x"20202020",
         17035 => x"41707020",
         17036 => x"41646472",
         17037 => x"65737320",
         17038 => x"20202020",
         17039 => x"20202020",
         17040 => x"20202020",
         17041 => x"203d2025",
         17042 => x"30386c78",
         17043 => x"0a000000",
         17044 => x"5a505520",
         17045 => x"496e7465",
         17046 => x"72727570",
         17047 => x"74204861",
         17048 => x"6e646c65",
         17049 => x"72000000",
         17050 => x"55415254",
         17051 => x"31205458",
         17052 => x"20696e74",
         17053 => x"65727275",
         17054 => x"70740000",
         17055 => x"55415254",
         17056 => x"31205258",
         17057 => x"20696e74",
         17058 => x"65727275",
         17059 => x"70740000",
         17060 => x"55415254",
         17061 => x"30205458",
         17062 => x"20696e74",
         17063 => x"65727275",
         17064 => x"70740000",
         17065 => x"55415254",
         17066 => x"30205258",
         17067 => x"20696e74",
         17068 => x"65727275",
         17069 => x"70740000",
         17070 => x"494f4354",
         17071 => x"4c205752",
         17072 => x"20696e74",
         17073 => x"65727275",
         17074 => x"70740000",
         17075 => x"494f4354",
         17076 => x"4c205244",
         17077 => x"20696e74",
         17078 => x"65727275",
         17079 => x"70740000",
         17080 => x"50533220",
         17081 => x"696e7465",
         17082 => x"72727570",
         17083 => x"74000000",
         17084 => x"54696d65",
         17085 => x"7220696e",
         17086 => x"74657272",
         17087 => x"75707400",
         17088 => x"53657474",
         17089 => x"696e6720",
         17090 => x"75702074",
         17091 => x"696d6572",
         17092 => x"2e2e2e00",
         17093 => x"456e6162",
         17094 => x"6c696e67",
         17095 => x"2074696d",
         17096 => x"65722e2e",
         17097 => x"2e000000",
         17098 => x"6175746f",
         17099 => x"65786563",
         17100 => x"2e626174",
         17101 => x"00000000",
         17102 => x"7a4f535f",
         17103 => x"7a70752e",
         17104 => x"68737400",
         17105 => x"4661696c",
         17106 => x"65642074",
         17107 => x"6f20696e",
         17108 => x"69746961",
         17109 => x"6c697365",
         17110 => x"20736420",
         17111 => x"63617264",
         17112 => x"20302c20",
         17113 => x"706c6561",
         17114 => x"73652069",
         17115 => x"6e697420",
         17116 => x"6d616e75",
         17117 => x"616c6c79",
         17118 => x"2e000000",
         17119 => x"2a200000",
         17120 => x"25643a5c",
         17121 => x"25730000",
         17122 => x"303a0000",
         17123 => x"42616420",
         17124 => x"636f6d6d",
         17125 => x"616e642e",
         17126 => x"00000000",
         17127 => x"5a505500",
         17128 => x"62696e00",
         17129 => x"25643a5c",
         17130 => x"25735c25",
         17131 => x"732e2573",
         17132 => x"00000000",
         17133 => x"436f6c64",
         17134 => x"20726562",
         17135 => x"6f6f7469",
         17136 => x"6e672e2e",
         17137 => x"2e000000",
         17138 => x"52657374",
         17139 => x"61727469",
         17140 => x"6e672061",
         17141 => x"70706c69",
         17142 => x"63617469",
         17143 => x"6f6e2e2e",
         17144 => x"2e000000",
         17145 => x"43616c6c",
         17146 => x"696e6720",
         17147 => x"636f6465",
         17148 => x"20402025",
         17149 => x"30386c78",
         17150 => x"202e2e2e",
         17151 => x"0a000000",
         17152 => x"43616c6c",
         17153 => x"20726574",
         17154 => x"75726e65",
         17155 => x"6420636f",
         17156 => x"64652028",
         17157 => x"2564292e",
         17158 => x"0a000000",
         17159 => x"45786563",
         17160 => x"7574696e",
         17161 => x"6720636f",
         17162 => x"64652040",
         17163 => x"20253038",
         17164 => x"6c78202e",
         17165 => x"2e2e0a00",
         17166 => x"2530386c",
         17167 => x"58202530",
         17168 => x"386c582d",
         17169 => x"00000000",
         17170 => x"2530386c",
         17171 => x"58202530",
         17172 => x"34582d00",
         17173 => x"436f6d70",
         17174 => x"6172696e",
         17175 => x"672e2e2e",
         17176 => x"00000000",
         17177 => x"2530386c",
         17178 => x"78282530",
         17179 => x"3878292d",
         17180 => x"3e253038",
         17181 => x"6c782825",
         17182 => x"30387829",
         17183 => x"0a000000",
         17184 => x"436f7079",
         17185 => x"696e672e",
         17186 => x"2e2e0000",
         17187 => x"2530386c",
         17188 => x"58202530",
         17189 => x"32582d00",
         17190 => x"436c6561",
         17191 => x"72696e67",
         17192 => x"2e2e2e2e",
         17193 => x"00000000",
         17194 => x"44756d70",
         17195 => x"204d656d",
         17196 => x"6f727900",
         17197 => x"0a436f6d",
         17198 => x"706c6574",
         17199 => x"652e0000",
         17200 => x"25643a5c",
         17201 => x"25735c25",
         17202 => x"73000000",
         17203 => x"4d656d6f",
         17204 => x"72792065",
         17205 => x"78686175",
         17206 => x"73746564",
         17207 => x"2c206361",
         17208 => x"6e6e6f74",
         17209 => x"2070726f",
         17210 => x"63657373",
         17211 => x"20636f6d",
         17212 => x"6d616e64",
         17213 => x"2e000000",
         17214 => x"3f3f3f00",
         17215 => x"25642f25",
         17216 => x"642f2564",
         17217 => x"2025643a",
         17218 => x"25643a25",
         17219 => x"642e2564",
         17220 => x"25640a00",
         17221 => x"536f4320",
         17222 => x"436f6e66",
         17223 => x"69677572",
         17224 => x"6174696f",
         17225 => x"6e000000",
         17226 => x"3a0a4465",
         17227 => x"76696365",
         17228 => x"7320696d",
         17229 => x"706c656d",
         17230 => x"656e7465",
         17231 => x"643a0000",
         17232 => x"41646472",
         17233 => x"65737365",
         17234 => x"733a0000",
         17235 => x"20202020",
         17236 => x"43505520",
         17237 => x"52657365",
         17238 => x"74205665",
         17239 => x"63746f72",
         17240 => x"20416464",
         17241 => x"72657373",
         17242 => x"203d2025",
         17243 => x"3038580a",
         17244 => x"00000000",
         17245 => x"20202020",
         17246 => x"43505520",
         17247 => x"4d656d6f",
         17248 => x"72792053",
         17249 => x"74617274",
         17250 => x"20416464",
         17251 => x"72657373",
         17252 => x"203d2025",
         17253 => x"3038580a",
         17254 => x"00000000",
         17255 => x"20202020",
         17256 => x"53746163",
         17257 => x"6b205374",
         17258 => x"61727420",
         17259 => x"41646472",
         17260 => x"65737320",
         17261 => x"20202020",
         17262 => x"203d2025",
         17263 => x"3038580a",
         17264 => x"00000000",
         17265 => x"4d697363",
         17266 => x"3a000000",
         17267 => x"20202020",
         17268 => x"5a505520",
         17269 => x"49642020",
         17270 => x"20202020",
         17271 => x"20202020",
         17272 => x"20202020",
         17273 => x"20202020",
         17274 => x"203d2025",
         17275 => x"3034580a",
         17276 => x"00000000",
         17277 => x"20202020",
         17278 => x"53797374",
         17279 => x"656d2043",
         17280 => x"6c6f636b",
         17281 => x"20467265",
         17282 => x"71202020",
         17283 => x"20202020",
         17284 => x"203d2025",
         17285 => x"642e2530",
         17286 => x"34644d48",
         17287 => x"7a0a0000",
         17288 => x"20202020",
         17289 => x"57697368",
         17290 => x"626f6e65",
         17291 => x"20534452",
         17292 => x"414d2043",
         17293 => x"6c6f636b",
         17294 => x"20467265",
         17295 => x"713d2025",
         17296 => x"642e2530",
         17297 => x"34644d48",
         17298 => x"7a0a0000",
         17299 => x"20202020",
         17300 => x"53445241",
         17301 => x"4d20436c",
         17302 => x"6f636b20",
         17303 => x"46726571",
         17304 => x"20202020",
         17305 => x"20202020",
         17306 => x"203d2025",
         17307 => x"642e2530",
         17308 => x"34644d48",
         17309 => x"7a0a0000",
         17310 => x"20202020",
         17311 => x"53504900",
         17312 => x"20202020",
         17313 => x"50533200",
         17314 => x"20202020",
         17315 => x"494f4354",
         17316 => x"4c000000",
         17317 => x"20202020",
         17318 => x"57422049",
         17319 => x"32430000",
         17320 => x"20202020",
         17321 => x"57495348",
         17322 => x"424f4e45",
         17323 => x"20425553",
         17324 => x"00000000",
         17325 => x"20202020",
         17326 => x"494e5452",
         17327 => x"20435452",
         17328 => x"4c202843",
         17329 => x"68616e6e",
         17330 => x"656c733d",
         17331 => x"25303264",
         17332 => x"292e0a00",
         17333 => x"20202020",
         17334 => x"54494d45",
         17335 => x"52312020",
         17336 => x"20202854",
         17337 => x"696d6572",
         17338 => x"7320203d",
         17339 => x"25303264",
         17340 => x"292e0a00",
         17341 => x"20202020",
         17342 => x"53442043",
         17343 => x"41524420",
         17344 => x"20202844",
         17345 => x"65766963",
         17346 => x"6573203d",
         17347 => x"25303264",
         17348 => x"292e0a00",
         17349 => x"20202020",
         17350 => x"52414d20",
         17351 => x"20202020",
         17352 => x"20202825",
         17353 => x"3038583a",
         17354 => x"25303858",
         17355 => x"292e0a00",
         17356 => x"20202020",
         17357 => x"4252414d",
         17358 => x"20202020",
         17359 => x"20202825",
         17360 => x"3038583a",
         17361 => x"25303858",
         17362 => x"292e0a00",
         17363 => x"20202020",
         17364 => x"494e534e",
         17365 => x"20425241",
         17366 => x"4d202825",
         17367 => x"3038583a",
         17368 => x"25303858",
         17369 => x"292e0a00",
         17370 => x"20202020",
         17371 => x"53445241",
         17372 => x"4d202020",
         17373 => x"20202825",
         17374 => x"3038583a",
         17375 => x"25303858",
         17376 => x"292e0a00",
         17377 => x"20202020",
         17378 => x"57422053",
         17379 => x"4452414d",
         17380 => x"20202825",
         17381 => x"3038583a",
         17382 => x"25303858",
         17383 => x"292e0a00",
         17384 => x"20286672",
         17385 => x"6f6d2053",
         17386 => x"6f432063",
         17387 => x"6f6e6669",
         17388 => x"67290000",
         17389 => x"556e6b6e",
         17390 => x"6f776e00",
         17391 => x"45564f6d",
         17392 => x"00000000",
         17393 => x"536d616c",
         17394 => x"6c000000",
         17395 => x"4d656469",
         17396 => x"756d0000",
         17397 => x"466c6578",
         17398 => x"00000000",
         17399 => x"45564f00",
         17400 => x"0000f13c",
         17401 => x"01000000",
         17402 => x"00000002",
         17403 => x"0000f138",
         17404 => x"01000000",
         17405 => x"00000003",
         17406 => x"0000f134",
         17407 => x"01000000",
         17408 => x"00000004",
         17409 => x"0000f130",
         17410 => x"01000000",
         17411 => x"00000005",
         17412 => x"0000f12c",
         17413 => x"01000000",
         17414 => x"00000006",
         17415 => x"0000f128",
         17416 => x"01000000",
         17417 => x"00000007",
         17418 => x"0000f124",
         17419 => x"01000000",
         17420 => x"00000001",
         17421 => x"0000f120",
         17422 => x"01000000",
         17423 => x"00000008",
         17424 => x"0000f11c",
         17425 => x"01000000",
         17426 => x"0000000b",
         17427 => x"0000f118",
         17428 => x"01000000",
         17429 => x"00000009",
         17430 => x"0000f114",
         17431 => x"01000000",
         17432 => x"0000000a",
         17433 => x"0000f110",
         17434 => x"04000000",
         17435 => x"0000000d",
         17436 => x"0000f10c",
         17437 => x"04000000",
         17438 => x"0000000c",
         17439 => x"0000f108",
         17440 => x"04000000",
         17441 => x"0000000e",
         17442 => x"0000f104",
         17443 => x"03000000",
         17444 => x"0000000f",
         17445 => x"0000f100",
         17446 => x"04000000",
         17447 => x"0000000f",
         17448 => x"0000f0fc",
         17449 => x"04000000",
         17450 => x"00000010",
         17451 => x"0000f0f8",
         17452 => x"04000000",
         17453 => x"00000011",
         17454 => x"0000f0f4",
         17455 => x"03000000",
         17456 => x"00000012",
         17457 => x"0000f0f0",
         17458 => x"03000000",
         17459 => x"00000013",
         17460 => x"0000f0ec",
         17461 => x"03000000",
         17462 => x"00000014",
         17463 => x"0000f0e8",
         17464 => x"03000000",
         17465 => x"00000015",
         17466 => x"1b5b4400",
         17467 => x"1b5b4300",
         17468 => x"1b5b4200",
         17469 => x"1b5b4100",
         17470 => x"1b5b367e",
         17471 => x"1b5b357e",
         17472 => x"1b5b347e",
         17473 => x"1b304600",
         17474 => x"1b5b337e",
         17475 => x"1b5b327e",
         17476 => x"1b5b317e",
         17477 => x"10000000",
         17478 => x"0e000000",
         17479 => x"0d000000",
         17480 => x"0b000000",
         17481 => x"08000000",
         17482 => x"06000000",
         17483 => x"05000000",
         17484 => x"04000000",
         17485 => x"03000000",
         17486 => x"02000000",
         17487 => x"01000000",
         17488 => x"48697374",
         17489 => x"6f727920",
         17490 => x"68656170",
         17491 => x"3a253038",
         17492 => x"6c780a00",
         17493 => x"43616e6e",
         17494 => x"6f74206f",
         17495 => x"70656e2f",
         17496 => x"63726561",
         17497 => x"74652068",
         17498 => x"6973746f",
         17499 => x"72792066",
         17500 => x"696c652c",
         17501 => x"20646973",
         17502 => x"61626c69",
         17503 => x"6e672e00",
         17504 => x"68697374",
         17505 => x"6f727900",
         17506 => x"68697374",
         17507 => x"00000000",
         17508 => x"21000000",
         17509 => x"48697374",
         17510 => x"6f727920",
         17511 => x"62756666",
         17512 => x"65724025",
         17513 => x"30386c78",
         17514 => x"0a000000",
         17515 => x"2530366c",
         17516 => x"75202025",
         17517 => x"730a0000",
         17518 => x"4661696c",
         17519 => x"65642074",
         17520 => x"6f207265",
         17521 => x"73657420",
         17522 => x"74686520",
         17523 => x"68697374",
         17524 => x"6f727920",
         17525 => x"66696c65",
         17526 => x"20746f20",
         17527 => x"454f462e",
         17528 => x"00000000",
         17529 => x"3e25730a",
         17530 => x"00000000",
         17531 => x"1b5b317e",
         17532 => x"00000000",
         17533 => x"1b5b4100",
         17534 => x"1b5b4200",
         17535 => x"1b5b4300",
         17536 => x"1b5b4400",
         17537 => x"1b5b3130",
         17538 => x"7e000000",
         17539 => x"1b5b3131",
         17540 => x"7e000000",
         17541 => x"1b5b3132",
         17542 => x"7e000000",
         17543 => x"1b5b3133",
         17544 => x"7e000000",
         17545 => x"1b5b3134",
         17546 => x"7e000000",
         17547 => x"1b5b3135",
         17548 => x"7e000000",
         17549 => x"1b5b3137",
         17550 => x"7e000000",
         17551 => x"1b5b3138",
         17552 => x"7e000000",
         17553 => x"1b5b3139",
         17554 => x"7e000000",
         17555 => x"1b5b3230",
         17556 => x"7e000000",
         17557 => x"1b5b327e",
         17558 => x"00000000",
         17559 => x"1b5b337e",
         17560 => x"00000000",
         17561 => x"1b5b4600",
         17562 => x"1b5b357e",
         17563 => x"00000000",
         17564 => x"1b5b367e",
         17565 => x"00000000",
         17566 => x"583a2564",
         17567 => x"2c25642c",
         17568 => x"25642c25",
         17569 => x"642c2564",
         17570 => x"2c25643a",
         17571 => x"25303278",
         17572 => x"00000000",
         17573 => x"443a2564",
         17574 => x"2d25642d",
         17575 => x"25643a25",
         17576 => x"633a2564",
         17577 => x"2c25642c",
         17578 => x"25643a00",
         17579 => x"25642c00",
         17580 => x"4b3a2564",
         17581 => x"3a000000",
         17582 => x"25303278",
         17583 => x"2c000000",
         17584 => x"25635b25",
         17585 => x"643b2564",
         17586 => x"52000000",
         17587 => x"5265706f",
         17588 => x"72742043",
         17589 => x"7572736f",
         17590 => x"723a0000",
         17591 => x"55703a25",
         17592 => x"30327820",
         17593 => x"25303278",
         17594 => x"00000000",
         17595 => x"44773a25",
         17596 => x"30327820",
         17597 => x"25303278",
         17598 => x"00000000",
         17599 => x"48643a25",
         17600 => x"30327820",
         17601 => x"00000000",
         17602 => x"4e6f2074",
         17603 => x"65737420",
         17604 => x"64656669",
         17605 => x"6e65642e",
         17606 => x"00000000",
         17607 => x"53440000",
         17608 => x"222a3a3c",
         17609 => x"3e3f7c7f",
         17610 => x"00000000",
         17611 => x"2b2c3b3d",
         17612 => x"5b5d0000",
         17613 => x"46415400",
         17614 => x"46415433",
         17615 => x"32000000",
         17616 => x"ebfe904d",
         17617 => x"53444f53",
         17618 => x"352e3000",
         17619 => x"4e4f204e",
         17620 => x"414d4520",
         17621 => x"20202046",
         17622 => x"41542020",
         17623 => x"20202000",
         17624 => x"4e4f204e",
         17625 => x"414d4520",
         17626 => x"20202046",
         17627 => x"41543332",
         17628 => x"20202000",
         17629 => x"0000f31c",
         17630 => x"00000000",
         17631 => x"00000000",
         17632 => x"00000000",
         17633 => x"01030507",
         17634 => x"090e1012",
         17635 => x"1416181c",
         17636 => x"1e000000",
         17637 => x"809a4541",
         17638 => x"8e418f80",
         17639 => x"45454549",
         17640 => x"49498e8f",
         17641 => x"9092924f",
         17642 => x"994f5555",
         17643 => x"59999a9b",
         17644 => x"9c9d9e9f",
         17645 => x"41494f55",
         17646 => x"a5a5a6a7",
         17647 => x"a8a9aaab",
         17648 => x"acadaeaf",
         17649 => x"b0b1b2b3",
         17650 => x"b4b5b6b7",
         17651 => x"b8b9babb",
         17652 => x"bcbdbebf",
         17653 => x"c0c1c2c3",
         17654 => x"c4c5c6c7",
         17655 => x"c8c9cacb",
         17656 => x"cccdcecf",
         17657 => x"d0d1d2d3",
         17658 => x"d4d5d6d7",
         17659 => x"d8d9dadb",
         17660 => x"dcdddedf",
         17661 => x"e0e1e2e3",
         17662 => x"e4e5e6e7",
         17663 => x"e8e9eaeb",
         17664 => x"ecedeeef",
         17665 => x"f0f1f2f3",
         17666 => x"f4f5f6f7",
         17667 => x"f8f9fafb",
         17668 => x"fcfdfeff",
         17669 => x"2b2e2c3b",
         17670 => x"3d5b5d2f",
         17671 => x"5c222a3a",
         17672 => x"3c3e3f7c",
         17673 => x"7f000000",
         17674 => x"00010004",
         17675 => x"00100040",
         17676 => x"01000200",
         17677 => x"00000000",
         17678 => x"00010002",
         17679 => x"00040008",
         17680 => x"00100020",
         17681 => x"00000000",
         17682 => x"00c700fc",
         17683 => x"00e900e2",
         17684 => x"00e400e0",
         17685 => x"00e500e7",
         17686 => x"00ea00eb",
         17687 => x"00e800ef",
         17688 => x"00ee00ec",
         17689 => x"00c400c5",
         17690 => x"00c900e6",
         17691 => x"00c600f4",
         17692 => x"00f600f2",
         17693 => x"00fb00f9",
         17694 => x"00ff00d6",
         17695 => x"00dc00a2",
         17696 => x"00a300a5",
         17697 => x"20a70192",
         17698 => x"00e100ed",
         17699 => x"00f300fa",
         17700 => x"00f100d1",
         17701 => x"00aa00ba",
         17702 => x"00bf2310",
         17703 => x"00ac00bd",
         17704 => x"00bc00a1",
         17705 => x"00ab00bb",
         17706 => x"25912592",
         17707 => x"25932502",
         17708 => x"25242561",
         17709 => x"25622556",
         17710 => x"25552563",
         17711 => x"25512557",
         17712 => x"255d255c",
         17713 => x"255b2510",
         17714 => x"25142534",
         17715 => x"252c251c",
         17716 => x"2500253c",
         17717 => x"255e255f",
         17718 => x"255a2554",
         17719 => x"25692566",
         17720 => x"25602550",
         17721 => x"256c2567",
         17722 => x"25682564",
         17723 => x"25652559",
         17724 => x"25582552",
         17725 => x"2553256b",
         17726 => x"256a2518",
         17727 => x"250c2588",
         17728 => x"2584258c",
         17729 => x"25902580",
         17730 => x"03b100df",
         17731 => x"039303c0",
         17732 => x"03a303c3",
         17733 => x"00b503c4",
         17734 => x"03a60398",
         17735 => x"03a903b4",
         17736 => x"221e03c6",
         17737 => x"03b52229",
         17738 => x"226100b1",
         17739 => x"22652264",
         17740 => x"23202321",
         17741 => x"00f72248",
         17742 => x"00b02219",
         17743 => x"00b7221a",
         17744 => x"207f00b2",
         17745 => x"25a000a0",
         17746 => x"0061031a",
         17747 => x"00e00317",
         17748 => x"00f80307",
         17749 => x"00ff0001",
         17750 => x"01780100",
         17751 => x"01300132",
         17752 => x"01060139",
         17753 => x"0110014a",
         17754 => x"012e0179",
         17755 => x"01060180",
         17756 => x"004d0243",
         17757 => x"01810182",
         17758 => x"01820184",
         17759 => x"01840186",
         17760 => x"01870187",
         17761 => x"0189018a",
         17762 => x"018b018b",
         17763 => x"018d018e",
         17764 => x"018f0190",
         17765 => x"01910191",
         17766 => x"01930194",
         17767 => x"01f60196",
         17768 => x"01970198",
         17769 => x"0198023d",
         17770 => x"019b019c",
         17771 => x"019d0220",
         17772 => x"019f01a0",
         17773 => x"01a001a2",
         17774 => x"01a201a4",
         17775 => x"01a401a6",
         17776 => x"01a701a7",
         17777 => x"01a901aa",
         17778 => x"01ab01ac",
         17779 => x"01ac01ae",
         17780 => x"01af01af",
         17781 => x"01b101b2",
         17782 => x"01b301b3",
         17783 => x"01b501b5",
         17784 => x"01b701b8",
         17785 => x"01b801ba",
         17786 => x"01bb01bc",
         17787 => x"01bc01be",
         17788 => x"01f701c0",
         17789 => x"01c101c2",
         17790 => x"01c301c4",
         17791 => x"01c501c4",
         17792 => x"01c701c8",
         17793 => x"01c701ca",
         17794 => x"01cb01ca",
         17795 => x"01cd0110",
         17796 => x"01dd0001",
         17797 => x"018e01de",
         17798 => x"011201f3",
         17799 => x"000301f1",
         17800 => x"01f401f4",
         17801 => x"01f80128",
         17802 => x"02220112",
         17803 => x"023a0009",
         17804 => x"2c65023b",
         17805 => x"023b023d",
         17806 => x"2c66023f",
         17807 => x"02400241",
         17808 => x"02410246",
         17809 => x"010a0253",
         17810 => x"00400181",
         17811 => x"01860255",
         17812 => x"0189018a",
         17813 => x"0258018f",
         17814 => x"025a0190",
         17815 => x"025c025d",
         17816 => x"025e025f",
         17817 => x"01930261",
         17818 => x"02620194",
         17819 => x"02640265",
         17820 => x"02660267",
         17821 => x"01970196",
         17822 => x"026a2c62",
         17823 => x"026c026d",
         17824 => x"026e019c",
         17825 => x"02700271",
         17826 => x"019d0273",
         17827 => x"0274019f",
         17828 => x"02760277",
         17829 => x"02780279",
         17830 => x"027a027b",
         17831 => x"027c2c64",
         17832 => x"027e027f",
         17833 => x"01a60281",
         17834 => x"028201a9",
         17835 => x"02840285",
         17836 => x"02860287",
         17837 => x"01ae0244",
         17838 => x"01b101b2",
         17839 => x"0245028d",
         17840 => x"028e028f",
         17841 => x"02900291",
         17842 => x"01b7037b",
         17843 => x"000303fd",
         17844 => x"03fe03ff",
         17845 => x"03ac0004",
         17846 => x"03860388",
         17847 => x"0389038a",
         17848 => x"03b10311",
         17849 => x"03c20002",
         17850 => x"03a303a3",
         17851 => x"03c40308",
         17852 => x"03cc0003",
         17853 => x"038c038e",
         17854 => x"038f03d8",
         17855 => x"011803f2",
         17856 => x"000a03f9",
         17857 => x"03f303f4",
         17858 => x"03f503f6",
         17859 => x"03f703f7",
         17860 => x"03f903fa",
         17861 => x"03fa0430",
         17862 => x"03200450",
         17863 => x"07100460",
         17864 => x"0122048a",
         17865 => x"013604c1",
         17866 => x"010e04cf",
         17867 => x"000104c0",
         17868 => x"04d00144",
         17869 => x"05610426",
         17870 => x"00000000",
         17871 => x"1d7d0001",
         17872 => x"2c631e00",
         17873 => x"01961ea0",
         17874 => x"015a1f00",
         17875 => x"06081f10",
         17876 => x"06061f20",
         17877 => x"06081f30",
         17878 => x"06081f40",
         17879 => x"06061f51",
         17880 => x"00071f59",
         17881 => x"1f521f5b",
         17882 => x"1f541f5d",
         17883 => x"1f561f5f",
         17884 => x"1f600608",
         17885 => x"1f70000e",
         17886 => x"1fba1fbb",
         17887 => x"1fc81fc9",
         17888 => x"1fca1fcb",
         17889 => x"1fda1fdb",
         17890 => x"1ff81ff9",
         17891 => x"1fea1feb",
         17892 => x"1ffa1ffb",
         17893 => x"1f800608",
         17894 => x"1f900608",
         17895 => x"1fa00608",
         17896 => x"1fb00004",
         17897 => x"1fb81fb9",
         17898 => x"1fb21fbc",
         17899 => x"1fcc0001",
         17900 => x"1fc31fd0",
         17901 => x"06021fe0",
         17902 => x"06021fe5",
         17903 => x"00011fec",
         17904 => x"1ff30001",
         17905 => x"1ffc214e",
         17906 => x"00012132",
         17907 => x"21700210",
         17908 => x"21840001",
         17909 => x"218324d0",
         17910 => x"051a2c30",
         17911 => x"042f2c60",
         17912 => x"01022c67",
         17913 => x"01062c75",
         17914 => x"01022c80",
         17915 => x"01642d00",
         17916 => x"0826ff41",
         17917 => x"031a0000",
         17918 => x"00000000",
         17919 => x"0000e6f8",
         17920 => x"01020100",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"0000e700",
         17924 => x"01040100",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"0000e708",
         17928 => x"01140300",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"0000e710",
         17932 => x"012b0300",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"0000e718",
         17936 => x"01300300",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"0000e720",
         17940 => x"013c0400",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"0000e728",
         17944 => x"013d0400",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"0000e730",
         17948 => x"013f0400",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"0000e738",
         17952 => x"01400400",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"0000e740",
         17956 => x"01410400",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"0000e744",
         17960 => x"01420400",
         17961 => x"00000000",
         17962 => x"00000000",
         17963 => x"0000e748",
         17964 => x"01430400",
         17965 => x"00000000",
         17966 => x"00000000",
         17967 => x"0000e74c",
         17968 => x"01500500",
         17969 => x"00000000",
         17970 => x"00000000",
         17971 => x"0000e750",
         17972 => x"01510500",
         17973 => x"00000000",
         17974 => x"00000000",
         17975 => x"0000e754",
         17976 => x"01540500",
         17977 => x"00000000",
         17978 => x"00000000",
         17979 => x"0000e758",
         17980 => x"01550500",
         17981 => x"00000000",
         17982 => x"00000000",
         17983 => x"0000e75c",
         17984 => x"01790700",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"0000e764",
         17988 => x"01780700",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"0000e768",
         17992 => x"01820800",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"0000e770",
         17996 => x"01830800",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"0000e778",
         18000 => x"01850800",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"0000e780",
         18004 => x"01870800",
         18005 => x"00000000",
         18006 => x"00000000",
         18007 => x"0000e788",
         18008 => x"01880800",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"0000e78c",
         18012 => x"01890800",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"0000e790",
         18016 => x"018c0900",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"0000e798",
         18020 => x"018d0900",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"0000e7a0",
         18024 => x"018e0900",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"0000e7a8",
         18028 => x"018f0900",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00007fff",
         18034 => x"00000000",
         18035 => x"00007fff",
         18036 => x"00010000",
         18037 => x"00007fff",
         18038 => x"00010000",
         18039 => x"00810000",
         18040 => x"01000000",
         18041 => x"017fffff",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00007800",
         18045 => x"00000000",
         18046 => x"05f5e100",
         18047 => x"05f5e100",
         18048 => x"05f5e100",
         18049 => x"00000000",
         18050 => x"01010101",
         18051 => x"01010101",
         18052 => x"01011001",
         18053 => x"01000000",
         18054 => x"00000000",
         18055 => x"00000000",
         18056 => x"00000000",
         18057 => x"00000000",
         18058 => x"00000000",
         18059 => x"00000000",
         18060 => x"00000000",
         18061 => x"00000000",
         18062 => x"00000000",
         18063 => x"00000000",
         18064 => x"00000000",
         18065 => x"00000000",
         18066 => x"00000000",
         18067 => x"00000000",
         18068 => x"00000000",
         18069 => x"00000000",
         18070 => x"00000000",
         18071 => x"00000000",
         18072 => x"00000000",
         18073 => x"00000000",
         18074 => x"00000000",
         18075 => x"00000000",
         18076 => x"00000000",
         18077 => x"00000000",
         18078 => x"0000f180",
         18079 => x"01000000",
         18080 => x"0000f188",
         18081 => x"01000000",
         18082 => x"0000f190",
         18083 => x"02000000",
         18084 => x"0001fd80",
         18085 => x"1bfc5ffd",
         18086 => x"f03b3a0d",
         18087 => x"797a405b",
         18088 => x"5df0f0f0",
         18089 => x"71727374",
         18090 => x"75767778",
         18091 => x"696a6b6c",
         18092 => x"6d6e6f70",
         18093 => x"61626364",
         18094 => x"65666768",
         18095 => x"31323334",
         18096 => x"35363738",
         18097 => x"5cf32d20",
         18098 => x"30392c2e",
         18099 => x"f67ff3f4",
         18100 => x"f1f23f2f",
         18101 => x"08f0f0f0",
         18102 => x"f0f0f0f0",
         18103 => x"80818283",
         18104 => x"84f0f0f0",
         18105 => x"1bfc58fd",
         18106 => x"f03a3b0d",
         18107 => x"595a405b",
         18108 => x"5df0f0f0",
         18109 => x"51525354",
         18110 => x"55565758",
         18111 => x"494a4b4c",
         18112 => x"4d4e4f50",
         18113 => x"41424344",
         18114 => x"45464748",
         18115 => x"31323334",
         18116 => x"35363738",
         18117 => x"5cf32d20",
         18118 => x"30392c2e",
         18119 => x"f67ff3f4",
         18120 => x"f1f23f2f",
         18121 => x"08f0f0f0",
         18122 => x"f0f0f0f0",
         18123 => x"80818283",
         18124 => x"84f0f0f0",
         18125 => x"1bfc58fd",
         18126 => x"f02b2a0d",
         18127 => x"595a607b",
         18128 => x"7df0f0f0",
         18129 => x"51525354",
         18130 => x"55565758",
         18131 => x"494a4b4c",
         18132 => x"4d4e4f50",
         18133 => x"41424344",
         18134 => x"45464748",
         18135 => x"21222324",
         18136 => x"25262728",
         18137 => x"7c7e3d20",
         18138 => x"20293c3e",
         18139 => x"f7e2e0e1",
         18140 => x"f9f83f2f",
         18141 => x"fbf0f0f0",
         18142 => x"f0f0f0f0",
         18143 => x"85868788",
         18144 => x"89f0f0f0",
         18145 => x"1bfe1efa",
         18146 => x"f0f0f0f0",
         18147 => x"191a001b",
         18148 => x"1df0f0f0",
         18149 => x"11121314",
         18150 => x"15161718",
         18151 => x"090a0b0c",
         18152 => x"0d0e0f10",
         18153 => x"01020304",
         18154 => x"05060708",
         18155 => x"f0f0f0f0",
         18156 => x"f0f0f0f0",
         18157 => x"f01ef0f0",
         18158 => x"f01ff0f0",
         18159 => x"f0f0f0f0",
         18160 => x"f0f0f01c",
         18161 => x"f0f0f0f0",
         18162 => x"f0f0f0f0",
         18163 => x"80818283",
         18164 => x"84f0f0f0",
         18165 => x"bff0cfc9",
         18166 => x"f0b54dcd",
         18167 => x"3577d7b3",
         18168 => x"b7f0f0f0",
         18169 => x"7c704131",
         18170 => x"39a678dd",
         18171 => x"3d5d6c56",
         18172 => x"1d33d5b1",
         18173 => x"466ed948",
         18174 => x"74434c73",
         18175 => x"3f367e3b",
         18176 => x"7a1e5fa2",
         18177 => x"d39fd100",
         18178 => x"9da3d0b9",
         18179 => x"c6c5c2c1",
         18180 => x"c3c4bbbe",
         18181 => x"f0f0f0f0",
         18182 => x"f0f0f0f0",
         18183 => x"80818283",
         18184 => x"84f0f0f0",
         18185 => x"00000000",
         18186 => x"00000000",
         18187 => x"00000000",
         18188 => x"00000000",
         18189 => x"00000000",
         18190 => x"00000000",
         18191 => x"00000000",
         18192 => x"00000000",
         18193 => x"00000000",
         18194 => x"00000000",
         18195 => x"00000000",
         18196 => x"00000000",
         18197 => x"00000000",
         18198 => x"00000000",
         18199 => x"00000000",
         18200 => x"00000000",
         18201 => x"00000000",
         18202 => x"00000000",
         18203 => x"00000000",
         18204 => x"00000000",
         18205 => x"00000000",
         18206 => x"00000000",
         18207 => x"00000000",
         18208 => x"00000000",
         18209 => x"00000000",
         18210 => x"00010000",
         18211 => x"00000000",
         18212 => x"f8000000",
         18213 => x"0000f1ec",
         18214 => x"f3000000",
         18215 => x"0000f1f4",
         18216 => x"f4000000",
         18217 => x"0000f1f8",
         18218 => x"f1000000",
         18219 => x"0000f1fc",
         18220 => x"f2000000",
         18221 => x"0000f200",
         18222 => x"80000000",
         18223 => x"0000f204",
         18224 => x"81000000",
         18225 => x"0000f20c",
         18226 => x"82000000",
         18227 => x"0000f214",
         18228 => x"83000000",
         18229 => x"0000f21c",
         18230 => x"84000000",
         18231 => x"0000f224",
         18232 => x"85000000",
         18233 => x"0000f22c",
         18234 => x"86000000",
         18235 => x"0000f234",
         18236 => x"87000000",
         18237 => x"0000f23c",
         18238 => x"88000000",
         18239 => x"0000f244",
         18240 => x"89000000",
         18241 => x"0000f24c",
         18242 => x"f6000000",
         18243 => x"0000f254",
         18244 => x"7f000000",
         18245 => x"0000f25c",
         18246 => x"f9000000",
         18247 => x"0000f264",
         18248 => x"e0000000",
         18249 => x"0000f268",
         18250 => x"e1000000",
         18251 => x"0000f270",
         18252 => x"71000000",
         18253 => x"00000000",
         18254 => x"00000000",
         18255 => x"00000000",
         18256 => x"00000000",
         18257 => x"00000000",
         18258 => x"00000000",
         18259 => x"00000000",
         18260 => x"00000000",
         18261 => x"00000000",
         18262 => x"00000000",
         18263 => x"00000000",
         18264 => x"00000000",
         18265 => x"00000000",
         18266 => x"00000000",
         18267 => x"00000000",
         18268 => x"00000000",
         18269 => x"00000000",
         18270 => x"00000000",
         18271 => x"00000000",
         18272 => x"00000000",
         18273 => x"00000000",
         18274 => x"00000000",
         18275 => x"00000000",
         18276 => x"00000000",
         18277 => x"00000000",
         18278 => x"00000000",
         18279 => x"00000000",
         18280 => x"00000000",
         18281 => x"00000000",
         18282 => x"00000000",
         18283 => x"00000000",
         18284 => x"00000000",
         18285 => x"00000000",
         18286 => x"00000000",
         18287 => x"00000000",
         18288 => x"00000000",
         18289 => x"00000000",
         18290 => x"00000000",
         18291 => x"00000000",
         18292 => x"00000000",
         18293 => x"00000000",
         18294 => x"00000000",
         18295 => x"00000000",
         18296 => x"00000000",
         18297 => x"00000000",
         18298 => x"00000000",
         18299 => x"00000000",
         18300 => x"00000000",
         18301 => x"00000000",
         18302 => x"00000000",
         18303 => x"00000000",
         18304 => x"00000000",
         18305 => x"00000000",
         18306 => x"00000000",
         18307 => x"00000000",
         18308 => x"00000000",
         18309 => x"00000000",
         18310 => x"00000000",
         18311 => x"00000000",
         18312 => x"00000000",
         18313 => x"00000000",
         18314 => x"00000000",
         18315 => x"00000000",
         18316 => x"00000000",
         18317 => x"00000000",
         18318 => x"00000000",
         18319 => x"00000000",
         18320 => x"00000000",
         18321 => x"00000000",
         18322 => x"00000000",
         18323 => x"00000000",
         18324 => x"00000000",
         18325 => x"00000000",
         18326 => x"00000000",
         18327 => x"00000000",
         18328 => x"00000000",
         18329 => x"00000000",
         18330 => x"00000000",
         18331 => x"00000000",
         18332 => x"00000000",
         18333 => x"00000000",
         18334 => x"00000000",
         18335 => x"00000000",
         18336 => x"00000000",
         18337 => x"00000000",
         18338 => x"00000000",
         18339 => x"00000000",
         18340 => x"00000000",
         18341 => x"00000000",
         18342 => x"00000000",
         18343 => x"00000000",
         18344 => x"00000000",
         18345 => x"00000000",
         18346 => x"00000000",
         18347 => x"00000000",
         18348 => x"00000000",
         18349 => x"00000000",
         18350 => x"00000000",
         18351 => x"00000000",
         18352 => x"00000000",
         18353 => x"00000000",
         18354 => x"00000000",
         18355 => x"00000000",
         18356 => x"00000000",
         18357 => x"00000000",
         18358 => x"00000000",
         18359 => x"00000000",
         18360 => x"00000000",
         18361 => x"00000000",
         18362 => x"00000000",
         18363 => x"00000000",
         18364 => x"00000000",
         18365 => x"00000000",
         18366 => x"00000000",
         18367 => x"00000000",
         18368 => x"00000000",
         18369 => x"00000000",
         18370 => x"00000000",
         18371 => x"00000000",
         18372 => x"00000000",
         18373 => x"00000000",
         18374 => x"00000000",
         18375 => x"00000000",
         18376 => x"00000000",
         18377 => x"00000000",
         18378 => x"00000000",
         18379 => x"00000000",
         18380 => x"00000000",
         18381 => x"00000000",
         18382 => x"00000000",
         18383 => x"00000000",
         18384 => x"00000000",
         18385 => x"00000000",
         18386 => x"00000000",
         18387 => x"00000000",
         18388 => x"00000000",
         18389 => x"00000000",
         18390 => x"00000000",
         18391 => x"00000000",
         18392 => x"00000000",
         18393 => x"00000000",
         18394 => x"00000000",
         18395 => x"00000000",
         18396 => x"00000000",
         18397 => x"00000000",
         18398 => x"00000000",
         18399 => x"00000000",
         18400 => x"00000000",
         18401 => x"00000000",
         18402 => x"00000000",
         18403 => x"00000000",
         18404 => x"00000000",
         18405 => x"00000000",
         18406 => x"00000000",
         18407 => x"00000000",
         18408 => x"00000000",
         18409 => x"00000000",
         18410 => x"00000000",
         18411 => x"00000000",
         18412 => x"00000000",
         18413 => x"00000000",
         18414 => x"00000000",
         18415 => x"00000000",
         18416 => x"00000000",
         18417 => x"00000000",
         18418 => x"00000000",
         18419 => x"00000000",
         18420 => x"00000000",
         18421 => x"00000000",
         18422 => x"00000000",
         18423 => x"00000000",
         18424 => x"00000000",
         18425 => x"00000000",
         18426 => x"00000000",
         18427 => x"00000000",
         18428 => x"00000000",
         18429 => x"00000000",
         18430 => x"00000000",
         18431 => x"00000000",
         18432 => x"00000000",
         18433 => x"00000000",
         18434 => x"00000000",
         18435 => x"00000000",
         18436 => x"00000000",
         18437 => x"00000000",
         18438 => x"00000000",
         18439 => x"00000000",
         18440 => x"00000000",
         18441 => x"00000000",
         18442 => x"00000000",
         18443 => x"00000000",
         18444 => x"00000000",
         18445 => x"00000000",
         18446 => x"00000000",
         18447 => x"00000000",
         18448 => x"00000000",
         18449 => x"00000000",
         18450 => x"00000000",
         18451 => x"00000000",
         18452 => x"00000000",
         18453 => x"00000000",
         18454 => x"00000000",
         18455 => x"00000000",
         18456 => x"00000000",
         18457 => x"00000000",
         18458 => x"00000000",
         18459 => x"00000000",
         18460 => x"00000000",
         18461 => x"00000000",
         18462 => x"00000000",
         18463 => x"00000000",
         18464 => x"00000000",
         18465 => x"00000000",
         18466 => x"00000000",
         18467 => x"00000000",
         18468 => x"00000000",
         18469 => x"00000000",
         18470 => x"00000000",
         18471 => x"00000000",
         18472 => x"00000000",
         18473 => x"00000000",
         18474 => x"00000000",
         18475 => x"00000000",
         18476 => x"00000000",
         18477 => x"00000000",
         18478 => x"00000000",
         18479 => x"00000000",
         18480 => x"00000000",
         18481 => x"00000000",
         18482 => x"00000000",
         18483 => x"00000000",
         18484 => x"00000000",
         18485 => x"00000000",
         18486 => x"00000000",
         18487 => x"00000000",
         18488 => x"00000000",
         18489 => x"00000000",
         18490 => x"00000000",
         18491 => x"00000000",
         18492 => x"00000000",
         18493 => x"00000000",
         18494 => x"00000000",
         18495 => x"00000000",
         18496 => x"00000000",
         18497 => x"00000000",
         18498 => x"00000000",
         18499 => x"00000000",
         18500 => x"00000000",
         18501 => x"00000000",
         18502 => x"00000000",
         18503 => x"00000000",
         18504 => x"00000000",
         18505 => x"00000000",
         18506 => x"00000000",
         18507 => x"00000000",
         18508 => x"00000000",
         18509 => x"00000000",
         18510 => x"00000000",
         18511 => x"00000000",
         18512 => x"00000000",
         18513 => x"00000000",
         18514 => x"00000000",
         18515 => x"00000000",
         18516 => x"00000000",
         18517 => x"00000000",
         18518 => x"00000000",
         18519 => x"00000000",
         18520 => x"00000000",
         18521 => x"00000000",
         18522 => x"00000000",
         18523 => x"00000000",
         18524 => x"00000000",
         18525 => x"00000000",
         18526 => x"00000000",
         18527 => x"00000000",
         18528 => x"00000000",
         18529 => x"00000000",
         18530 => x"00000000",
         18531 => x"00000000",
         18532 => x"00000000",
         18533 => x"00000000",
         18534 => x"00000000",
         18535 => x"00000000",
         18536 => x"00000000",
         18537 => x"00000000",
         18538 => x"00000000",
         18539 => x"00000000",
         18540 => x"00000000",
         18541 => x"00000000",
         18542 => x"00000000",
         18543 => x"00000000",
         18544 => x"00000000",
         18545 => x"00000000",
         18546 => x"00000000",
         18547 => x"00000000",
         18548 => x"00000000",
         18549 => x"00000000",
         18550 => x"00000000",
         18551 => x"00000000",
         18552 => x"00000000",
         18553 => x"00000000",
         18554 => x"00000000",
         18555 => x"00000000",
         18556 => x"00000000",
         18557 => x"00000000",
         18558 => x"00000000",
         18559 => x"00000000",
         18560 => x"00000000",
         18561 => x"00000000",
         18562 => x"00000000",
         18563 => x"00000000",
         18564 => x"00000000",
         18565 => x"00000000",
         18566 => x"00000000",
         18567 => x"00000000",
         18568 => x"00000000",
         18569 => x"00000000",
         18570 => x"00000000",
         18571 => x"00000000",
         18572 => x"00000000",
         18573 => x"00000000",
         18574 => x"00000000",
         18575 => x"00000000",
         18576 => x"00000000",
         18577 => x"00000000",
         18578 => x"00000000",
         18579 => x"00000000",
         18580 => x"00000000",
         18581 => x"00000000",
         18582 => x"00000000",
         18583 => x"00000000",
         18584 => x"00000000",
         18585 => x"00000000",
         18586 => x"00000000",
         18587 => x"00000000",
         18588 => x"00000000",
         18589 => x"00000000",
         18590 => x"00000000",
         18591 => x"00000000",
         18592 => x"00000000",
         18593 => x"00000000",
         18594 => x"00000000",
         18595 => x"00000000",
         18596 => x"00000000",
         18597 => x"00000000",
         18598 => x"00000000",
         18599 => x"00000000",
         18600 => x"00000000",
         18601 => x"00000000",
         18602 => x"00000000",
         18603 => x"00000000",
         18604 => x"00000000",
         18605 => x"00000000",
         18606 => x"00000000",
         18607 => x"00000000",
         18608 => x"00000000",
         18609 => x"00000000",
         18610 => x"00000000",
         18611 => x"00000000",
         18612 => x"00000000",
         18613 => x"00000000",
         18614 => x"00000000",
         18615 => x"00000000",
         18616 => x"00000000",
         18617 => x"00000000",
         18618 => x"00000000",
         18619 => x"00000000",
         18620 => x"00000000",
         18621 => x"00000000",
         18622 => x"00000000",
         18623 => x"00000000",
         18624 => x"00000000",
         18625 => x"00000000",
         18626 => x"00000000",
         18627 => x"00000000",
         18628 => x"00000000",
         18629 => x"00000000",
         18630 => x"00000000",
         18631 => x"00000000",
         18632 => x"00000000",
         18633 => x"00000000",
         18634 => x"00000000",
         18635 => x"00000000",
         18636 => x"00000000",
         18637 => x"00000000",
         18638 => x"00000000",
         18639 => x"00000000",
         18640 => x"00000000",
         18641 => x"00000000",
         18642 => x"00000000",
         18643 => x"00000000",
         18644 => x"00000000",
         18645 => x"00000000",
         18646 => x"00000000",
         18647 => x"00000000",
         18648 => x"00000000",
         18649 => x"00000000",
         18650 => x"00000000",
         18651 => x"00000000",
         18652 => x"00000000",
         18653 => x"00000000",
         18654 => x"00000000",
         18655 => x"00000000",
         18656 => x"00000000",
         18657 => x"00000000",
         18658 => x"00000000",
         18659 => x"00000000",
         18660 => x"00000000",
         18661 => x"00000000",
         18662 => x"00000000",
         18663 => x"00000000",
         18664 => x"00000000",
         18665 => x"00000000",
         18666 => x"00000000",
         18667 => x"00000000",
         18668 => x"00000000",
         18669 => x"00000000",
         18670 => x"00000000",
         18671 => x"00000000",
         18672 => x"00000000",
         18673 => x"00000000",
         18674 => x"00000000",
         18675 => x"00000000",
         18676 => x"00000000",
         18677 => x"00000000",
         18678 => x"00000000",
         18679 => x"00000000",
         18680 => x"00000000",
         18681 => x"00000000",
         18682 => x"00000000",
         18683 => x"00000000",
         18684 => x"00000000",
         18685 => x"00000000",
         18686 => x"00000000",
         18687 => x"00000000",
         18688 => x"00000000",
         18689 => x"00000000",
         18690 => x"00000000",
         18691 => x"00000000",
         18692 => x"00000000",
         18693 => x"00000000",
         18694 => x"00000000",
         18695 => x"00000000",
         18696 => x"00000000",
         18697 => x"00000000",
         18698 => x"00000000",
         18699 => x"00000000",
         18700 => x"00000000",
         18701 => x"00000000",
         18702 => x"00000000",
         18703 => x"00000000",
         18704 => x"00000000",
         18705 => x"00000000",
         18706 => x"00000000",
         18707 => x"00000000",
         18708 => x"00000000",
         18709 => x"00000000",
         18710 => x"00000000",
         18711 => x"00000000",
         18712 => x"00000000",
         18713 => x"00000000",
         18714 => x"00000000",
         18715 => x"00000000",
         18716 => x"00000000",
         18717 => x"00000000",
         18718 => x"00000000",
         18719 => x"00000000",
         18720 => x"00000000",
         18721 => x"00000000",
         18722 => x"00000000",
         18723 => x"00000000",
         18724 => x"00000000",
         18725 => x"00000000",
         18726 => x"00000000",
         18727 => x"00000000",
         18728 => x"00000000",
         18729 => x"00000000",
         18730 => x"00000000",
         18731 => x"00000000",
         18732 => x"00000000",
         18733 => x"00000000",
         18734 => x"00000000",
         18735 => x"00000000",
         18736 => x"00000000",
         18737 => x"00000000",
         18738 => x"00000000",
         18739 => x"00000000",
         18740 => x"00000000",
         18741 => x"00000000",
         18742 => x"00000000",
         18743 => x"00000000",
         18744 => x"00000000",
         18745 => x"00000000",
         18746 => x"00000000",
         18747 => x"00000000",
         18748 => x"00000000",
         18749 => x"00000000",
         18750 => x"00000000",
         18751 => x"00000000",
         18752 => x"00000000",
         18753 => x"00000000",
         18754 => x"00000000",
         18755 => x"00000000",
         18756 => x"00000000",
         18757 => x"00000000",
         18758 => x"00000000",
         18759 => x"00000000",
         18760 => x"00000000",
         18761 => x"00000000",
         18762 => x"00000000",
         18763 => x"00000000",
         18764 => x"00000000",
         18765 => x"00000000",
         18766 => x"00000000",
         18767 => x"00000000",
         18768 => x"00000000",
         18769 => x"00000000",
         18770 => x"00000000",
         18771 => x"00000000",
         18772 => x"00000000",
         18773 => x"00000000",
         18774 => x"00000000",
         18775 => x"00000000",
         18776 => x"00000000",
         18777 => x"00000000",
         18778 => x"00000000",
         18779 => x"00000000",
         18780 => x"00000000",
         18781 => x"00000000",
         18782 => x"00000000",
         18783 => x"00000000",
         18784 => x"00000000",
         18785 => x"00000000",
         18786 => x"00000000",
         18787 => x"00000000",
         18788 => x"00000000",
         18789 => x"00000000",
         18790 => x"00000000",
         18791 => x"00000000",
         18792 => x"00000000",
         18793 => x"00000000",
         18794 => x"00000000",
         18795 => x"00000000",
         18796 => x"00000000",
         18797 => x"00000000",
         18798 => x"00000000",
         18799 => x"00000000",
         18800 => x"00000000",
         18801 => x"00000000",
         18802 => x"00000000",
         18803 => x"00000000",
         18804 => x"00000000",
         18805 => x"00000000",
         18806 => x"00000000",
         18807 => x"00000000",
         18808 => x"00000000",
         18809 => x"00000000",
         18810 => x"00000000",
         18811 => x"00000000",
         18812 => x"00000000",
         18813 => x"00000000",
         18814 => x"00000000",
         18815 => x"00000000",
         18816 => x"00000000",
         18817 => x"00000000",
         18818 => x"00000000",
         18819 => x"00000000",
         18820 => x"00000000",
         18821 => x"00000000",
         18822 => x"00000000",
         18823 => x"00000000",
         18824 => x"00000000",
         18825 => x"00000000",
         18826 => x"00000000",
         18827 => x"00000000",
         18828 => x"00000000",
         18829 => x"00000000",
         18830 => x"00000000",
         18831 => x"00000000",
         18832 => x"00000000",
         18833 => x"00000000",
         18834 => x"00000000",
         18835 => x"00000000",
         18836 => x"00000000",
         18837 => x"00000000",
         18838 => x"00000000",
         18839 => x"00000000",
         18840 => x"00000000",
         18841 => x"00000000",
         18842 => x"00000000",
         18843 => x"00000000",
         18844 => x"00000000",
         18845 => x"00000000",
         18846 => x"00000000",
         18847 => x"00000000",
         18848 => x"00000000",
         18849 => x"00000000",
         18850 => x"00000000",
         18851 => x"00000000",
         18852 => x"00000000",
         18853 => x"00000000",
         18854 => x"00000000",
         18855 => x"00000000",
         18856 => x"00000000",
         18857 => x"00000000",
         18858 => x"00000000",
         18859 => x"00000000",
         18860 => x"00000000",
         18861 => x"00000000",
         18862 => x"00000000",
         18863 => x"00000000",
         18864 => x"00000000",
         18865 => x"00000000",
         18866 => x"00000000",
         18867 => x"00000000",
         18868 => x"00000000",
         18869 => x"00000000",
         18870 => x"00000000",
         18871 => x"00000000",
         18872 => x"00000000",
         18873 => x"00000000",
         18874 => x"00000000",
         18875 => x"00000000",
         18876 => x"00000000",
         18877 => x"00000000",
         18878 => x"00000000",
         18879 => x"00000000",
         18880 => x"00000000",
         18881 => x"00000000",
         18882 => x"00000000",
         18883 => x"00000000",
         18884 => x"00000000",
         18885 => x"00000000",
         18886 => x"00000000",
         18887 => x"00000000",
         18888 => x"00000000",
         18889 => x"00000000",
         18890 => x"00000000",
         18891 => x"00000000",
         18892 => x"00000000",
         18893 => x"00000000",
         18894 => x"00000000",
         18895 => x"00000000",
         18896 => x"00000000",
         18897 => x"00000000",
         18898 => x"00000000",
         18899 => x"00000000",
         18900 => x"00000000",
         18901 => x"00000000",
         18902 => x"00000000",
         18903 => x"00000000",
         18904 => x"00000000",
         18905 => x"00000000",
         18906 => x"00000000",
         18907 => x"00000000",
         18908 => x"00000000",
         18909 => x"00000000",
         18910 => x"00000000",
         18911 => x"00000000",
         18912 => x"00000000",
         18913 => x"00000000",
         18914 => x"00000000",
         18915 => x"00000000",
         18916 => x"00000000",
         18917 => x"00000000",
         18918 => x"00000000",
         18919 => x"00000000",
         18920 => x"00000000",
         18921 => x"00000000",
         18922 => x"00000000",
         18923 => x"00000000",
         18924 => x"00000000",
         18925 => x"00000000",
         18926 => x"00000000",
         18927 => x"00000000",
         18928 => x"00000000",
         18929 => x"00000000",
         18930 => x"00000000",
         18931 => x"00000000",
         18932 => x"00000000",
         18933 => x"00000000",
         18934 => x"00000000",
         18935 => x"00000000",
         18936 => x"00000000",
         18937 => x"00000000",
         18938 => x"00000000",
         18939 => x"00000000",
         18940 => x"00000000",
         18941 => x"00000000",
         18942 => x"00000000",
         18943 => x"00000000",
         18944 => x"00000000",
         18945 => x"00000000",
         18946 => x"00000000",
         18947 => x"00000000",
         18948 => x"00000000",
         18949 => x"00000000",
         18950 => x"00000000",
         18951 => x"00000000",
         18952 => x"00000000",
         18953 => x"00000000",
         18954 => x"00000000",
         18955 => x"00000000",
         18956 => x"00000000",
         18957 => x"00000000",
         18958 => x"00000000",
         18959 => x"00000000",
         18960 => x"00000000",
         18961 => x"00000000",
         18962 => x"00000000",
         18963 => x"00000000",
         18964 => x"00000000",
         18965 => x"00000000",
         18966 => x"00000000",
         18967 => x"00000000",
         18968 => x"00000000",
         18969 => x"00000000",
         18970 => x"00000000",
         18971 => x"00000000",
         18972 => x"00000000",
         18973 => x"00000000",
         18974 => x"00000000",
         18975 => x"00000000",
         18976 => x"00000000",
         18977 => x"00000000",
         18978 => x"00000000",
         18979 => x"00000000",
         18980 => x"00000000",
         18981 => x"00000000",
         18982 => x"00000000",
         18983 => x"00000000",
         18984 => x"00000000",
         18985 => x"00000000",
         18986 => x"00000000",
         18987 => x"00000000",
         18988 => x"00000000",
         18989 => x"00000000",
         18990 => x"00000000",
         18991 => x"00000000",
         18992 => x"00000000",
         18993 => x"00000000",
         18994 => x"00000000",
         18995 => x"00000000",
         18996 => x"00000000",
         18997 => x"00000000",
         18998 => x"00000000",
         18999 => x"00000000",
         19000 => x"00000000",
         19001 => x"00000000",
         19002 => x"00000000",
         19003 => x"00000000",
         19004 => x"00000000",
         19005 => x"00000000",
         19006 => x"00000000",
         19007 => x"00000000",
         19008 => x"00000000",
         19009 => x"00000000",
         19010 => x"00000000",
         19011 => x"00000000",
         19012 => x"00000000",
         19013 => x"00000000",
         19014 => x"00000000",
         19015 => x"00000000",
         19016 => x"00000000",
         19017 => x"00000000",
         19018 => x"00000000",
         19019 => x"00000000",
         19020 => x"00000000",
         19021 => x"00000000",
         19022 => x"00000000",
         19023 => x"00000000",
         19024 => x"00000000",
         19025 => x"00000000",
         19026 => x"00000000",
         19027 => x"00000000",
         19028 => x"00000000",
         19029 => x"00000000",
         19030 => x"00000000",
         19031 => x"00000000",
         19032 => x"00000000",
         19033 => x"00000000",
         19034 => x"00000000",
         19035 => x"00000000",
         19036 => x"00000000",
         19037 => x"00000000",
         19038 => x"00000000",
         19039 => x"00000000",
         19040 => x"00000000",
         19041 => x"00000000",
         19042 => x"00000000",
         19043 => x"00000000",
         19044 => x"00000000",
         19045 => x"00000000",
         19046 => x"00000000",
         19047 => x"00000000",
         19048 => x"00000000",
         19049 => x"00000000",
         19050 => x"00000000",
         19051 => x"00000000",
         19052 => x"00000000",
         19053 => x"00000000",
         19054 => x"00000000",
         19055 => x"00000000",
         19056 => x"00000000",
         19057 => x"00000000",
         19058 => x"00000000",
         19059 => x"00000000",
         19060 => x"00000000",
         19061 => x"00000000",
         19062 => x"00000000",
         19063 => x"00000000",
         19064 => x"00000000",
         19065 => x"00000000",
         19066 => x"00000000",
         19067 => x"00000000",
         19068 => x"00000000",
         19069 => x"00000000",
         19070 => x"00000000",
         19071 => x"00000000",
         19072 => x"00000000",
         19073 => x"00000000",
         19074 => x"00000000",
         19075 => x"00000000",
         19076 => x"00000000",
         19077 => x"00000000",
         19078 => x"00000000",
         19079 => x"00000000",
         19080 => x"00000000",
         19081 => x"00000000",
         19082 => x"00000000",
         19083 => x"00000000",
         19084 => x"00000000",
         19085 => x"00000000",
         19086 => x"00000000",
         19087 => x"00000000",
         19088 => x"00000000",
         19089 => x"00000000",
         19090 => x"00000000",
         19091 => x"00000000",
         19092 => x"00000000",
         19093 => x"00000000",
         19094 => x"00000000",
         19095 => x"00000000",
         19096 => x"00000000",
         19097 => x"00000000",
         19098 => x"00000000",
         19099 => x"00000000",
         19100 => x"00000000",
         19101 => x"00000000",
         19102 => x"00000000",
         19103 => x"00000000",
         19104 => x"00000000",
         19105 => x"00000000",
         19106 => x"00000000",
         19107 => x"00000000",
         19108 => x"00000000",
         19109 => x"00000000",
         19110 => x"00000000",
         19111 => x"00000000",
         19112 => x"00000000",
         19113 => x"00000000",
         19114 => x"00000000",
         19115 => x"00000000",
         19116 => x"00000000",
         19117 => x"00000000",
         19118 => x"00000000",
         19119 => x"00000000",
         19120 => x"00000000",
         19121 => x"00000000",
         19122 => x"00000000",
         19123 => x"00000000",
         19124 => x"00000000",
         19125 => x"00000000",
         19126 => x"00000000",
         19127 => x"00000000",
         19128 => x"00000000",
         19129 => x"00000000",
         19130 => x"00000000",
         19131 => x"00000000",
         19132 => x"00000000",
         19133 => x"00000000",
         19134 => x"00000000",
         19135 => x"00000000",
         19136 => x"00000000",
         19137 => x"00000000",
         19138 => x"00000000",
         19139 => x"00000000",
         19140 => x"00000000",
         19141 => x"00000000",
         19142 => x"00000000",
         19143 => x"00000000",
         19144 => x"00000000",
         19145 => x"00000000",
         19146 => x"00000000",
         19147 => x"00000000",
         19148 => x"00000000",
         19149 => x"00000000",
         19150 => x"00000000",
         19151 => x"00000000",
         19152 => x"00000000",
         19153 => x"00000000",
         19154 => x"00000000",
         19155 => x"00000000",
         19156 => x"00000000",
         19157 => x"00000000",
         19158 => x"00000000",
         19159 => x"00000000",
         19160 => x"00000000",
         19161 => x"00000000",
         19162 => x"00000000",
         19163 => x"00000000",
         19164 => x"00000000",
         19165 => x"00000000",
         19166 => x"00000000",
         19167 => x"00000000",
         19168 => x"00000000",
         19169 => x"00000000",
         19170 => x"00000000",
         19171 => x"00000000",
         19172 => x"00000000",
         19173 => x"00000000",
         19174 => x"00000000",
         19175 => x"00000000",
         19176 => x"00000000",
         19177 => x"00000000",
         19178 => x"00000000",
         19179 => x"00000000",
         19180 => x"00000000",
         19181 => x"00000000",
         19182 => x"00000000",
         19183 => x"00000000",
         19184 => x"00000000",
         19185 => x"00000000",
         19186 => x"00000000",
         19187 => x"00000000",
         19188 => x"00000000",
         19189 => x"00000000",
         19190 => x"00000000",
         19191 => x"00000000",
         19192 => x"00000000",
         19193 => x"00000000",
         19194 => x"00000000",
         19195 => x"00000000",
         19196 => x"00000000",
         19197 => x"00000000",
         19198 => x"00000000",
         19199 => x"00000000",
         19200 => x"00000000",
         19201 => x"00000000",
         19202 => x"00000000",
         19203 => x"00000000",
         19204 => x"00000000",
         19205 => x"00000000",
         19206 => x"00000000",
         19207 => x"00000000",
         19208 => x"00000000",
         19209 => x"00000000",
         19210 => x"00000000",
         19211 => x"00000000",
         19212 => x"00000000",
         19213 => x"00000000",
         19214 => x"00000000",
         19215 => x"00000000",
         19216 => x"00000000",
         19217 => x"00000000",
         19218 => x"00000000",
         19219 => x"00000000",
         19220 => x"00000000",
         19221 => x"00000000",
         19222 => x"00000000",
         19223 => x"00000000",
         19224 => x"00000000",
         19225 => x"00000000",
         19226 => x"00000000",
         19227 => x"00000000",
         19228 => x"00000000",
         19229 => x"00000000",
         19230 => x"00000000",
         19231 => x"00000000",
         19232 => x"00000000",
         19233 => x"00000000",
         19234 => x"00000000",
         19235 => x"00000000",
         19236 => x"00000000",
         19237 => x"00000000",
         19238 => x"00000000",
         19239 => x"00000000",
         19240 => x"00000000",
         19241 => x"00000000",
         19242 => x"00000000",
         19243 => x"00000000",
         19244 => x"00000000",
         19245 => x"00000000",
         19246 => x"00000000",
         19247 => x"00000000",
         19248 => x"00000000",
         19249 => x"00000000",
         19250 => x"00000000",
         19251 => x"00000000",
         19252 => x"00000000",
         19253 => x"00000000",
         19254 => x"00000000",
         19255 => x"00000000",
         19256 => x"00000000",
         19257 => x"00000000",
         19258 => x"00000000",
         19259 => x"00000000",
         19260 => x"00000000",
         19261 => x"00000000",
         19262 => x"00000000",
         19263 => x"00000000",
         19264 => x"00000000",
         19265 => x"00000000",
         19266 => x"00000000",
         19267 => x"00000000",
         19268 => x"00000000",
         19269 => x"00000000",
         19270 => x"00000000",
         19271 => x"00000000",
         19272 => x"00000000",
         19273 => x"00000000",
         19274 => x"00000000",
         19275 => x"00000000",
         19276 => x"00000000",
         19277 => x"00000000",
         19278 => x"00000000",
         19279 => x"00000000",
         19280 => x"00000000",
         19281 => x"00000000",
         19282 => x"00000000",
         19283 => x"00000000",
         19284 => x"00000000",
         19285 => x"00000000",
         19286 => x"00000000",
         19287 => x"00000000",
         19288 => x"00000000",
         19289 => x"00000000",
         19290 => x"00000000",
         19291 => x"00000000",
         19292 => x"00000000",
         19293 => x"00000000",
         19294 => x"00000000",
         19295 => x"00000000",
         19296 => x"00000000",
         19297 => x"00000000",
         19298 => x"00000000",
         19299 => x"00000000",
         19300 => x"00000000",
         19301 => x"00000000",
         19302 => x"00000000",
         19303 => x"00000000",
         19304 => x"00000000",
         19305 => x"00000000",
         19306 => x"00000000",
         19307 => x"00000000",
         19308 => x"00000000",
         19309 => x"00000000",
         19310 => x"00000000",
         19311 => x"00000000",
         19312 => x"00000000",
         19313 => x"00000000",
         19314 => x"00000000",
         19315 => x"00000000",
         19316 => x"00000000",
         19317 => x"00000000",
         19318 => x"00000000",
         19319 => x"00000000",
         19320 => x"00000000",
         19321 => x"00000000",
         19322 => x"00000000",
         19323 => x"00000000",
         19324 => x"00000000",
         19325 => x"00000000",
         19326 => x"00000000",
         19327 => x"00000000",
         19328 => x"00000000",
         19329 => x"00000000",
         19330 => x"00000000",
         19331 => x"00000000",
         19332 => x"00000000",
         19333 => x"00000000",
         19334 => x"00000000",
         19335 => x"00000000",
         19336 => x"00000000",
         19337 => x"00000000",
         19338 => x"00000000",
         19339 => x"00000000",
         19340 => x"00000000",
         19341 => x"00000000",
         19342 => x"00000000",
         19343 => x"00000000",
         19344 => x"00000000",
         19345 => x"00000000",
         19346 => x"00000000",
         19347 => x"00000000",
         19348 => x"00000000",
         19349 => x"00000000",
         19350 => x"00000000",
         19351 => x"00000000",
         19352 => x"00000000",
         19353 => x"00000000",
         19354 => x"00000000",
         19355 => x"00000000",
         19356 => x"00000000",
         19357 => x"00000000",
         19358 => x"00000000",
         19359 => x"00000000",
         19360 => x"00000000",
         19361 => x"00000000",
         19362 => x"00000000",
         19363 => x"00000000",
         19364 => x"00000000",
         19365 => x"00000000",
         19366 => x"00000000",
         19367 => x"00000000",
         19368 => x"00000000",
         19369 => x"00000000",
         19370 => x"00000000",
         19371 => x"00000000",
         19372 => x"00000000",
         19373 => x"00000000",
         19374 => x"00000000",
         19375 => x"00000000",
         19376 => x"00000000",
         19377 => x"00000000",
         19378 => x"00000000",
         19379 => x"00000000",
         19380 => x"00000000",
         19381 => x"00000000",
         19382 => x"00000000",
         19383 => x"00000000",
         19384 => x"00000000",
         19385 => x"00000000",
         19386 => x"00000000",
         19387 => x"00000000",
         19388 => x"00000000",
         19389 => x"00000000",
         19390 => x"00000000",
         19391 => x"00000000",
         19392 => x"00000000",
         19393 => x"00000000",
         19394 => x"00000000",
         19395 => x"00000000",
         19396 => x"00000000",
         19397 => x"00000000",
         19398 => x"00000000",
         19399 => x"00000000",
         19400 => x"00000000",
         19401 => x"00000000",
         19402 => x"00000000",
         19403 => x"00000000",
         19404 => x"00000000",
         19405 => x"00000000",
         19406 => x"00000000",
         19407 => x"00000000",
         19408 => x"00000000",
         19409 => x"00000000",
         19410 => x"00000000",
         19411 => x"00000000",
         19412 => x"00000000",
         19413 => x"00000000",
         19414 => x"00000000",
         19415 => x"00000000",
         19416 => x"00000000",
         19417 => x"00000000",
         19418 => x"00000000",
         19419 => x"00000000",
         19420 => x"00000000",
         19421 => x"00000000",
         19422 => x"00000000",
         19423 => x"00000000",
         19424 => x"00000000",
         19425 => x"00000000",
         19426 => x"00000000",
         19427 => x"00000000",
         19428 => x"00000000",
         19429 => x"00000000",
         19430 => x"00000000",
         19431 => x"00000000",
         19432 => x"00000000",
         19433 => x"00000000",
         19434 => x"00000000",
         19435 => x"00000000",
         19436 => x"00000000",
         19437 => x"00000000",
         19438 => x"00000000",
         19439 => x"00000000",
         19440 => x"00000000",
         19441 => x"00000000",
         19442 => x"00000000",
         19443 => x"00000000",
         19444 => x"00000000",
         19445 => x"00000000",
         19446 => x"00000000",
         19447 => x"00000000",
         19448 => x"00000000",
         19449 => x"00000000",
         19450 => x"00000000",
         19451 => x"00000000",
         19452 => x"00000000",
         19453 => x"00000000",
         19454 => x"00000000",
         19455 => x"00000000",
         19456 => x"00000000",
         19457 => x"00000000",
         19458 => x"00000000",
         19459 => x"00000000",
         19460 => x"00000000",
         19461 => x"00000000",
         19462 => x"00000000",
         19463 => x"00000000",
         19464 => x"00000000",
         19465 => x"00000000",
         19466 => x"00000000",
         19467 => x"00000000",
         19468 => x"00000000",
         19469 => x"00000000",
         19470 => x"00000000",
         19471 => x"00000000",
         19472 => x"00000000",
         19473 => x"00000000",
         19474 => x"00000000",
         19475 => x"00000000",
         19476 => x"00000000",
         19477 => x"00000000",
         19478 => x"00000000",
         19479 => x"00000000",
         19480 => x"00000000",
         19481 => x"00000000",
         19482 => x"00000000",
         19483 => x"00000000",
         19484 => x"00000000",
         19485 => x"00000000",
         19486 => x"00000000",
         19487 => x"00000000",
         19488 => x"00000000",
         19489 => x"00000000",
         19490 => x"00000000",
         19491 => x"00000000",
         19492 => x"00000000",
         19493 => x"00000000",
         19494 => x"00000000",
         19495 => x"00000000",
         19496 => x"00000000",
         19497 => x"00000000",
         19498 => x"00000000",
         19499 => x"00000000",
         19500 => x"00000000",
         19501 => x"00000000",
         19502 => x"00000000",
         19503 => x"00000000",
         19504 => x"00000000",
         19505 => x"00000000",
         19506 => x"00000000",
         19507 => x"00000000",
         19508 => x"00000000",
         19509 => x"00000000",
         19510 => x"00000000",
         19511 => x"00000000",
         19512 => x"00000000",
         19513 => x"00000000",
         19514 => x"00000000",
         19515 => x"00000000",
         19516 => x"00000000",
         19517 => x"00000000",
         19518 => x"00000000",
         19519 => x"00000000",
         19520 => x"00000000",
         19521 => x"00000000",
         19522 => x"00000000",
         19523 => x"00000000",
         19524 => x"00000000",
         19525 => x"00000000",
         19526 => x"00000000",
         19527 => x"00000000",
         19528 => x"00000000",
         19529 => x"00000000",
         19530 => x"00000000",
         19531 => x"00000000",
         19532 => x"00000000",
         19533 => x"00000000",
         19534 => x"00000000",
         19535 => x"00000000",
         19536 => x"00000000",
         19537 => x"00000000",
         19538 => x"00000000",
         19539 => x"00000000",
         19540 => x"00000000",
         19541 => x"00000000",
         19542 => x"00000000",
         19543 => x"00000000",
         19544 => x"00000000",
         19545 => x"00000000",
         19546 => x"00000000",
         19547 => x"00000000",
         19548 => x"00000000",
         19549 => x"00000000",
         19550 => x"00000000",
         19551 => x"00000000",
         19552 => x"00000000",
         19553 => x"00000000",
         19554 => x"00000000",
         19555 => x"00000000",
         19556 => x"00000000",
         19557 => x"00000000",
         19558 => x"00000000",
         19559 => x"00000000",
         19560 => x"00000000",
         19561 => x"00000000",
         19562 => x"00000000",
         19563 => x"00000000",
         19564 => x"00000000",
         19565 => x"00000000",
         19566 => x"00000000",
         19567 => x"00000000",
         19568 => x"00000000",
         19569 => x"00000000",
         19570 => x"00000000",
         19571 => x"00000000",
         19572 => x"00000000",
         19573 => x"00000000",
         19574 => x"00000000",
         19575 => x"00000000",
         19576 => x"00000000",
         19577 => x"00000000",
         19578 => x"00000000",
         19579 => x"00000000",
         19580 => x"00000000",
         19581 => x"00000000",
         19582 => x"00000000",
         19583 => x"00000000",
         19584 => x"00000000",
         19585 => x"00000000",
         19586 => x"00000000",
         19587 => x"00000000",
         19588 => x"00000000",
         19589 => x"00000000",
         19590 => x"00000000",
         19591 => x"00000000",
         19592 => x"00000000",
         19593 => x"00000000",
         19594 => x"00000000",
         19595 => x"00000000",
         19596 => x"00000000",
         19597 => x"00000000",
         19598 => x"00000000",
         19599 => x"00000000",
         19600 => x"00000000",
         19601 => x"00000000",
         19602 => x"00000000",
         19603 => x"00000000",
         19604 => x"00000000",
         19605 => x"00000000",
         19606 => x"00000000",
         19607 => x"00000000",
         19608 => x"00000000",
         19609 => x"00000000",
         19610 => x"00000000",
         19611 => x"00000000",
         19612 => x"00000000",
         19613 => x"00000000",
         19614 => x"00000000",
         19615 => x"00000000",
         19616 => x"00000000",
         19617 => x"00000000",
         19618 => x"00000000",
         19619 => x"00000000",
         19620 => x"00000000",
         19621 => x"00000000",
         19622 => x"00000000",
         19623 => x"00000000",
         19624 => x"00000000",
         19625 => x"00000000",
         19626 => x"00000000",
         19627 => x"00000000",
         19628 => x"00000000",
         19629 => x"00000000",
         19630 => x"00000000",
         19631 => x"00000000",
         19632 => x"00000000",
         19633 => x"00000000",
         19634 => x"00000000",
         19635 => x"00000000",
         19636 => x"00000000",
         19637 => x"00000000",
         19638 => x"00000000",
         19639 => x"00000000",
         19640 => x"00000000",
         19641 => x"00000000",
         19642 => x"00000000",
         19643 => x"00000000",
         19644 => x"00000000",
         19645 => x"00000000",
         19646 => x"00000000",
         19647 => x"00000000",
         19648 => x"00000000",
         19649 => x"00000000",
         19650 => x"00000000",
         19651 => x"00000000",
         19652 => x"00000000",
         19653 => x"00000000",
         19654 => x"00000000",
         19655 => x"00000000",
         19656 => x"00000000",
         19657 => x"00000000",
         19658 => x"00000000",
         19659 => x"00000000",
         19660 => x"00000000",
         19661 => x"00000000",
         19662 => x"00000000",
         19663 => x"00000000",
         19664 => x"00000000",
         19665 => x"00000000",
         19666 => x"00000000",
         19667 => x"00000000",
         19668 => x"00000000",
         19669 => x"00000000",
         19670 => x"00000000",
         19671 => x"00000000",
         19672 => x"00000000",
         19673 => x"00000000",
         19674 => x"00000000",
         19675 => x"00000000",
         19676 => x"00000000",
         19677 => x"00000000",
         19678 => x"00000000",
         19679 => x"00000000",
         19680 => x"00000000",
         19681 => x"00000000",
         19682 => x"00000000",
         19683 => x"00000000",
         19684 => x"00000000",
         19685 => x"00000000",
         19686 => x"00000000",
         19687 => x"00000000",
         19688 => x"00000000",
         19689 => x"00000000",
         19690 => x"00000000",
         19691 => x"00000000",
         19692 => x"00000000",
         19693 => x"00000000",
         19694 => x"00000000",
         19695 => x"00000000",
         19696 => x"00000000",
         19697 => x"00000000",
         19698 => x"00000000",
         19699 => x"00000000",
         19700 => x"00000000",
         19701 => x"00000000",
         19702 => x"00000000",
         19703 => x"00000000",
         19704 => x"00000000",
         19705 => x"00000000",
         19706 => x"00000000",
         19707 => x"00000000",
         19708 => x"00000000",
         19709 => x"00000000",
         19710 => x"00000000",
         19711 => x"00000000",
         19712 => x"00000000",
         19713 => x"00000000",
         19714 => x"00000000",
         19715 => x"00000000",
         19716 => x"00000000",
         19717 => x"00000000",
         19718 => x"00000000",
         19719 => x"00000000",
         19720 => x"00000000",
         19721 => x"00000000",
         19722 => x"00000000",
         19723 => x"00000000",
         19724 => x"00000000",
         19725 => x"00000000",
         19726 => x"00000000",
         19727 => x"00000000",
         19728 => x"00000000",
         19729 => x"00000000",
         19730 => x"00000000",
         19731 => x"00000000",
         19732 => x"00000000",
         19733 => x"00000000",
         19734 => x"00000000",
         19735 => x"00000000",
         19736 => x"00000000",
         19737 => x"00000000",
         19738 => x"00000000",
         19739 => x"00000000",
         19740 => x"00000000",
         19741 => x"00000000",
         19742 => x"00000000",
         19743 => x"00000000",
         19744 => x"00000000",
         19745 => x"00000000",
         19746 => x"00000000",
         19747 => x"00000000",
         19748 => x"00000000",
         19749 => x"00000000",
         19750 => x"00000000",
         19751 => x"00000000",
         19752 => x"00000000",
         19753 => x"00000000",
         19754 => x"00000000",
         19755 => x"00000000",
         19756 => x"00000000",
         19757 => x"00000000",
         19758 => x"00000000",
         19759 => x"00000000",
         19760 => x"00000000",
         19761 => x"00000000",
         19762 => x"00000000",
         19763 => x"00000000",
         19764 => x"00000000",
         19765 => x"00000000",
         19766 => x"00000000",
         19767 => x"00000000",
         19768 => x"00000000",
         19769 => x"00000000",
         19770 => x"00000000",
         19771 => x"00000000",
         19772 => x"00000000",
         19773 => x"00000000",
         19774 => x"00000000",
         19775 => x"00000000",
         19776 => x"00000000",
         19777 => x"00000000",
         19778 => x"00000000",
         19779 => x"00000000",
         19780 => x"00000000",
         19781 => x"00000000",
         19782 => x"00000000",
         19783 => x"00000000",
         19784 => x"00000000",
         19785 => x"00000000",
         19786 => x"00000000",
         19787 => x"00000000",
         19788 => x"00000000",
         19789 => x"00000000",
         19790 => x"00000000",
         19791 => x"00000000",
         19792 => x"00000000",
         19793 => x"00000000",
         19794 => x"00000000",
         19795 => x"00000000",
         19796 => x"00000000",
         19797 => x"00000000",
         19798 => x"00000000",
         19799 => x"00000000",
         19800 => x"00000000",
         19801 => x"00000000",
         19802 => x"00000000",
         19803 => x"00000000",
         19804 => x"00000000",
         19805 => x"00000000",
         19806 => x"00000000",
         19807 => x"00000000",
         19808 => x"00000000",
         19809 => x"00000000",
         19810 => x"00000000",
         19811 => x"00000000",
         19812 => x"00000000",
         19813 => x"00000000",
         19814 => x"00000000",
         19815 => x"00000000",
         19816 => x"00000000",
         19817 => x"00000000",
         19818 => x"00000000",
         19819 => x"00000000",
         19820 => x"00000000",
         19821 => x"00000000",
         19822 => x"00000000",
         19823 => x"00000000",
         19824 => x"00000000",
         19825 => x"00000000",
         19826 => x"00000000",
         19827 => x"00000000",
         19828 => x"00000000",
         19829 => x"00000000",
         19830 => x"00000000",
         19831 => x"00000000",
         19832 => x"00000000",
         19833 => x"00000000",
         19834 => x"00000000",
         19835 => x"00000000",
         19836 => x"00000000",
         19837 => x"00000000",
         19838 => x"00000000",
         19839 => x"00000000",
         19840 => x"00000000",
         19841 => x"00000000",
         19842 => x"00000000",
         19843 => x"00000000",
         19844 => x"00000000",
         19845 => x"00000000",
         19846 => x"00000000",
         19847 => x"00000000",
         19848 => x"00000000",
         19849 => x"00000000",
         19850 => x"00000000",
         19851 => x"00000000",
         19852 => x"00000000",
         19853 => x"00000000",
         19854 => x"00000000",
         19855 => x"00000000",
         19856 => x"00000000",
         19857 => x"00000000",
         19858 => x"00000000",
         19859 => x"00000000",
         19860 => x"00000000",
         19861 => x"00000000",
         19862 => x"00000000",
         19863 => x"00000000",
         19864 => x"00000000",
         19865 => x"00000000",
         19866 => x"00000000",
         19867 => x"00000000",
         19868 => x"00000000",
         19869 => x"00000000",
         19870 => x"00000000",
         19871 => x"00000000",
         19872 => x"00000000",
         19873 => x"00000000",
         19874 => x"00000000",
         19875 => x"00000000",
         19876 => x"00000000",
         19877 => x"00000000",
         19878 => x"00000000",
         19879 => x"00000000",
         19880 => x"00000000",
         19881 => x"00000000",
         19882 => x"00000000",
         19883 => x"00000000",
         19884 => x"00000000",
         19885 => x"00000000",
         19886 => x"00000000",
         19887 => x"00000000",
         19888 => x"00000000",
         19889 => x"00000000",
         19890 => x"00000000",
         19891 => x"00000000",
         19892 => x"00000000",
         19893 => x"00000000",
         19894 => x"00000000",
         19895 => x"00000000",
         19896 => x"00000000",
         19897 => x"00000000",
         19898 => x"00000000",
         19899 => x"00000000",
         19900 => x"00000000",
         19901 => x"00000000",
         19902 => x"00000000",
         19903 => x"00000000",
         19904 => x"00000000",
         19905 => x"00000000",
         19906 => x"00000000",
         19907 => x"00000000",
         19908 => x"00000000",
         19909 => x"00000000",
         19910 => x"00000000",
         19911 => x"00000000",
         19912 => x"00000000",
         19913 => x"00000000",
         19914 => x"00000000",
         19915 => x"00000000",
         19916 => x"00000000",
         19917 => x"00000000",
         19918 => x"00000000",
         19919 => x"00000000",
         19920 => x"00000000",
         19921 => x"00000000",
         19922 => x"00000000",
         19923 => x"00000000",
         19924 => x"00000000",
         19925 => x"00000000",
         19926 => x"00000000",
         19927 => x"00000000",
         19928 => x"00000000",
         19929 => x"00000000",
         19930 => x"00000000",
         19931 => x"00000000",
         19932 => x"00000000",
         19933 => x"00000000",
         19934 => x"00000000",
         19935 => x"00000000",
         19936 => x"00000000",
         19937 => x"00000000",
         19938 => x"00000000",
         19939 => x"00000000",
         19940 => x"00000000",
         19941 => x"00000000",
         19942 => x"00000000",
         19943 => x"00000000",
         19944 => x"00000000",
         19945 => x"00000000",
         19946 => x"00000000",
         19947 => x"00000000",
         19948 => x"00000000",
         19949 => x"00000000",
         19950 => x"00000000",
         19951 => x"00000000",
         19952 => x"00000000",
         19953 => x"00000000",
         19954 => x"00000000",
         19955 => x"00000000",
         19956 => x"00000000",
         19957 => x"00000000",
         19958 => x"00000000",
         19959 => x"00000000",
         19960 => x"00000000",
         19961 => x"00000000",
         19962 => x"00000000",
         19963 => x"00000000",
         19964 => x"00000000",
         19965 => x"00000000",
         19966 => x"00000000",
         19967 => x"00000000",
         19968 => x"00000000",
         19969 => x"00000000",
         19970 => x"00000000",
         19971 => x"00000000",
         19972 => x"00000000",
         19973 => x"00000000",
         19974 => x"00000000",
         19975 => x"00000000",
         19976 => x"00000000",
         19977 => x"00000000",
         19978 => x"00000000",
         19979 => x"00000000",
         19980 => x"00000000",
         19981 => x"00000000",
         19982 => x"00000000",
         19983 => x"00000000",
         19984 => x"00000000",
         19985 => x"00000000",
         19986 => x"00000000",
         19987 => x"00000000",
         19988 => x"00000000",
         19989 => x"00000000",
         19990 => x"00000000",
         19991 => x"00000000",
         19992 => x"00000000",
         19993 => x"00000000",
         19994 => x"00000000",
         19995 => x"00000000",
         19996 => x"00000000",
         19997 => x"00000000",
         19998 => x"00000000",
         19999 => x"00000000",
         20000 => x"00000000",
         20001 => x"00000000",
         20002 => x"00000000",
         20003 => x"00000000",
         20004 => x"00000000",
         20005 => x"00000000",
         20006 => x"00000000",
         20007 => x"00000000",
         20008 => x"00000000",
         20009 => x"00000000",
         20010 => x"00000000",
         20011 => x"00000000",
         20012 => x"00000000",
         20013 => x"00000000",
         20014 => x"00000000",
         20015 => x"00000000",
         20016 => x"00000000",
         20017 => x"00000000",
         20018 => x"00000000",
         20019 => x"00000000",
         20020 => x"00000000",
         20021 => x"00000000",
         20022 => x"00000000",
         20023 => x"00000000",
         20024 => x"00000000",
         20025 => x"00000000",
         20026 => x"00000000",
         20027 => x"00000000",
         20028 => x"00000000",
         20029 => x"00000000",
         20030 => x"00000000",
         20031 => x"00000000",
         20032 => x"00000000",
         20033 => x"00000000",
         20034 => x"00000000",
         20035 => x"00000000",
         20036 => x"00000000",
         20037 => x"00000000",
         20038 => x"00000000",
         20039 => x"00000000",
         20040 => x"00000000",
         20041 => x"00000000",
         20042 => x"00000000",
         20043 => x"00000000",
         20044 => x"00000000",
         20045 => x"00000000",
         20046 => x"00000000",
         20047 => x"00000000",
         20048 => x"00000000",
         20049 => x"00000000",
         20050 => x"00000000",
         20051 => x"00000000",
         20052 => x"00000000",
         20053 => x"00000000",
         20054 => x"00000000",
         20055 => x"00000000",
         20056 => x"00000000",
         20057 => x"00000000",
         20058 => x"00000000",
         20059 => x"00000000",
         20060 => x"00000000",
         20061 => x"00000000",
         20062 => x"00000000",
         20063 => x"00000000",
         20064 => x"00000000",
         20065 => x"00000000",
         20066 => x"00000000",
         20067 => x"00000000",
         20068 => x"00000000",
         20069 => x"00000000",
         20070 => x"00000000",
         20071 => x"00000000",
         20072 => x"00000000",
         20073 => x"00000000",
         20074 => x"00000000",
         20075 => x"00000000",
         20076 => x"00000000",
         20077 => x"00000000",
         20078 => x"00000000",
         20079 => x"00000000",
         20080 => x"00000000",
         20081 => x"00000000",
         20082 => x"00000000",
         20083 => x"00000000",
         20084 => x"00000000",
         20085 => x"00000000",
         20086 => x"00000000",
         20087 => x"00000000",
         20088 => x"00000000",
         20089 => x"00000000",
         20090 => x"00000000",
         20091 => x"00000000",
         20092 => x"00000000",
         20093 => x"00000000",
         20094 => x"00000000",
         20095 => x"00000000",
         20096 => x"00000000",
         20097 => x"00000000",
         20098 => x"00000000",
         20099 => x"00000000",
         20100 => x"00000000",
         20101 => x"00000000",
         20102 => x"00000000",
         20103 => x"00000000",
         20104 => x"00000000",
         20105 => x"00000000",
         20106 => x"00000000",
         20107 => x"00000000",
         20108 => x"00000000",
         20109 => x"00000000",
         20110 => x"00000000",
         20111 => x"00000000",
         20112 => x"00000000",
         20113 => x"00000000",
         20114 => x"00000000",
         20115 => x"00000000",
         20116 => x"00000000",
         20117 => x"00000000",
         20118 => x"00000000",
         20119 => x"00000000",
         20120 => x"00000000",
         20121 => x"00000000",
         20122 => x"00000000",
         20123 => x"00000000",
         20124 => x"00000000",
         20125 => x"00000000",
         20126 => x"00000000",
         20127 => x"00000000",
         20128 => x"00000000",
         20129 => x"00000000",
         20130 => x"00000000",
         20131 => x"00000000",
         20132 => x"00000000",
         20133 => x"00000000",
         20134 => x"00000000",
         20135 => x"00000000",
         20136 => x"00000000",
         20137 => x"00000000",
         20138 => x"00000000",
         20139 => x"00000000",
         20140 => x"00000000",
         20141 => x"00000000",
         20142 => x"00000000",
         20143 => x"00000000",
         20144 => x"00000000",
         20145 => x"00000000",
         20146 => x"00000000",
         20147 => x"00000000",
         20148 => x"00000000",
         20149 => x"00000000",
         20150 => x"00000000",
         20151 => x"00000000",
         20152 => x"00000000",
         20153 => x"00000000",
         20154 => x"00000000",
         20155 => x"00000000",
         20156 => x"00000000",
         20157 => x"00000000",
         20158 => x"00000000",
         20159 => x"00000000",
         20160 => x"00000000",
         20161 => x"00000000",
         20162 => x"00000000",
         20163 => x"00000000",
         20164 => x"00000000",
         20165 => x"00000000",
         20166 => x"00000000",
         20167 => x"00000000",
         20168 => x"00000000",
         20169 => x"00000000",
         20170 => x"00000000",
         20171 => x"00000000",
         20172 => x"00000000",
         20173 => x"00000000",
         20174 => x"00000000",
         20175 => x"00000000",
         20176 => x"00000000",
         20177 => x"00000000",
         20178 => x"00000000",
         20179 => x"00000000",
         20180 => x"00000000",
         20181 => x"00000000",
         20182 => x"00000000",
         20183 => x"00000000",
         20184 => x"00000000",
         20185 => x"00000000",
         20186 => x"00000000",
         20187 => x"00000000",
         20188 => x"00000000",
         20189 => x"00000000",
         20190 => x"00000000",
         20191 => x"00000000",
         20192 => x"00000000",
         20193 => x"00000000",
         20194 => x"00000000",
         20195 => x"00000000",
         20196 => x"00000000",
         20197 => x"00000000",
         20198 => x"00000000",
         20199 => x"00000000",
         20200 => x"00000000",
         20201 => x"00000000",
         20202 => x"00000000",
         20203 => x"00000000",
         20204 => x"00000000",
         20205 => x"00000000",
         20206 => x"00000000",
         20207 => x"00000000",
         20208 => x"00000000",
         20209 => x"00000000",
         20210 => x"00000000",
         20211 => x"00000000",
         20212 => x"00000000",
         20213 => x"00000000",
         20214 => x"00000000",
         20215 => x"00000000",
         20216 => x"00000000",
         20217 => x"00000000",
         20218 => x"00000000",
         20219 => x"00000000",
         20220 => x"00000000",
         20221 => x"00000000",
         20222 => x"00000000",
         20223 => x"00000000",
         20224 => x"00000000",
         20225 => x"00000000",
         20226 => x"00000000",
         20227 => x"00000000",
         20228 => x"00000000",
         20229 => x"00000000",
         20230 => x"00000000",
         20231 => x"00000000",
         20232 => x"00000000",
         20233 => x"00000000",
         20234 => x"00000000",
         20235 => x"00000000",
         20236 => x"00000000",
         20237 => x"00000000",
         20238 => x"00000000",
         20239 => x"00000000",
         20240 => x"00000000",
         20241 => x"00000000",
         20242 => x"00000000",
         20243 => x"00000000",
         20244 => x"00000000",
         20245 => x"00000000",
         20246 => x"00000000",
         20247 => x"00000000",
         20248 => x"00000000",
         20249 => x"00000000",
         20250 => x"00000000",
         20251 => x"00000000",
         20252 => x"00000000",
         20253 => x"00003219",
         20254 => x"50000100",
         20255 => x"00000000",
         20256 => x"cce0f2f3",
         20257 => x"cecff6f7",
         20258 => x"f8f9fafb",
         20259 => x"fcfdfeff",
         20260 => x"e1c1c2c3",
         20261 => x"c4c5c6e2",
         20262 => x"e3e4e5e6",
         20263 => x"ebeeeff4",
         20264 => x"00616263",
         20265 => x"64656667",
         20266 => x"68696b6a",
         20267 => x"2f2a2e2d",
         20268 => x"20212223",
         20269 => x"24252627",
         20270 => x"28294f2c",
         20271 => x"512b5749",
         20272 => x"55010203",
         20273 => x"04050607",
         20274 => x"08090a0b",
         20275 => x"0c0d0e0f",
         20276 => x"10111213",
         20277 => x"14151617",
         20278 => x"18191a52",
         20279 => x"5954be3c",
         20280 => x"c7818283",
         20281 => x"84858687",
         20282 => x"88898a8b",
         20283 => x"8c8d8e8f",
         20284 => x"90919293",
         20285 => x"94959697",
         20286 => x"98999abc",
         20287 => x"8040a5c0",
         20288 => x"00000000",
         20289 => x"00000000",
         20290 => x"00000000",
         20291 => x"00000000",
         20292 => x"00000000",
         20293 => x"00000000",
         20294 => x"00000000",
         20295 => x"00000000",
         20296 => x"00000000",
         20297 => x"00000000",
         20298 => x"00000000",
         20299 => x"00000000",
         20300 => x"00000000",
         20301 => x"00000000",
         20302 => x"00000000",
         20303 => x"00000000",
         20304 => x"00000000",
         20305 => x"00000000",
         20306 => x"00000000",
         20307 => x"00000000",
         20308 => x"00000000",
         20309 => x"00000000",
         20310 => x"00000000",
         20311 => x"00000000",
         20312 => x"00000000",
         20313 => x"00000000",
         20314 => x"00000000",
         20315 => x"00000000",
         20316 => x"00000000",
         20317 => x"00000000",
         20318 => x"00020003",
         20319 => x"00040101",
         20320 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

