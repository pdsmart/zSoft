-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b93",
             1 => x"99040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b92",
            73 => x"fd040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b92e0",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b81e8",
           162 => x"b4738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"92e50400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80eb",
           171 => x"b62d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80ed",
           179 => x"f22d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"94040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b4040b0b",
           272 => x"0b8cc404",
           273 => x"0b0b0b8c",
           274 => x"d4040b0b",
           275 => x"0b8ce404",
           276 => x"0b0b0b8c",
           277 => x"f4040b0b",
           278 => x"0b8d8404",
           279 => x"0b0b0b8d",
           280 => x"94040b0b",
           281 => x"0b8da404",
           282 => x"0b0b0b8d",
           283 => x"b4040b0b",
           284 => x"0b8dc404",
           285 => x"0b0b0b8d",
           286 => x"d4040b0b",
           287 => x"0b8de404",
           288 => x"0b0b0b8d",
           289 => x"f4040b0b",
           290 => x"0b8e8304",
           291 => x"0b0b0b8e",
           292 => x"92040b0b",
           293 => x"0b8ea104",
           294 => x"0b0b0b8e",
           295 => x"b1040b0b",
           296 => x"0b8ec104",
           297 => x"0b0b0b8e",
           298 => x"d1040b0b",
           299 => x"0b8ee104",
           300 => x"0b0b0b8e",
           301 => x"f1040b0b",
           302 => x"0b8f8104",
           303 => x"0b0b0b8f",
           304 => x"91040b0b",
           305 => x"0b8fa104",
           306 => x"0b0b0b8f",
           307 => x"b1040b0b",
           308 => x"0b8fc104",
           309 => x"0b0b0b8f",
           310 => x"d1040b0b",
           311 => x"0b8fe104",
           312 => x"0b0b0b8f",
           313 => x"f1040b0b",
           314 => x"0b908104",
           315 => x"0b0b0b90",
           316 => x"91040b0b",
           317 => x"0b90a104",
           318 => x"0b0b0b90",
           319 => x"b1040b0b",
           320 => x"0b90c104",
           321 => x"0b0b0b90",
           322 => x"d1040b0b",
           323 => x"0b90e104",
           324 => x"0b0b0b90",
           325 => x"f1040b0b",
           326 => x"0b918104",
           327 => x"0b0b0b91",
           328 => x"91040b0b",
           329 => x"0b91a104",
           330 => x"0b0b0b91",
           331 => x"b1040b0b",
           332 => x"0b91c104",
           333 => x"0b0b0b91",
           334 => x"d1040b0b",
           335 => x"0b91e104",
           336 => x"0b0b0b91",
           337 => x"f1040b0b",
           338 => x"0b928104",
           339 => x"0b0b0b92",
           340 => x"90040b0b",
           341 => x"0b929f04",
           342 => x"0b0b0b92",
           343 => x"ae04ffff",
           344 => x"ffffffff",
           345 => x"ffffffff",
           346 => x"ffffffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"048287d8",
           386 => x"0cbe972d",
           387 => x"8287d808",
           388 => x"82a09004",
           389 => x"8287d80c",
           390 => x"80cbc32d",
           391 => x"8287d808",
           392 => x"82a09004",
           393 => x"8287d80c",
           394 => x"80cc822d",
           395 => x"8287d808",
           396 => x"82a09004",
           397 => x"8287d80c",
           398 => x"80cca02d",
           399 => x"8287d808",
           400 => x"82a09004",
           401 => x"8287d80c",
           402 => x"80d2de2d",
           403 => x"8287d808",
           404 => x"82a09004",
           405 => x"8287d80c",
           406 => x"80d3dc2d",
           407 => x"8287d808",
           408 => x"82a09004",
           409 => x"8287d80c",
           410 => x"80ccc32d",
           411 => x"8287d808",
           412 => x"82a09004",
           413 => x"8287d80c",
           414 => x"80d3f92d",
           415 => x"8287d808",
           416 => x"82a09004",
           417 => x"8287d80c",
           418 => x"80d5eb2d",
           419 => x"8287d808",
           420 => x"82a09004",
           421 => x"8287d80c",
           422 => x"80d2842d",
           423 => x"8287d808",
           424 => x"82a09004",
           425 => x"8287d80c",
           426 => x"80ccf52d",
           427 => x"8287d808",
           428 => x"82a09004",
           429 => x"8287d80c",
           430 => x"80d29a2d",
           431 => x"8287d808",
           432 => x"82a09004",
           433 => x"8287d80c",
           434 => x"80d2be2d",
           435 => x"8287d808",
           436 => x"82a09004",
           437 => x"8287d80c",
           438 => x"80c0a02d",
           439 => x"8287d808",
           440 => x"82a09004",
           441 => x"8287d80c",
           442 => x"80c0ef2d",
           443 => x"8287d808",
           444 => x"82a09004",
           445 => x"8287d80c",
           446 => x"b8d32d82",
           447 => x"87d80882",
           448 => x"a0900482",
           449 => x"87d80cba",
           450 => x"ca2d8287",
           451 => x"d80882a0",
           452 => x"90048287",
           453 => x"d80cbbfd",
           454 => x"2d8287d8",
           455 => x"0882a090",
           456 => x"048287d8",
           457 => x"0c81ab97",
           458 => x"2d8287d8",
           459 => x"0882a090",
           460 => x"048287d8",
           461 => x"0c81b888",
           462 => x"2d8287d8",
           463 => x"0882a090",
           464 => x"048287d8",
           465 => x"0c81affc",
           466 => x"2d8287d8",
           467 => x"0882a090",
           468 => x"048287d8",
           469 => x"0c81b2f9",
           470 => x"2d8287d8",
           471 => x"0882a090",
           472 => x"048287d8",
           473 => x"0c81bd97",
           474 => x"2d8287d8",
           475 => x"0882a090",
           476 => x"048287d8",
           477 => x"0c81c5f7",
           478 => x"2d8287d8",
           479 => x"0882a090",
           480 => x"048287d8",
           481 => x"0c81b6ea",
           482 => x"2d8287d8",
           483 => x"0882a090",
           484 => x"048287d8",
           485 => x"0c81c0b6",
           486 => x"2d8287d8",
           487 => x"0882a090",
           488 => x"048287d8",
           489 => x"0c81c1d5",
           490 => x"2d8287d8",
           491 => x"0882a090",
           492 => x"048287d8",
           493 => x"0c81c1f4",
           494 => x"2d8287d8",
           495 => x"0882a090",
           496 => x"048287d8",
           497 => x"0c81c9de",
           498 => x"2d8287d8",
           499 => x"0882a090",
           500 => x"048287d8",
           501 => x"0c81c7c4",
           502 => x"2d8287d8",
           503 => x"0882a090",
           504 => x"048287d8",
           505 => x"0c81ccb2",
           506 => x"2d8287d8",
           507 => x"0882a090",
           508 => x"048287d8",
           509 => x"0c81c2f8",
           510 => x"2d8287d8",
           511 => x"0882a090",
           512 => x"048287d8",
           513 => x"0c81cfb2",
           514 => x"2d8287d8",
           515 => x"0882a090",
           516 => x"048287d8",
           517 => x"0c81d0b3",
           518 => x"2d8287d8",
           519 => x"0882a090",
           520 => x"048287d8",
           521 => x"0c81b8e8",
           522 => x"2d8287d8",
           523 => x"0882a090",
           524 => x"048287d8",
           525 => x"0c81b8c1",
           526 => x"2d8287d8",
           527 => x"0882a090",
           528 => x"048287d8",
           529 => x"0c81b9ec",
           530 => x"2d8287d8",
           531 => x"0882a090",
           532 => x"048287d8",
           533 => x"0c81c3cf",
           534 => x"2d8287d8",
           535 => x"0882a090",
           536 => x"048287d8",
           537 => x"0c81d1a4",
           538 => x"2d8287d8",
           539 => x"0882a090",
           540 => x"048287d8",
           541 => x"0c81d3ae",
           542 => x"2d8287d8",
           543 => x"0882a090",
           544 => x"048287d8",
           545 => x"0c81d6f0",
           546 => x"2d8287d8",
           547 => x"0882a090",
           548 => x"048287d8",
           549 => x"0c81aab6",
           550 => x"2d8287d8",
           551 => x"0882a090",
           552 => x"048287d8",
           553 => x"0c81d9dc",
           554 => x"2d8287d8",
           555 => x"0882a090",
           556 => x"048287d8",
           557 => x"0c81e891",
           558 => x"2d8287d8",
           559 => x"0882a090",
           560 => x"048287d8",
           561 => x"0c81e5fd",
           562 => x"2d8287d8",
           563 => x"0882a090",
           564 => x"048287d8",
           565 => x"0c80fbf2",
           566 => x"2d8287d8",
           567 => x"0882a090",
           568 => x"048287d8",
           569 => x"0c80fddc",
           570 => x"2d8287d8",
           571 => x"0882a090",
           572 => x"048287d8",
           573 => x"0c80ffc0",
           574 => x"2d8287d8",
           575 => x"0882a090",
           576 => x"048287d8",
           577 => x"0cb8fc2d",
           578 => x"8287d808",
           579 => x"82a09004",
           580 => x"8287d80c",
           581 => x"baa02d82",
           582 => x"87d80882",
           583 => x"a0900482",
           584 => x"87d80cbd",
           585 => x"8d2d8287",
           586 => x"d80882a0",
           587 => x"90048287",
           588 => x"d80c9af4",
           589 => x"2d8287d8",
           590 => x"0882a090",
           591 => x"043c0400",
           592 => x"00101010",
           593 => x"10101010",
           594 => x"10101010",
           595 => x"10101010",
           596 => x"10101010",
           597 => x"10101010",
           598 => x"10101010",
           599 => x"10101010",
           600 => x"53510400",
           601 => x"007381ff",
           602 => x"06738306",
           603 => x"09810583",
           604 => x"05101010",
           605 => x"2b0772fc",
           606 => x"060c5151",
           607 => x"04727280",
           608 => x"728106ff",
           609 => x"05097206",
           610 => x"05711052",
           611 => x"720a100a",
           612 => x"5372ed38",
           613 => x"51515351",
           614 => x"048287cc",
           615 => x"70829f88",
           616 => x"278e3880",
           617 => x"71708405",
           618 => x"530c0b0b",
           619 => x"0b939c04",
           620 => x"8c8151b7",
           621 => x"ad040082",
           622 => x"87d80802",
           623 => x"8287d80c",
           624 => x"fe3d0d82",
           625 => x"87d80888",
           626 => x"05088287",
           627 => x"d808fc05",
           628 => x"0c8287d8",
           629 => x"08fc0508",
           630 => x"52713382",
           631 => x"87d808fc",
           632 => x"05088105",
           633 => x"8287d808",
           634 => x"fc050c70",
           635 => x"81ff0651",
           636 => x"5170802e",
           637 => x"8338da39",
           638 => x"8287d808",
           639 => x"fc0508ff",
           640 => x"058287d8",
           641 => x"08fc050c",
           642 => x"8287d808",
           643 => x"fc050882",
           644 => x"87d80888",
           645 => x"05083170",
           646 => x"8287cc0c",
           647 => x"51843d0d",
           648 => x"8287d80c",
           649 => x"048287d8",
           650 => x"08028287",
           651 => x"d80cfe3d",
           652 => x"0d8287d8",
           653 => x"08880508",
           654 => x"8287d808",
           655 => x"fc050c82",
           656 => x"87d8088c",
           657 => x"05085271",
           658 => x"338287d8",
           659 => x"088c0508",
           660 => x"81058287",
           661 => x"d8088c05",
           662 => x"0c8287d8",
           663 => x"08fc0508",
           664 => x"53517072",
           665 => x"348287d8",
           666 => x"08fc0508",
           667 => x"81058287",
           668 => x"d808fc05",
           669 => x"0c7081ff",
           670 => x"06517080",
           671 => x"2e8438ff",
           672 => x"be398287",
           673 => x"d8088805",
           674 => x"08708287",
           675 => x"cc0c5184",
           676 => x"3d0d8287",
           677 => x"d80c0482",
           678 => x"87d80802",
           679 => x"8287d80c",
           680 => x"fd3d0d82",
           681 => x"87d80888",
           682 => x"05088287",
           683 => x"d808fc05",
           684 => x"0c8287d8",
           685 => x"088c0508",
           686 => x"8287d808",
           687 => x"f8050c82",
           688 => x"87d80890",
           689 => x"0508802e",
           690 => x"80e53882",
           691 => x"87d80890",
           692 => x"05088105",
           693 => x"8287d808",
           694 => x"90050c82",
           695 => x"87d80890",
           696 => x"0508ff05",
           697 => x"8287d808",
           698 => x"90050c82",
           699 => x"87d80890",
           700 => x"0508802e",
           701 => x"ba388287",
           702 => x"d808f805",
           703 => x"08517033",
           704 => x"8287d808",
           705 => x"f8050881",
           706 => x"058287d8",
           707 => x"08f8050c",
           708 => x"8287d808",
           709 => x"fc050852",
           710 => x"52717134",
           711 => x"8287d808",
           712 => x"fc050881",
           713 => x"058287d8",
           714 => x"08fc050c",
           715 => x"ffad3982",
           716 => x"87d80888",
           717 => x"05087082",
           718 => x"87cc0c51",
           719 => x"853d0d82",
           720 => x"87d80c04",
           721 => x"8287d808",
           722 => x"028287d8",
           723 => x"0cfd3d0d",
           724 => x"8287d808",
           725 => x"90050880",
           726 => x"2e81f438",
           727 => x"8287d808",
           728 => x"8c050852",
           729 => x"71338287",
           730 => x"d8088c05",
           731 => x"08810582",
           732 => x"87d8088c",
           733 => x"050c8287",
           734 => x"d8088805",
           735 => x"08703372",
           736 => x"81ff0653",
           737 => x"54545171",
           738 => x"712e8438",
           739 => x"80ce3982",
           740 => x"87d80888",
           741 => x"05085271",
           742 => x"338287d8",
           743 => x"08880508",
           744 => x"81058287",
           745 => x"d8088805",
           746 => x"0c7081ff",
           747 => x"06515170",
           748 => x"8d38800b",
           749 => x"8287d808",
           750 => x"fc050c81",
           751 => x"9b398287",
           752 => x"d8089005",
           753 => x"08ff0582",
           754 => x"87d80890",
           755 => x"050c8287",
           756 => x"d8089005",
           757 => x"08802e84",
           758 => x"38ff8139",
           759 => x"8287d808",
           760 => x"90050880",
           761 => x"2e80e838",
           762 => x"8287d808",
           763 => x"88050870",
           764 => x"33525370",
           765 => x"8d38ff0b",
           766 => x"8287d808",
           767 => x"fc050c80",
           768 => x"d7398287",
           769 => x"d8088c05",
           770 => x"08ff0582",
           771 => x"87d8088c",
           772 => x"050c8287",
           773 => x"d8088c05",
           774 => x"08703352",
           775 => x"52708c38",
           776 => x"810b8287",
           777 => x"d808fc05",
           778 => x"0cae3982",
           779 => x"87d80888",
           780 => x"05087033",
           781 => x"8287d808",
           782 => x"8c050870",
           783 => x"33727131",
           784 => x"708287d8",
           785 => x"08fc050c",
           786 => x"53555252",
           787 => x"538a3980",
           788 => x"0b8287d8",
           789 => x"08fc050c",
           790 => x"8287d808",
           791 => x"fc050882",
           792 => x"87cc0c85",
           793 => x"3d0d8287",
           794 => x"d80c0482",
           795 => x"87d80802",
           796 => x"8287d80c",
           797 => x"fe3d0d82",
           798 => x"87d80888",
           799 => x"05088287",
           800 => x"d808fc05",
           801 => x"0c8287d8",
           802 => x"08900508",
           803 => x"802e80d4",
           804 => x"388287d8",
           805 => x"08900508",
           806 => x"81058287",
           807 => x"d8089005",
           808 => x"0c8287d8",
           809 => x"08900508",
           810 => x"ff058287",
           811 => x"d8089005",
           812 => x"0c8287d8",
           813 => x"08900508",
           814 => x"802ea938",
           815 => x"8287d808",
           816 => x"8c050851",
           817 => x"708287d8",
           818 => x"08fc0508",
           819 => x"52527171",
           820 => x"348287d8",
           821 => x"08fc0508",
           822 => x"81058287",
           823 => x"d808fc05",
           824 => x"0cffbe39",
           825 => x"8287d808",
           826 => x"88050870",
           827 => x"8287cc0c",
           828 => x"51843d0d",
           829 => x"8287d80c",
           830 => x"04f93d0d",
           831 => x"79700870",
           832 => x"56565874",
           833 => x"802e80e3",
           834 => x"38953975",
           835 => x"0851f9a7",
           836 => x"3f8287cc",
           837 => x"0815780c",
           838 => x"85163354",
           839 => x"80cd3974",
           840 => x"335473a0",
           841 => x"2e098106",
           842 => x"86388115",
           843 => x"55f13980",
           844 => x"57769029",
           845 => x"8282cc05",
           846 => x"70085256",
           847 => x"f8f93f82",
           848 => x"87cc0853",
           849 => x"74527508",
           850 => x"51fbf93f",
           851 => x"8287cc08",
           852 => x"8b388416",
           853 => x"33547381",
           854 => x"2effb038",
           855 => x"81177081",
           856 => x"ff065854",
           857 => x"997727c9",
           858 => x"38ff5473",
           859 => x"8287cc0c",
           860 => x"893d0d04",
           861 => x"ff3d0d73",
           862 => x"52719326",
           863 => x"818e3871",
           864 => x"842981e8",
           865 => x"c4055271",
           866 => x"080481eb",
           867 => x"ac518180",
           868 => x"3981ebb8",
           869 => x"5180f939",
           870 => x"81ebcc51",
           871 => x"80f23981",
           872 => x"ebe05180",
           873 => x"eb3981eb",
           874 => x"f05180e4",
           875 => x"3981ec80",
           876 => x"5180dd39",
           877 => x"81ec9451",
           878 => x"80d63981",
           879 => x"eca45180",
           880 => x"cf3981ec",
           881 => x"bc5180c8",
           882 => x"3981ecd4",
           883 => x"5180c139",
           884 => x"81ecec51",
           885 => x"bb3981ed",
           886 => x"8851b539",
           887 => x"81ed9c51",
           888 => x"af3981ed",
           889 => x"c851a939",
           890 => x"81eddc51",
           891 => x"a33981ed",
           892 => x"fc519d39",
           893 => x"81ee9051",
           894 => x"973981ee",
           895 => x"a8519139",
           896 => x"81eec051",
           897 => x"8b3981ee",
           898 => x"d8518539",
           899 => x"81eee451",
           900 => x"b08e3f83",
           901 => x"3d0d04fb",
           902 => x"3d0d7779",
           903 => x"56567487",
           904 => x"e7268a38",
           905 => x"74527587",
           906 => x"e8295191",
           907 => x"3987e852",
           908 => x"745180cf",
           909 => x"b63f8287",
           910 => x"cc085275",
           911 => x"5180cfab",
           912 => x"3f8287cc",
           913 => x"08547953",
           914 => x"755281ee",
           915 => x"f451b5b4",
           916 => x"3f873d0d",
           917 => x"04ec3d0d",
           918 => x"66028405",
           919 => x"80e30533",
           920 => x"5b578068",
           921 => x"7830707a",
           922 => x"07732551",
           923 => x"57595978",
           924 => x"567787ff",
           925 => x"26833881",
           926 => x"56747607",
           927 => x"7081ff06",
           928 => x"51559356",
           929 => x"74818238",
           930 => x"81537652",
           931 => x"8c3d7052",
           932 => x"56818e83",
           933 => x"3f8287cc",
           934 => x"08578287",
           935 => x"cc08b938",
           936 => x"8287cc08",
           937 => x"87c09888",
           938 => x"0c8287cc",
           939 => x"0859963d",
           940 => x"d4055484",
           941 => x"80537752",
           942 => x"75518192",
           943 => x"bf3f8287",
           944 => x"cc085782",
           945 => x"87cc0890",
           946 => x"387a5574",
           947 => x"802e8938",
           948 => x"74197519",
           949 => x"5959d739",
           950 => x"963dd805",
           951 => x"51819aa8",
           952 => x"3f763070",
           953 => x"78078025",
           954 => x"7b30709f",
           955 => x"2a720651",
           956 => x"57515674",
           957 => x"802e9038",
           958 => x"81ef9853",
           959 => x"87c09888",
           960 => x"08527851",
           961 => x"fe913f76",
           962 => x"56758287",
           963 => x"cc0c963d",
           964 => x"0d04f93d",
           965 => x"0d7b0284",
           966 => x"05b30533",
           967 => x"5758ff57",
           968 => x"80537a52",
           969 => x"7951fead",
           970 => x"3f8287cc",
           971 => x"08a43875",
           972 => x"802e8838",
           973 => x"75812e98",
           974 => x"38983960",
           975 => x"557f5482",
           976 => x"87cc537e",
           977 => x"527d5177",
           978 => x"2d8287cc",
           979 => x"08578339",
           980 => x"77047682",
           981 => x"87cc0c89",
           982 => x"3d0d04f3",
           983 => x"3d0d7f61",
           984 => x"63028c05",
           985 => x"80cf0533",
           986 => x"73731568",
           987 => x"415f5c5c",
           988 => x"5e5e5e7a",
           989 => x"5281efa0",
           990 => x"51b3893f",
           991 => x"81efa851",
           992 => x"ad9e3f80",
           993 => x"55747927",
           994 => x"80f4387b",
           995 => x"902e8938",
           996 => x"7ba02ea4",
           997 => x"3880c139",
           998 => x"74185372",
           999 => x"7a278d38",
          1000 => x"72225281",
          1001 => x"efac51b2",
          1002 => x"db3f8839",
          1003 => x"81efb851",
          1004 => x"acee3f82",
          1005 => x"1555bf39",
          1006 => x"74185372",
          1007 => x"7a278d38",
          1008 => x"72085281",
          1009 => x"efa051b2",
          1010 => x"bb3f8839",
          1011 => x"81efb451",
          1012 => x"acce3f84",
          1013 => x"15559f39",
          1014 => x"74185372",
          1015 => x"7a278d38",
          1016 => x"72335281",
          1017 => x"efc051b2",
          1018 => x"9b3f8839",
          1019 => x"81efc851",
          1020 => x"acae3f81",
          1021 => x"1555a051",
          1022 => x"abc93fff",
          1023 => x"883981ef",
          1024 => x"cc51ac9c",
          1025 => x"3f805574",
          1026 => x"7927bb38",
          1027 => x"74187033",
          1028 => x"55538056",
          1029 => x"727a2783",
          1030 => x"38815680",
          1031 => x"539f7427",
          1032 => x"83388153",
          1033 => x"75730670",
          1034 => x"81ff0651",
          1035 => x"5372802e",
          1036 => x"8b387380",
          1037 => x"fe268538",
          1038 => x"73518339",
          1039 => x"a051ab83",
          1040 => x"3f811555",
          1041 => x"c23981ef",
          1042 => x"d051abd4",
          1043 => x"3f781879",
          1044 => x"1c5c58a0",
          1045 => x"9a3f8287",
          1046 => x"cc08982b",
          1047 => x"70982c51",
          1048 => x"5776a02e",
          1049 => x"098106aa",
          1050 => x"38a0843f",
          1051 => x"8287cc08",
          1052 => x"982b7098",
          1053 => x"2c70a032",
          1054 => x"7030729b",
          1055 => x"32703070",
          1056 => x"72077375",
          1057 => x"07065158",
          1058 => x"58595751",
          1059 => x"57807324",
          1060 => x"d838769b",
          1061 => x"2e098106",
          1062 => x"85388053",
          1063 => x"8c397c1e",
          1064 => x"53727826",
          1065 => x"fdcd38ff",
          1066 => x"53728287",
          1067 => x"cc0c8f3d",
          1068 => x"0d04fc3d",
          1069 => x"0d029b05",
          1070 => x"3381efd4",
          1071 => x"5381efdc",
          1072 => x"5255b0c0",
          1073 => x"3f8286a4",
          1074 => x"2251a8dc",
          1075 => x"3f81efe8",
          1076 => x"5481eff4",
          1077 => x"538286a5",
          1078 => x"335281ef",
          1079 => x"fc51b0a4",
          1080 => x"3f74802e",
          1081 => x"8438a4a9",
          1082 => x"3f863d0d",
          1083 => x"04fe3d0d",
          1084 => x"87c09680",
          1085 => x"0853a9b9",
          1086 => x"3f81519b",
          1087 => x"903f81f0",
          1088 => x"98519d83",
          1089 => x"3f80519b",
          1090 => x"843f7281",
          1091 => x"2a708106",
          1092 => x"51527180",
          1093 => x"2e923881",
          1094 => x"519af23f",
          1095 => x"81f0b451",
          1096 => x"9ce53f80",
          1097 => x"519ae63f",
          1098 => x"72822a70",
          1099 => x"81065152",
          1100 => x"71802e92",
          1101 => x"3881519a",
          1102 => x"d43f81f0",
          1103 => x"c8519cc7",
          1104 => x"3f80519a",
          1105 => x"c83f7283",
          1106 => x"2a708106",
          1107 => x"51527180",
          1108 => x"2e923881",
          1109 => x"519ab63f",
          1110 => x"81f0d851",
          1111 => x"9ca93f80",
          1112 => x"519aaa3f",
          1113 => x"72842a70",
          1114 => x"81065152",
          1115 => x"71802e92",
          1116 => x"3881519a",
          1117 => x"983f81f0",
          1118 => x"ec519c8b",
          1119 => x"3f80519a",
          1120 => x"8c3f7285",
          1121 => x"2a708106",
          1122 => x"51527180",
          1123 => x"2e923881",
          1124 => x"5199fa3f",
          1125 => x"81f18051",
          1126 => x"9bed3f80",
          1127 => x"5199ee3f",
          1128 => x"72862a70",
          1129 => x"81065152",
          1130 => x"71802e92",
          1131 => x"38815199",
          1132 => x"dc3f81f1",
          1133 => x"94519bcf",
          1134 => x"3f805199",
          1135 => x"d03f7287",
          1136 => x"2a708106",
          1137 => x"51527180",
          1138 => x"2e923881",
          1139 => x"5199be3f",
          1140 => x"81f1a851",
          1141 => x"9bb13f80",
          1142 => x"5199b23f",
          1143 => x"72882a70",
          1144 => x"81065152",
          1145 => x"71802e92",
          1146 => x"38815199",
          1147 => x"a03f81f1",
          1148 => x"bc519b93",
          1149 => x"3f805199",
          1150 => x"943fa7bd",
          1151 => x"3f843d0d",
          1152 => x"04fb3d0d",
          1153 => x"77028405",
          1154 => x"a3053370",
          1155 => x"55565680",
          1156 => x"527551f4",
          1157 => x"d63f0b0b",
          1158 => x"8282c833",
          1159 => x"5473a938",
          1160 => x"815381f1",
          1161 => x"fc52829e",
          1162 => x"ac518186",
          1163 => x"ea3f8287",
          1164 => x"cc083070",
          1165 => x"8287cc08",
          1166 => x"07802582",
          1167 => x"71315151",
          1168 => x"54730b0b",
          1169 => x"8282c834",
          1170 => x"0b0b8282",
          1171 => x"c8335473",
          1172 => x"812e0981",
          1173 => x"06af3882",
          1174 => x"9eac5374",
          1175 => x"52755181",
          1176 => x"c19b3f82",
          1177 => x"87cc0880",
          1178 => x"2e8b3882",
          1179 => x"87cc0851",
          1180 => x"a7ae3f91",
          1181 => x"39829eac",
          1182 => x"5181938c",
          1183 => x"3f820b0b",
          1184 => x"0b8282c8",
          1185 => x"340b0b82",
          1186 => x"82c83354",
          1187 => x"73822e09",
          1188 => x"81068c38",
          1189 => x"81f28c53",
          1190 => x"74527551",
          1191 => x"b9ba3f80",
          1192 => x"0b8287cc",
          1193 => x"0c873d0d",
          1194 => x"04ce3d0d",
          1195 => x"80707182",
          1196 => x"9ea80c5f",
          1197 => x"5d81527c",
          1198 => x"5180d5b7",
          1199 => x"3f8287cc",
          1200 => x"0881ff06",
          1201 => x"59787d2e",
          1202 => x"098106a1",
          1203 => x"3881f298",
          1204 => x"52963d70",
          1205 => x"5259acc2",
          1206 => x"3f7c5378",
          1207 => x"528288d8",
          1208 => x"518184d2",
          1209 => x"3f8287cc",
          1210 => x"087d2e88",
          1211 => x"3881f29c",
          1212 => x"5191b439",
          1213 => x"81705f5d",
          1214 => x"81f2d451",
          1215 => x"a6a23f96",
          1216 => x"3d70465a",
          1217 => x"80f85279",
          1218 => x"51fdf63f",
          1219 => x"b43dff84",
          1220 => x"0551f3e5",
          1221 => x"3f8287cc",
          1222 => x"08902b70",
          1223 => x"902c5159",
          1224 => x"7880c12e",
          1225 => x"89d13878",
          1226 => x"80c12480",
          1227 => x"d93878ab",
          1228 => x"2e83b838",
          1229 => x"78ab24a4",
          1230 => x"3878822e",
          1231 => x"81b33878",
          1232 => x"82248a38",
          1233 => x"78802eff",
          1234 => x"af388ee1",
          1235 => x"3978842e",
          1236 => x"82833878",
          1237 => x"942e82ad",
          1238 => x"388ed239",
          1239 => x"78bd2e84",
          1240 => x"fa3878bd",
          1241 => x"24903878",
          1242 => x"b02e83a5",
          1243 => x"3878bc2e",
          1244 => x"8483388e",
          1245 => x"b83978bf",
          1246 => x"2e85c138",
          1247 => x"7880c02e",
          1248 => x"86b7388e",
          1249 => x"a8397880",
          1250 => x"d52e8d88",
          1251 => x"387880d5",
          1252 => x"24b03878",
          1253 => x"80d02e8c",
          1254 => x"c1387880",
          1255 => x"d0249238",
          1256 => x"7880c22e",
          1257 => x"89f23878",
          1258 => x"80c32e8b",
          1259 => x"94388dfd",
          1260 => x"397880d1",
          1261 => x"2e8cb238",
          1262 => x"7880d42e",
          1263 => x"8cba388d",
          1264 => x"ec397881",
          1265 => x"822e8dc6",
          1266 => x"38788182",
          1267 => x"24923878",
          1268 => x"80f82e8c",
          1269 => x"db387880",
          1270 => x"f92e8cf7",
          1271 => x"388dce39",
          1272 => x"7881832e",
          1273 => x"8db53878",
          1274 => x"81852e8d",
          1275 => x"ba388dbd",
          1276 => x"39b43dff",
          1277 => x"801153ff",
          1278 => x"840551ab",
          1279 => x"fc3f8287",
          1280 => x"cc088838",
          1281 => x"81f2d851",
          1282 => x"8f9d39b4",
          1283 => x"3dfefc11",
          1284 => x"53ff8405",
          1285 => x"51abe23f",
          1286 => x"8287cc08",
          1287 => x"802e8838",
          1288 => x"81632583",
          1289 => x"38804302",
          1290 => x"80cb0533",
          1291 => x"520280cf",
          1292 => x"05335180",
          1293 => x"d2bd3f82",
          1294 => x"87cc0881",
          1295 => x"ff065978",
          1296 => x"8d3881f2",
          1297 => x"e851a3d8",
          1298 => x"3f815efd",
          1299 => x"ab3981f2",
          1300 => x"f851879d",
          1301 => x"39b43dff",
          1302 => x"801153ff",
          1303 => x"840551ab",
          1304 => x"983f8287",
          1305 => x"cc08802e",
          1306 => x"fd8e3880",
          1307 => x"53805202",
          1308 => x"80cf0533",
          1309 => x"5180d6c8",
          1310 => x"3f8287cc",
          1311 => x"085281f3",
          1312 => x"90518c84",
          1313 => x"39b43dff",
          1314 => x"801153ff",
          1315 => x"840551aa",
          1316 => x"e83f8287",
          1317 => x"cc08802e",
          1318 => x"87386389",
          1319 => x"26fcd938",
          1320 => x"b43dfefc",
          1321 => x"1153ff84",
          1322 => x"0551aacd",
          1323 => x"3f8287cc",
          1324 => x"08863882",
          1325 => x"87cc0843",
          1326 => x"635381f3",
          1327 => x"98527951",
          1328 => x"a8d83f02",
          1329 => x"80cb0533",
          1330 => x"53795263",
          1331 => x"84b42982",
          1332 => x"88d80551",
          1333 => x"8180df3f",
          1334 => x"8287cc08",
          1335 => x"818c3881",
          1336 => x"f2e851a2",
          1337 => x"bb3f815d",
          1338 => x"fc8e39b4",
          1339 => x"3dff8405",
          1340 => x"518f893f",
          1341 => x"8287cc08",
          1342 => x"b53dff84",
          1343 => x"05525b90",
          1344 => x"9f3f8153",
          1345 => x"8287cc08",
          1346 => x"527a51f2",
          1347 => x"c83f80d1",
          1348 => x"39b43dff",
          1349 => x"8405518e",
          1350 => x"e33f8287",
          1351 => x"cc08b53d",
          1352 => x"ff840552",
          1353 => x"5b8ff93f",
          1354 => x"8287cc08",
          1355 => x"b53dff84",
          1356 => x"05525a8f",
          1357 => x"eb3f8287",
          1358 => x"cc08b53d",
          1359 => x"ff840552",
          1360 => x"598fdd3f",
          1361 => x"8285f058",
          1362 => x"8287dc57",
          1363 => x"80568055",
          1364 => x"8287cc08",
          1365 => x"81ff0654",
          1366 => x"78537952",
          1367 => x"7a51f3b2",
          1368 => x"3f8287cc",
          1369 => x"08802efb",
          1370 => x"8f388287",
          1371 => x"cc0851f0",
          1372 => x"833ffb84",
          1373 => x"39b43dff",
          1374 => x"801153ff",
          1375 => x"840551a8",
          1376 => x"f83f8287",
          1377 => x"cc08802e",
          1378 => x"faee38b4",
          1379 => x"3dfefc11",
          1380 => x"53ff8405",
          1381 => x"51a8e23f",
          1382 => x"8287cc08",
          1383 => x"802efad8",
          1384 => x"38b43dfe",
          1385 => x"f81153ff",
          1386 => x"840551a8",
          1387 => x"cc3f8287",
          1388 => x"cc088638",
          1389 => x"8287cc08",
          1390 => x"4281f39c",
          1391 => x"51a0e13f",
          1392 => x"63635c5a",
          1393 => x"797b2781",
          1394 => x"e9386159",
          1395 => x"787a7084",
          1396 => x"055c0c7a",
          1397 => x"7a26f538",
          1398 => x"81d839b4",
          1399 => x"3dff8011",
          1400 => x"53ff8405",
          1401 => x"51a8923f",
          1402 => x"8287cc08",
          1403 => x"802efa88",
          1404 => x"38b43dfe",
          1405 => x"fc1153ff",
          1406 => x"840551a7",
          1407 => x"fc3f8287",
          1408 => x"cc08802e",
          1409 => x"f9f238b4",
          1410 => x"3dfef811",
          1411 => x"53ff8405",
          1412 => x"51a7e63f",
          1413 => x"8287cc08",
          1414 => x"802ef9dc",
          1415 => x"3881f3ac",
          1416 => x"519ffd3f",
          1417 => x"635a7963",
          1418 => x"27818738",
          1419 => x"61597970",
          1420 => x"81055b33",
          1421 => x"79346181",
          1422 => x"0542eb39",
          1423 => x"b43dff80",
          1424 => x"1153ff84",
          1425 => x"0551a7b1",
          1426 => x"3f8287cc",
          1427 => x"08802ef9",
          1428 => x"a738b43d",
          1429 => x"fefc1153",
          1430 => x"ff840551",
          1431 => x"a79b3f82",
          1432 => x"87cc0880",
          1433 => x"2ef99138",
          1434 => x"b43dfef8",
          1435 => x"1153ff84",
          1436 => x"0551a785",
          1437 => x"3f8287cc",
          1438 => x"08802ef8",
          1439 => x"fb3881f3",
          1440 => x"b8519f9c",
          1441 => x"3f635a79",
          1442 => x"6327a738",
          1443 => x"6170337b",
          1444 => x"335e5a5b",
          1445 => x"787c2e91",
          1446 => x"3878557a",
          1447 => x"54793353",
          1448 => x"795281f3",
          1449 => x"c851a4dc",
          1450 => x"3f811a62",
          1451 => x"8105435a",
          1452 => x"d63981f2",
          1453 => x"e45182b9",
          1454 => x"39b43dff",
          1455 => x"801153ff",
          1456 => x"840551a6",
          1457 => x"b43f8287",
          1458 => x"cc0880df",
          1459 => x"388286b8",
          1460 => x"33597880",
          1461 => x"2e893882",
          1462 => x"85f00844",
          1463 => x"80cd3982",
          1464 => x"86b93359",
          1465 => x"78802e88",
          1466 => x"388285f8",
          1467 => x"0844bc39",
          1468 => x"8286ba33",
          1469 => x"5978802e",
          1470 => x"88388286",
          1471 => x"800844ab",
          1472 => x"398286bb",
          1473 => x"33597880",
          1474 => x"2e883882",
          1475 => x"86880844",
          1476 => x"9a398286",
          1477 => x"b6335978",
          1478 => x"802e8838",
          1479 => x"82869008",
          1480 => x"44893982",
          1481 => x"86a008fc",
          1482 => x"800544b4",
          1483 => x"3dfefc11",
          1484 => x"53ff8405",
          1485 => x"51a5c23f",
          1486 => x"8287cc08",
          1487 => x"80de3882",
          1488 => x"86b83359",
          1489 => x"78802e89",
          1490 => x"388285f4",
          1491 => x"084380cc",
          1492 => x"398286b9",
          1493 => x"33597880",
          1494 => x"2e883882",
          1495 => x"85fc0843",
          1496 => x"bb398286",
          1497 => x"ba335978",
          1498 => x"802e8838",
          1499 => x"82868408",
          1500 => x"43aa3982",
          1501 => x"86bb3359",
          1502 => x"78802e88",
          1503 => x"3882868c",
          1504 => x"08439939",
          1505 => x"8286b633",
          1506 => x"5978802e",
          1507 => x"88388286",
          1508 => x"94084388",
          1509 => x"398286a0",
          1510 => x"08880543",
          1511 => x"b43dfef8",
          1512 => x"1153ff84",
          1513 => x"0551a4d1",
          1514 => x"3f8287cc",
          1515 => x"08802ea7",
          1516 => x"3880625c",
          1517 => x"5c7a882e",
          1518 => x"8338815c",
          1519 => x"7a903270",
          1520 => x"30707207",
          1521 => x"9f2a707f",
          1522 => x"0651515a",
          1523 => x"5a78802e",
          1524 => x"88387aa0",
          1525 => x"2e833888",
          1526 => x"4281f3e4",
          1527 => x"519cc13f",
          1528 => x"a0556354",
          1529 => x"61536252",
          1530 => x"6351eeef",
          1531 => x"3f81f3f4",
          1532 => x"519cad3f",
          1533 => x"f68239b4",
          1534 => x"3dff8011",
          1535 => x"53ff8405",
          1536 => x"51a3f63f",
          1537 => x"8287cc08",
          1538 => x"802ef5ec",
          1539 => x"38b43dfe",
          1540 => x"fc1153ff",
          1541 => x"840551a3",
          1542 => x"e03f8287",
          1543 => x"cc08802e",
          1544 => x"a4386359",
          1545 => x"0280cb05",
          1546 => x"33793463",
          1547 => x"810544b4",
          1548 => x"3dfefc11",
          1549 => x"53ff8405",
          1550 => x"51a3be3f",
          1551 => x"8287cc08",
          1552 => x"e138f5b4",
          1553 => x"39637033",
          1554 => x"545281f4",
          1555 => x"8051a1b4",
          1556 => x"3f80f852",
          1557 => x"7951a286",
          1558 => x"3f794579",
          1559 => x"335978ae",
          1560 => x"2ef59538",
          1561 => x"9f79279f",
          1562 => x"38b43dfe",
          1563 => x"fc1153ff",
          1564 => x"840551a3",
          1565 => x"843f8287",
          1566 => x"cc08802e",
          1567 => x"91386359",
          1568 => x"0280cb05",
          1569 => x"33793463",
          1570 => x"810544ff",
          1571 => x"b83981f4",
          1572 => x"8c519b8c",
          1573 => x"3fffae39",
          1574 => x"b43dfef4",
          1575 => x"1153ff84",
          1576 => x"0551a4c7",
          1577 => x"3f8287cc",
          1578 => x"08802ef4",
          1579 => x"cb38b43d",
          1580 => x"fef01153",
          1581 => x"ff840551",
          1582 => x"a4b13f82",
          1583 => x"87cc0880",
          1584 => x"2ea53860",
          1585 => x"5902be05",
          1586 => x"22797082",
          1587 => x"055b2378",
          1588 => x"41b43dfe",
          1589 => x"f01153ff",
          1590 => x"840551a4",
          1591 => x"8e3f8287",
          1592 => x"cc08e038",
          1593 => x"f4923960",
          1594 => x"70225452",
          1595 => x"81f49451",
          1596 => x"a0923f80",
          1597 => x"f8527951",
          1598 => x"a0e43f79",
          1599 => x"45793359",
          1600 => x"78ae2ef3",
          1601 => x"f338789f",
          1602 => x"26873860",
          1603 => x"820541d7",
          1604 => x"39b43dfe",
          1605 => x"f01153ff",
          1606 => x"840551a3",
          1607 => x"ce3f8287",
          1608 => x"cc08802e",
          1609 => x"92386059",
          1610 => x"02be0522",
          1611 => x"79708205",
          1612 => x"5b237841",
          1613 => x"ffb13981",
          1614 => x"f48c5199",
          1615 => x"e33fffa7",
          1616 => x"39b43dfe",
          1617 => x"f41153ff",
          1618 => x"840551a3",
          1619 => x"9e3f8287",
          1620 => x"cc08802e",
          1621 => x"f3a238b4",
          1622 => x"3dfef011",
          1623 => x"53ff8405",
          1624 => x"51a3883f",
          1625 => x"8287cc08",
          1626 => x"802ea038",
          1627 => x"6060710c",
          1628 => x"59608405",
          1629 => x"41b43dfe",
          1630 => x"f01153ff",
          1631 => x"840551a2",
          1632 => x"ea3f8287",
          1633 => x"cc08e538",
          1634 => x"f2ee3960",
          1635 => x"70085452",
          1636 => x"81f4a051",
          1637 => x"9eee3f80",
          1638 => x"f8527951",
          1639 => x"9fc03f79",
          1640 => x"45793359",
          1641 => x"78ae2ef2",
          1642 => x"cf389f79",
          1643 => x"279b38b4",
          1644 => x"3dfef011",
          1645 => x"53ff8405",
          1646 => x"51a2b03f",
          1647 => x"8287cc08",
          1648 => x"802e8d38",
          1649 => x"6060710c",
          1650 => x"59608405",
          1651 => x"41ffbc39",
          1652 => x"81f48c51",
          1653 => x"98ca3fff",
          1654 => x"b23981f4",
          1655 => x"ac5198c0",
          1656 => x"3f825197",
          1657 => x"a73ff290",
          1658 => x"3981f4c4",
          1659 => x"5198b13f",
          1660 => x"a25196fc",
          1661 => x"3ff28139",
          1662 => x"81f4dc51",
          1663 => x"98a23f84",
          1664 => x"80810b87",
          1665 => x"c094840c",
          1666 => x"8480810b",
          1667 => x"87c09494",
          1668 => x"0cf1e539",
          1669 => x"81f4f051",
          1670 => x"98863f8c",
          1671 => x"80830b87",
          1672 => x"c094840c",
          1673 => x"8c80830b",
          1674 => x"87c09494",
          1675 => x"0cf1c939",
          1676 => x"b43dff80",
          1677 => x"1153ff84",
          1678 => x"05519fbd",
          1679 => x"3f8287cc",
          1680 => x"08802ef1",
          1681 => x"b3386352",
          1682 => x"81f58451",
          1683 => x"9db63f63",
          1684 => x"597804b4",
          1685 => x"3dff8011",
          1686 => x"53ff8405",
          1687 => x"519f9a3f",
          1688 => x"8287cc08",
          1689 => x"802ef190",
          1690 => x"38635281",
          1691 => x"f5a0519d",
          1692 => x"933f6359",
          1693 => x"782d8287",
          1694 => x"cc08802e",
          1695 => x"f0fa3882",
          1696 => x"87cc0852",
          1697 => x"81f5bc51",
          1698 => x"9cfa3ff0",
          1699 => x"eb3981f5",
          1700 => x"d851978c",
          1701 => x"3fde823f",
          1702 => x"f0de3981",
          1703 => x"f5f45196",
          1704 => x"ff3f8059",
          1705 => x"ffab3990",
          1706 => x"e83ff0cc",
          1707 => x"39794579",
          1708 => x"33597880",
          1709 => x"2ef0c138",
          1710 => x"7d7d0659",
          1711 => x"78802e81",
          1712 => x"ce38b43d",
          1713 => x"ff840551",
          1714 => x"83b23f82",
          1715 => x"87cc085b",
          1716 => x"815c7b82",
          1717 => x"2eb1387b",
          1718 => x"82248938",
          1719 => x"7b812e8c",
          1720 => x"3880ca39",
          1721 => x"7b832eae",
          1722 => x"3880c239",
          1723 => x"81f68856",
          1724 => x"7a5581f6",
          1725 => x"8c548053",
          1726 => x"81f69052",
          1727 => x"b43dffb0",
          1728 => x"05519c96",
          1729 => x"3fb83981",
          1730 => x"f6b052b4",
          1731 => x"3dffb005",
          1732 => x"519c873f",
          1733 => x"a9397a55",
          1734 => x"81f68c54",
          1735 => x"805381f6",
          1736 => x"a052b43d",
          1737 => x"ffb00551",
          1738 => x"9bf03f92",
          1739 => x"397a5480",
          1740 => x"5381f6ac",
          1741 => x"52b43dff",
          1742 => x"b005519b",
          1743 => x"dd3f8285",
          1744 => x"f0588287",
          1745 => x"dc578056",
          1746 => x"64558054",
          1747 => x"82a08053",
          1748 => x"82a08052",
          1749 => x"b43dffb0",
          1750 => x"0551e7b6",
          1751 => x"3f8287cc",
          1752 => x"088287cc",
          1753 => x"08097030",
          1754 => x"70720780",
          1755 => x"25515b5b",
          1756 => x"5f805a7b",
          1757 => x"83268338",
          1758 => x"815a787a",
          1759 => x"06597880",
          1760 => x"2e8d3881",
          1761 => x"1c7081ff",
          1762 => x"065d597b",
          1763 => x"fec4387d",
          1764 => x"81327d81",
          1765 => x"32075978",
          1766 => x"8a387eff",
          1767 => x"2e098106",
          1768 => x"eed63881",
          1769 => x"f6b4519a",
          1770 => x"db3feecc",
          1771 => x"39fc3d0d",
          1772 => x"800b8287",
          1773 => x"dc3487c0",
          1774 => x"948c7008",
          1775 => x"54558784",
          1776 => x"80527251",
          1777 => x"b4a53f82",
          1778 => x"87cc0890",
          1779 => x"2b750855",
          1780 => x"53878480",
          1781 => x"527351b4",
          1782 => x"923f7282",
          1783 => x"87cc0807",
          1784 => x"750c87c0",
          1785 => x"949c7008",
          1786 => x"54558784",
          1787 => x"80527251",
          1788 => x"b3f93f82",
          1789 => x"87cc0890",
          1790 => x"2b750855",
          1791 => x"53878480",
          1792 => x"527351b3",
          1793 => x"e63f7282",
          1794 => x"87cc0807",
          1795 => x"750c8c80",
          1796 => x"830b87c0",
          1797 => x"94840c8c",
          1798 => x"80830b87",
          1799 => x"c094940c",
          1800 => x"bda50b82",
          1801 => x"9ed40c80",
          1802 => x"c0a00b82",
          1803 => x"9ed80c89",
          1804 => x"943f92fd",
          1805 => x"3f81f6c4",
          1806 => x"5193e53f",
          1807 => x"81f6d051",
          1808 => x"93de3fa1",
          1809 => x"ed5192a3",
          1810 => x"3f8151e8",
          1811 => x"e53fecd9",
          1812 => x"3f8004fe",
          1813 => x"3d0d8052",
          1814 => x"83537188",
          1815 => x"2b5287c0",
          1816 => x"3f8287cc",
          1817 => x"0881ff06",
          1818 => x"7207ff14",
          1819 => x"54527280",
          1820 => x"25e83871",
          1821 => x"8287cc0c",
          1822 => x"843d0d04",
          1823 => x"fc3d0d76",
          1824 => x"70085455",
          1825 => x"80735254",
          1826 => x"72742e81",
          1827 => x"8a387233",
          1828 => x"5170a02e",
          1829 => x"09810686",
          1830 => x"38811353",
          1831 => x"f1397233",
          1832 => x"5170a22e",
          1833 => x"09810686",
          1834 => x"38811353",
          1835 => x"81547252",
          1836 => x"73812e09",
          1837 => x"81069f38",
          1838 => x"84398112",
          1839 => x"52807233",
          1840 => x"525470a2",
          1841 => x"2e833881",
          1842 => x"5470802e",
          1843 => x"9d3873ea",
          1844 => x"38983981",
          1845 => x"12528072",
          1846 => x"33525470",
          1847 => x"a02e8338",
          1848 => x"81547080",
          1849 => x"2e843873",
          1850 => x"ea388072",
          1851 => x"33525470",
          1852 => x"a02e0981",
          1853 => x"06833881",
          1854 => x"5470a232",
          1855 => x"70307080",
          1856 => x"25760751",
          1857 => x"51517080",
          1858 => x"2e883880",
          1859 => x"72708105",
          1860 => x"54347175",
          1861 => x"0c725170",
          1862 => x"8287cc0c",
          1863 => x"863d0d04",
          1864 => x"fc3d0d76",
          1865 => x"53720880",
          1866 => x"2e913886",
          1867 => x"3dfc0552",
          1868 => x"72519bb7",
          1869 => x"3f8287cc",
          1870 => x"08853880",
          1871 => x"53833974",
          1872 => x"53728287",
          1873 => x"cc0c863d",
          1874 => x"0d04fc3d",
          1875 => x"0d768211",
          1876 => x"33ff0552",
          1877 => x"53815270",
          1878 => x"8b268198",
          1879 => x"38831333",
          1880 => x"ff055182",
          1881 => x"52709e26",
          1882 => x"818a3884",
          1883 => x"13335183",
          1884 => x"52709726",
          1885 => x"80fe3885",
          1886 => x"13335184",
          1887 => x"5270bb26",
          1888 => x"80f23886",
          1889 => x"13335185",
          1890 => x"5270bb26",
          1891 => x"80e63888",
          1892 => x"13225586",
          1893 => x"527487e7",
          1894 => x"2680d938",
          1895 => x"8a132254",
          1896 => x"87527387",
          1897 => x"e72680cc",
          1898 => x"38810b87",
          1899 => x"c0989c0c",
          1900 => x"722287c0",
          1901 => x"98bc0c82",
          1902 => x"133387c0",
          1903 => x"98b80c83",
          1904 => x"133387c0",
          1905 => x"98b40c84",
          1906 => x"133387c0",
          1907 => x"98b00c85",
          1908 => x"133387c0",
          1909 => x"98ac0c86",
          1910 => x"133387c0",
          1911 => x"98a80c74",
          1912 => x"87c098a4",
          1913 => x"0c7387c0",
          1914 => x"98a00c80",
          1915 => x"0b87c098",
          1916 => x"9c0c8052",
          1917 => x"718287cc",
          1918 => x"0c863d0d",
          1919 => x"04f33d0d",
          1920 => x"7f5b87c0",
          1921 => x"989c5d81",
          1922 => x"7d0c87c0",
          1923 => x"98bc085e",
          1924 => x"7d7b2387",
          1925 => x"c098b808",
          1926 => x"5a79821c",
          1927 => x"3487c098",
          1928 => x"b4085a79",
          1929 => x"831c3487",
          1930 => x"c098b008",
          1931 => x"5a79841c",
          1932 => x"3487c098",
          1933 => x"ac085a79",
          1934 => x"851c3487",
          1935 => x"c098a808",
          1936 => x"5a79861c",
          1937 => x"3487c098",
          1938 => x"a4085c7b",
          1939 => x"881c2387",
          1940 => x"c098a008",
          1941 => x"5a798a1c",
          1942 => x"23807d0c",
          1943 => x"7983ffff",
          1944 => x"06597b83",
          1945 => x"ffff0658",
          1946 => x"861b3357",
          1947 => x"851b3356",
          1948 => x"841b3355",
          1949 => x"831b3354",
          1950 => x"821b3353",
          1951 => x"7d83ffff",
          1952 => x"065281f6",
          1953 => x"e85194fc",
          1954 => x"3f8f3d0d",
          1955 => x"04ff3d0d",
          1956 => x"028f0533",
          1957 => x"7030709f",
          1958 => x"2a515252",
          1959 => x"708285ec",
          1960 => x"34833d0d",
          1961 => x"04fb3d0d",
          1962 => x"778285ec",
          1963 => x"337081ff",
          1964 => x"06575556",
          1965 => x"87c09484",
          1966 => x"5174802e",
          1967 => x"863887c0",
          1968 => x"94945170",
          1969 => x"0870962a",
          1970 => x"70810653",
          1971 => x"54527080",
          1972 => x"2e8c3871",
          1973 => x"912a7081",
          1974 => x"06515170",
          1975 => x"d7387281",
          1976 => x"32708106",
          1977 => x"51517080",
          1978 => x"2e8d3871",
          1979 => x"932a7081",
          1980 => x"06515170",
          1981 => x"ffbe3873",
          1982 => x"81ff0651",
          1983 => x"87c09480",
          1984 => x"5270802e",
          1985 => x"863887c0",
          1986 => x"94905275",
          1987 => x"720c7582",
          1988 => x"87cc0c87",
          1989 => x"3d0d04fb",
          1990 => x"3d0d029f",
          1991 => x"05338285",
          1992 => x"ec337081",
          1993 => x"ff065755",
          1994 => x"5687c094",
          1995 => x"84517480",
          1996 => x"2e863887",
          1997 => x"c0949451",
          1998 => x"70087096",
          1999 => x"2a708106",
          2000 => x"53545270",
          2001 => x"802e8c38",
          2002 => x"71912a70",
          2003 => x"81065151",
          2004 => x"70d73872",
          2005 => x"81327081",
          2006 => x"06515170",
          2007 => x"802e8d38",
          2008 => x"71932a70",
          2009 => x"81065151",
          2010 => x"70ffbe38",
          2011 => x"7381ff06",
          2012 => x"5187c094",
          2013 => x"80527080",
          2014 => x"2e863887",
          2015 => x"c0949052",
          2016 => x"75720c87",
          2017 => x"3d0d04f9",
          2018 => x"3d0d7954",
          2019 => x"80743370",
          2020 => x"81ff0653",
          2021 => x"53577077",
          2022 => x"2e80fc38",
          2023 => x"7181ff06",
          2024 => x"81158285",
          2025 => x"ec337081",
          2026 => x"ff065957",
          2027 => x"555887c0",
          2028 => x"94845175",
          2029 => x"802e8638",
          2030 => x"87c09494",
          2031 => x"51700870",
          2032 => x"962a7081",
          2033 => x"06535452",
          2034 => x"70802e8c",
          2035 => x"3871912a",
          2036 => x"70810651",
          2037 => x"5170d738",
          2038 => x"72813270",
          2039 => x"81065151",
          2040 => x"70802e8d",
          2041 => x"3871932a",
          2042 => x"70810651",
          2043 => x"5170ffbe",
          2044 => x"387481ff",
          2045 => x"065187c0",
          2046 => x"94805270",
          2047 => x"802e8638",
          2048 => x"87c09490",
          2049 => x"5277720c",
          2050 => x"81177433",
          2051 => x"7081ff06",
          2052 => x"53535770",
          2053 => x"ff863876",
          2054 => x"8287cc0c",
          2055 => x"893d0d04",
          2056 => x"fe3d0d82",
          2057 => x"85ec3370",
          2058 => x"81ff0654",
          2059 => x"5287c094",
          2060 => x"84517280",
          2061 => x"2e863887",
          2062 => x"c0949451",
          2063 => x"70087082",
          2064 => x"2a708106",
          2065 => x"51515170",
          2066 => x"802ee238",
          2067 => x"7181ff06",
          2068 => x"5187c094",
          2069 => x"80527080",
          2070 => x"2e863887",
          2071 => x"c0949052",
          2072 => x"71087081",
          2073 => x"ff068287",
          2074 => x"cc0c5184",
          2075 => x"3d0d04fe",
          2076 => x"3d0d8285",
          2077 => x"ec337081",
          2078 => x"ff065253",
          2079 => x"87c09484",
          2080 => x"5270802e",
          2081 => x"863887c0",
          2082 => x"94945271",
          2083 => x"0870822a",
          2084 => x"70810651",
          2085 => x"5151ff52",
          2086 => x"70802ea0",
          2087 => x"387281ff",
          2088 => x"065187c0",
          2089 => x"94805270",
          2090 => x"802e8638",
          2091 => x"87c09490",
          2092 => x"52710870",
          2093 => x"982b7098",
          2094 => x"2c515351",
          2095 => x"718287cc",
          2096 => x"0c843d0d",
          2097 => x"04ff3d0d",
          2098 => x"87c09e80",
          2099 => x"08709c2a",
          2100 => x"8a065151",
          2101 => x"70802e84",
          2102 => x"b43887c0",
          2103 => x"9ea40882",
          2104 => x"85f00c87",
          2105 => x"c09ea808",
          2106 => x"8285f40c",
          2107 => x"87c09e94",
          2108 => x"088285f8",
          2109 => x"0c87c09e",
          2110 => x"98088285",
          2111 => x"fc0c87c0",
          2112 => x"9e9c0882",
          2113 => x"86800c87",
          2114 => x"c09ea008",
          2115 => x"8286840c",
          2116 => x"87c09eac",
          2117 => x"08828688",
          2118 => x"0c87c09e",
          2119 => x"b0088286",
          2120 => x"8c0c87c0",
          2121 => x"9eb40882",
          2122 => x"86900c87",
          2123 => x"c09eb808",
          2124 => x"8286940c",
          2125 => x"87c09ebc",
          2126 => x"08828698",
          2127 => x"0c87c09e",
          2128 => x"c0088286",
          2129 => x"9c0c87c0",
          2130 => x"9ec40882",
          2131 => x"86a00c87",
          2132 => x"c09e8008",
          2133 => x"51708286",
          2134 => x"a42387c0",
          2135 => x"9e840882",
          2136 => x"86a80c87",
          2137 => x"c09e8808",
          2138 => x"8286ac0c",
          2139 => x"87c09e8c",
          2140 => x"088286b0",
          2141 => x"0c810b82",
          2142 => x"86b43480",
          2143 => x"0b87c09e",
          2144 => x"90087084",
          2145 => x"800a0651",
          2146 => x"52527080",
          2147 => x"2e833881",
          2148 => x"52718286",
          2149 => x"b534800b",
          2150 => x"87c09e90",
          2151 => x"08708880",
          2152 => x"0a065152",
          2153 => x"5270802e",
          2154 => x"83388152",
          2155 => x"718286b6",
          2156 => x"34800b87",
          2157 => x"c09e9008",
          2158 => x"7090800a",
          2159 => x"06515252",
          2160 => x"70802e83",
          2161 => x"38815271",
          2162 => x"8286b734",
          2163 => x"800b87c0",
          2164 => x"9e900870",
          2165 => x"88808006",
          2166 => x"51525270",
          2167 => x"802e8338",
          2168 => x"81527182",
          2169 => x"86b83480",
          2170 => x"0b87c09e",
          2171 => x"900870a0",
          2172 => x"80800651",
          2173 => x"52527080",
          2174 => x"2e833881",
          2175 => x"52718286",
          2176 => x"b934800b",
          2177 => x"87c09e90",
          2178 => x"08709080",
          2179 => x"80065152",
          2180 => x"5270802e",
          2181 => x"83388152",
          2182 => x"718286ba",
          2183 => x"34800b87",
          2184 => x"c09e9008",
          2185 => x"70848080",
          2186 => x"06515252",
          2187 => x"70802e83",
          2188 => x"38815271",
          2189 => x"8286bb34",
          2190 => x"800b87c0",
          2191 => x"9e900870",
          2192 => x"82808006",
          2193 => x"51525270",
          2194 => x"802e8338",
          2195 => x"81527182",
          2196 => x"86bc3480",
          2197 => x"0b87c09e",
          2198 => x"90087081",
          2199 => x"80800651",
          2200 => x"52527080",
          2201 => x"2e833881",
          2202 => x"52718286",
          2203 => x"bd34800b",
          2204 => x"87c09e90",
          2205 => x"087080c0",
          2206 => x"80065152",
          2207 => x"5270802e",
          2208 => x"83388152",
          2209 => x"718286be",
          2210 => x"34800b87",
          2211 => x"c09e9008",
          2212 => x"70a08006",
          2213 => x"51525270",
          2214 => x"802e8338",
          2215 => x"81527182",
          2216 => x"86bf3487",
          2217 => x"c09e9008",
          2218 => x"70988006",
          2219 => x"708a2a51",
          2220 => x"51517082",
          2221 => x"86c03480",
          2222 => x"0b87c09e",
          2223 => x"90087084",
          2224 => x"80065152",
          2225 => x"5270802e",
          2226 => x"83388152",
          2227 => x"718286c1",
          2228 => x"3487c09e",
          2229 => x"90087083",
          2230 => x"f0067084",
          2231 => x"2a515151",
          2232 => x"708286c2",
          2233 => x"34800b87",
          2234 => x"c09e9008",
          2235 => x"70880651",
          2236 => x"52527080",
          2237 => x"2e833881",
          2238 => x"52718286",
          2239 => x"c33487c0",
          2240 => x"9e900870",
          2241 => x"87065151",
          2242 => x"708286c4",
          2243 => x"34833d0d",
          2244 => x"04fb3d0d",
          2245 => x"81f78051",
          2246 => x"86863f82",
          2247 => x"86b43354",
          2248 => x"73802e88",
          2249 => x"3881f794",
          2250 => x"5185f53f",
          2251 => x"81f7a851",
          2252 => x"85ee3f82",
          2253 => x"86b63354",
          2254 => x"73802e93",
          2255 => x"38828690",
          2256 => x"08828694",
          2257 => x"08115452",
          2258 => x"81f7c051",
          2259 => x"8bb63f82",
          2260 => x"86bb3354",
          2261 => x"73802e93",
          2262 => x"38828688",
          2263 => x"0882868c",
          2264 => x"08115452",
          2265 => x"81f7dc51",
          2266 => x"8b9a3f82",
          2267 => x"86b83354",
          2268 => x"73802e93",
          2269 => x"388285f0",
          2270 => x"088285f4",
          2271 => x"08115452",
          2272 => x"81f7f851",
          2273 => x"8afe3f82",
          2274 => x"86b93354",
          2275 => x"73802e93",
          2276 => x"388285f8",
          2277 => x"088285fc",
          2278 => x"08115452",
          2279 => x"81f89451",
          2280 => x"8ae23f82",
          2281 => x"86ba3354",
          2282 => x"73802e93",
          2283 => x"38828680",
          2284 => x"08828684",
          2285 => x"08115452",
          2286 => x"81f8b051",
          2287 => x"8ac63f82",
          2288 => x"86bf3354",
          2289 => x"73802e8d",
          2290 => x"388286c0",
          2291 => x"335281f8",
          2292 => x"cc518ab0",
          2293 => x"3f8286c3",
          2294 => x"33547380",
          2295 => x"2e8d3882",
          2296 => x"86c43352",
          2297 => x"81f8ec51",
          2298 => x"8a9a3f82",
          2299 => x"86c13354",
          2300 => x"73802e8d",
          2301 => x"388286c2",
          2302 => x"335281f9",
          2303 => x"8c518a84",
          2304 => x"3f8286b5",
          2305 => x"33547380",
          2306 => x"2e883881",
          2307 => x"f9ac5184",
          2308 => x"8f3f8286",
          2309 => x"b7335473",
          2310 => x"802e8838",
          2311 => x"81f9c051",
          2312 => x"83fe3f82",
          2313 => x"86bc3354",
          2314 => x"73802e88",
          2315 => x"3881f9cc",
          2316 => x"5183ed3f",
          2317 => x"8286bd33",
          2318 => x"5473802e",
          2319 => x"883881f9",
          2320 => x"d85183dc",
          2321 => x"3f8286be",
          2322 => x"33547380",
          2323 => x"2e883881",
          2324 => x"f9e45183",
          2325 => x"cb3f81f9",
          2326 => x"f05183c4",
          2327 => x"3f828698",
          2328 => x"085281f9",
          2329 => x"fc51899c",
          2330 => x"3f82869c",
          2331 => x"085281fa",
          2332 => x"a4518990",
          2333 => x"3f8286a0",
          2334 => x"085281fa",
          2335 => x"cc518984",
          2336 => x"3f81faf4",
          2337 => x"5183993f",
          2338 => x"8286a422",
          2339 => x"5281fafc",
          2340 => x"5188f13f",
          2341 => x"8286a808",
          2342 => x"56bd84c0",
          2343 => x"527551a2",
          2344 => x"ca3f8287",
          2345 => x"cc08bd84",
          2346 => x"c0297671",
          2347 => x"31545482",
          2348 => x"87cc0852",
          2349 => x"81fba451",
          2350 => x"88ca3f82",
          2351 => x"86bb3354",
          2352 => x"73802ea8",
          2353 => x"388286ac",
          2354 => x"0856bd84",
          2355 => x"c0527551",
          2356 => x"a2993f82",
          2357 => x"87cc08bd",
          2358 => x"84c02976",
          2359 => x"71315454",
          2360 => x"8287cc08",
          2361 => x"5281fbd0",
          2362 => x"5188993f",
          2363 => x"8286b633",
          2364 => x"5473802e",
          2365 => x"a8388286",
          2366 => x"b00856bd",
          2367 => x"84c05275",
          2368 => x"51a1e83f",
          2369 => x"8287cc08",
          2370 => x"bd84c029",
          2371 => x"76713154",
          2372 => x"548287cc",
          2373 => x"085281fb",
          2374 => x"fc5187e8",
          2375 => x"3f81f2e4",
          2376 => x"5181fd3f",
          2377 => x"873d0d04",
          2378 => x"fe3d0d02",
          2379 => x"920533ff",
          2380 => x"05527184",
          2381 => x"26aa3871",
          2382 => x"842981e9",
          2383 => x"94055271",
          2384 => x"080481fc",
          2385 => x"a8519d39",
          2386 => x"81fcb051",
          2387 => x"973981fc",
          2388 => x"b8519139",
          2389 => x"81fcc051",
          2390 => x"8b3981fc",
          2391 => x"c4518539",
          2392 => x"81fccc51",
          2393 => x"81ba3f84",
          2394 => x"3d0d0471",
          2395 => x"88800c04",
          2396 => x"ff3d0d87",
          2397 => x"c0968470",
          2398 => x"08525280",
          2399 => x"720c7074",
          2400 => x"07708286",
          2401 => x"c80c720c",
          2402 => x"833d0d04",
          2403 => x"ff3d0d87",
          2404 => x"c0968470",
          2405 => x"088286c8",
          2406 => x"0c528072",
          2407 => x"0c730970",
          2408 => x"8286c808",
          2409 => x"06708286",
          2410 => x"c80c730c",
          2411 => x"51833d0d",
          2412 => x"04800b87",
          2413 => x"c096840c",
          2414 => x"048286c8",
          2415 => x"0887c096",
          2416 => x"840c04fe",
          2417 => x"3d0d0293",
          2418 => x"05335372",
          2419 => x"8a2e0981",
          2420 => x"0685388d",
          2421 => x"51ed3f82",
          2422 => x"9edc0852",
          2423 => x"71802e90",
          2424 => x"38727234",
          2425 => x"829edc08",
          2426 => x"8105829e",
          2427 => x"dc0c8f39",
          2428 => x"829ed408",
          2429 => x"5271802e",
          2430 => x"85387251",
          2431 => x"712d843d",
          2432 => x"0d04fe3d",
          2433 => x"0d029705",
          2434 => x"33829ed4",
          2435 => x"0876829e",
          2436 => x"d40c5451",
          2437 => x"ffad3f72",
          2438 => x"829ed40c",
          2439 => x"843d0d04",
          2440 => x"fd3d0d75",
          2441 => x"54733370",
          2442 => x"81ff0653",
          2443 => x"5371802e",
          2444 => x"8e387281",
          2445 => x"ff065181",
          2446 => x"1454ff87",
          2447 => x"3fe73985",
          2448 => x"3d0d04fc",
          2449 => x"3d0d7782",
          2450 => x"9ed40878",
          2451 => x"829ed40c",
          2452 => x"56547333",
          2453 => x"7081ff06",
          2454 => x"53537180",
          2455 => x"2e8e3872",
          2456 => x"81ff0651",
          2457 => x"811454fe",
          2458 => x"da3fe739",
          2459 => x"74829ed4",
          2460 => x"0c863d0d",
          2461 => x"04ec3d0d",
          2462 => x"66685959",
          2463 => x"78708105",
          2464 => x"5a335675",
          2465 => x"802e84f8",
          2466 => x"3875a52e",
          2467 => x"09810682",
          2468 => x"de388070",
          2469 => x"7a708105",
          2470 => x"5c33585b",
          2471 => x"5b75b02e",
          2472 => x"09810685",
          2473 => x"38815a8b",
          2474 => x"3975ad2e",
          2475 => x"0981068a",
          2476 => x"38825a78",
          2477 => x"7081055a",
          2478 => x"335675aa",
          2479 => x"2e098106",
          2480 => x"92387784",
          2481 => x"1971087b",
          2482 => x"7081055d",
          2483 => x"33595d59",
          2484 => x"539d39d0",
          2485 => x"16537289",
          2486 => x"2695387a",
          2487 => x"88297b10",
          2488 => x"057605d0",
          2489 => x"05797081",
          2490 => x"055b3357",
          2491 => x"5be53975",
          2492 => x"80ec3270",
          2493 => x"30707207",
          2494 => x"80257880",
          2495 => x"cc327030",
          2496 => x"70720780",
          2497 => x"25730753",
          2498 => x"54585155",
          2499 => x"5373802e",
          2500 => x"8c387984",
          2501 => x"07797081",
          2502 => x"055b3357",
          2503 => x"5a75802e",
          2504 => x"83de3875",
          2505 => x"5480e076",
          2506 => x"278938e0",
          2507 => x"167081ff",
          2508 => x"06555373",
          2509 => x"80cf2e81",
          2510 => x"aa387380",
          2511 => x"cf24a238",
          2512 => x"7380c32e",
          2513 => x"818e3873",
          2514 => x"80c3248b",
          2515 => x"387380c2",
          2516 => x"2e818c38",
          2517 => x"81993973",
          2518 => x"80c42e81",
          2519 => x"8a38818f",
          2520 => x"397380d5",
          2521 => x"2e818038",
          2522 => x"7380d524",
          2523 => x"8a387380",
          2524 => x"d32e8e38",
          2525 => x"80f93973",
          2526 => x"80d82e80",
          2527 => x"ee3880ef",
          2528 => x"39778419",
          2529 => x"71085659",
          2530 => x"53807433",
          2531 => x"54557275",
          2532 => x"2e8d3881",
          2533 => x"15701570",
          2534 => x"33515455",
          2535 => x"72f53879",
          2536 => x"812a5690",
          2537 => x"39748116",
          2538 => x"5653727b",
          2539 => x"278f38a0",
          2540 => x"51fc903f",
          2541 => x"75810653",
          2542 => x"72802ee9",
          2543 => x"387351fc",
          2544 => x"df3f7481",
          2545 => x"16565372",
          2546 => x"7b27fdb0",
          2547 => x"38a051fb",
          2548 => x"f23fef39",
          2549 => x"77841983",
          2550 => x"12335359",
          2551 => x"53933982",
          2552 => x"5c953988",
          2553 => x"5c91398a",
          2554 => x"5c8d3990",
          2555 => x"5c893975",
          2556 => x"51fbd03f",
          2557 => x"fd863979",
          2558 => x"822a7081",
          2559 => x"06515372",
          2560 => x"802e8838",
          2561 => x"77841959",
          2562 => x"53863984",
          2563 => x"18785458",
          2564 => x"72087480",
          2565 => x"c4327030",
          2566 => x"70720780",
          2567 => x"25515555",
          2568 => x"55748025",
          2569 => x"8d387280",
          2570 => x"2e883874",
          2571 => x"307a9007",
          2572 => x"5b55800b",
          2573 => x"8f3d5e57",
          2574 => x"7b527451",
          2575 => x"9dd43f82",
          2576 => x"87cc0881",
          2577 => x"ff067c53",
          2578 => x"7552549b",
          2579 => x"9e3f8287",
          2580 => x"cc085589",
          2581 => x"74279238",
          2582 => x"a7145375",
          2583 => x"80f82e84",
          2584 => x"38871453",
          2585 => x"7281ff06",
          2586 => x"54b01453",
          2587 => x"727d7081",
          2588 => x"055f3481",
          2589 => x"17753070",
          2590 => x"77079f2a",
          2591 => x"51545776",
          2592 => x"9f268538",
          2593 => x"72ffb138",
          2594 => x"79842a70",
          2595 => x"81065153",
          2596 => x"72802e8e",
          2597 => x"38963d77",
          2598 => x"05e00553",
          2599 => x"ad733481",
          2600 => x"1757767a",
          2601 => x"81065455",
          2602 => x"b0547283",
          2603 => x"38a05479",
          2604 => x"812a7081",
          2605 => x"06545672",
          2606 => x"9f388117",
          2607 => x"55767b27",
          2608 => x"97387351",
          2609 => x"f9fd3f75",
          2610 => x"81065372",
          2611 => x"8b387481",
          2612 => x"1656537a",
          2613 => x"7326eb38",
          2614 => x"963d7705",
          2615 => x"e00553ff",
          2616 => x"17ff1470",
          2617 => x"33535457",
          2618 => x"f9d93f76",
          2619 => x"f2387481",
          2620 => x"16565372",
          2621 => x"7b27fb84",
          2622 => x"38a051f9",
          2623 => x"c63fef39",
          2624 => x"963d0d04",
          2625 => x"fd3d0d86",
          2626 => x"3d707084",
          2627 => x"05520855",
          2628 => x"527351fa",
          2629 => x"e03f853d",
          2630 => x"0d04fe3d",
          2631 => x"0d74829e",
          2632 => x"dc0c853d",
          2633 => x"88055275",
          2634 => x"51faca3f",
          2635 => x"829edc08",
          2636 => x"53807334",
          2637 => x"800b829e",
          2638 => x"dc0c843d",
          2639 => x"0d04fd3d",
          2640 => x"0d829ed4",
          2641 => x"0876829e",
          2642 => x"d40c873d",
          2643 => x"88055377",
          2644 => x"5253faa1",
          2645 => x"3f72829e",
          2646 => x"d40c853d",
          2647 => x"0d04fb3d",
          2648 => x"0d777982",
          2649 => x"9ed80870",
          2650 => x"56545755",
          2651 => x"80547180",
          2652 => x"2e80e038",
          2653 => x"829ed808",
          2654 => x"52712d82",
          2655 => x"87cc0881",
          2656 => x"ff065372",
          2657 => x"802e80cb",
          2658 => x"38728d2e",
          2659 => x"b9387288",
          2660 => x"32703070",
          2661 => x"80255151",
          2662 => x"5273802e",
          2663 => x"8b387180",
          2664 => x"2e8638ff",
          2665 => x"14549739",
          2666 => x"9f7325c8",
          2667 => x"38ff1652",
          2668 => x"737225c0",
          2669 => x"38741452",
          2670 => x"72723481",
          2671 => x"14547251",
          2672 => x"f8813fff",
          2673 => x"af397315",
          2674 => x"52807234",
          2675 => x"8a51f7f3",
          2676 => x"3f815372",
          2677 => x"8287cc0c",
          2678 => x"873d0d04",
          2679 => x"fe3d0d82",
          2680 => x"9ed80875",
          2681 => x"829ed80c",
          2682 => x"77537652",
          2683 => x"53feef3f",
          2684 => x"72829ed8",
          2685 => x"0c843d0d",
          2686 => x"04f83d0d",
          2687 => x"7a7c5a56",
          2688 => x"80707a0c",
          2689 => x"58750870",
          2690 => x"33555373",
          2691 => x"a02e0981",
          2692 => x"06873881",
          2693 => x"13760ced",
          2694 => x"3973ad2e",
          2695 => x"0981068e",
          2696 => x"38817608",
          2697 => x"11770c76",
          2698 => x"08703356",
          2699 => x"545873b0",
          2700 => x"2e098106",
          2701 => x"80c23875",
          2702 => x"08810576",
          2703 => x"0c750870",
          2704 => x"33555373",
          2705 => x"80e22e8b",
          2706 => x"38905773",
          2707 => x"80f82e85",
          2708 => x"388f3982",
          2709 => x"57811376",
          2710 => x"0c750870",
          2711 => x"335553ac",
          2712 => x"398155a0",
          2713 => x"742780fa",
          2714 => x"38d01453",
          2715 => x"80558857",
          2716 => x"89732798",
          2717 => x"3880eb39",
          2718 => x"d0145380",
          2719 => x"55728926",
          2720 => x"80e03886",
          2721 => x"39805580",
          2722 => x"d9398a57",
          2723 => x"8055a074",
          2724 => x"2780c238",
          2725 => x"80e07427",
          2726 => x"8938e014",
          2727 => x"7081ff06",
          2728 => x"5553d014",
          2729 => x"7081ff06",
          2730 => x"55539074",
          2731 => x"278e38f9",
          2732 => x"147081ff",
          2733 => x"06555389",
          2734 => x"7427ca38",
          2735 => x"737727c5",
          2736 => x"38747729",
          2737 => x"14760881",
          2738 => x"05770c76",
          2739 => x"08703356",
          2740 => x"5455ffba",
          2741 => x"3977802e",
          2742 => x"84387430",
          2743 => x"5574790c",
          2744 => x"81557482",
          2745 => x"87cc0c8a",
          2746 => x"3d0d04f8",
          2747 => x"3d0d7a7c",
          2748 => x"5a568070",
          2749 => x"7a0c5875",
          2750 => x"08703355",
          2751 => x"5373a02e",
          2752 => x"09810687",
          2753 => x"38811376",
          2754 => x"0ced3973",
          2755 => x"ad2e0981",
          2756 => x"068e3881",
          2757 => x"76081177",
          2758 => x"0c760870",
          2759 => x"33565458",
          2760 => x"73b02e09",
          2761 => x"810680c2",
          2762 => x"38750881",
          2763 => x"05760c75",
          2764 => x"08703355",
          2765 => x"537380e2",
          2766 => x"2e8b3890",
          2767 => x"577380f8",
          2768 => x"2e85388f",
          2769 => x"39825781",
          2770 => x"13760c75",
          2771 => x"08703355",
          2772 => x"53ac3981",
          2773 => x"55a07427",
          2774 => x"80fa38d0",
          2775 => x"14538055",
          2776 => x"88578973",
          2777 => x"27983880",
          2778 => x"eb39d014",
          2779 => x"53805572",
          2780 => x"892680e0",
          2781 => x"38863980",
          2782 => x"5580d939",
          2783 => x"8a578055",
          2784 => x"a0742780",
          2785 => x"c23880e0",
          2786 => x"74278938",
          2787 => x"e0147081",
          2788 => x"ff065553",
          2789 => x"d0147081",
          2790 => x"ff065553",
          2791 => x"9074278e",
          2792 => x"38f91470",
          2793 => x"81ff0655",
          2794 => x"53897427",
          2795 => x"ca387377",
          2796 => x"27c53874",
          2797 => x"77291476",
          2798 => x"08810577",
          2799 => x"0c760870",
          2800 => x"33565455",
          2801 => x"ffba3977",
          2802 => x"802e8438",
          2803 => x"74305574",
          2804 => x"790c8155",
          2805 => x"748287cc",
          2806 => x"0c8a3d0d",
          2807 => x"04fd3d0d",
          2808 => x"76982b70",
          2809 => x"982c7998",
          2810 => x"2b70982c",
          2811 => x"72101370",
          2812 => x"822b5153",
          2813 => x"51545151",
          2814 => x"800b81fc",
          2815 => x"d8123355",
          2816 => x"53717425",
          2817 => x"9c3881fc",
          2818 => x"d4110812",
          2819 => x"02840597",
          2820 => x"05337133",
          2821 => x"52525270",
          2822 => x"722e0981",
          2823 => x"06833881",
          2824 => x"53728287",
          2825 => x"cc0c853d",
          2826 => x"0d04fc3d",
          2827 => x"0d780284",
          2828 => x"059f0533",
          2829 => x"71335455",
          2830 => x"5371802e",
          2831 => x"9f388851",
          2832 => x"f3813fa0",
          2833 => x"51f2fc3f",
          2834 => x"8851f2f7",
          2835 => x"3f7233ff",
          2836 => x"05527173",
          2837 => x"347181ff",
          2838 => x"0652de39",
          2839 => x"7651f3c0",
          2840 => x"3f737334",
          2841 => x"863d0d04",
          2842 => x"f63d0d7c",
          2843 => x"028405b7",
          2844 => x"05330288",
          2845 => x"05bb0533",
          2846 => x"8287a433",
          2847 => x"70842982",
          2848 => x"86cc0570",
          2849 => x"08515959",
          2850 => x"5a585974",
          2851 => x"802e8638",
          2852 => x"74519e83",
          2853 => x"3f8287a4",
          2854 => x"33708429",
          2855 => x"8286cc05",
          2856 => x"81197054",
          2857 => x"58565aa1",
          2858 => x"843f8287",
          2859 => x"cc08750c",
          2860 => x"8287a433",
          2861 => x"70842982",
          2862 => x"86cc0570",
          2863 => x"0851565a",
          2864 => x"74802ea7",
          2865 => x"38755378",
          2866 => x"527451ff",
          2867 => x"bbc93f82",
          2868 => x"87a43381",
          2869 => x"05557482",
          2870 => x"87a43474",
          2871 => x"81ff0655",
          2872 => x"93752787",
          2873 => x"38800b82",
          2874 => x"87a43477",
          2875 => x"802eb638",
          2876 => x"8287a008",
          2877 => x"5675802e",
          2878 => x"ac388287",
          2879 => x"9c335574",
          2880 => x"a4388c3d",
          2881 => x"fc055476",
          2882 => x"53785275",
          2883 => x"5180d8e9",
          2884 => x"3f8287a0",
          2885 => x"08528a51",
          2886 => x"818df63f",
          2887 => x"8287a008",
          2888 => x"5180dcc6",
          2889 => x"3f8c3d0d",
          2890 => x"04fd3d0d",
          2891 => x"8286cc53",
          2892 => x"93547208",
          2893 => x"5271802e",
          2894 => x"89387151",
          2895 => x"9cd93f80",
          2896 => x"730cff14",
          2897 => x"84145454",
          2898 => x"738025e6",
          2899 => x"38800b82",
          2900 => x"87a43482",
          2901 => x"87a00852",
          2902 => x"71802e95",
          2903 => x"38715180",
          2904 => x"dda63f82",
          2905 => x"87a00851",
          2906 => x"9cad3f80",
          2907 => x"0b8287a0",
          2908 => x"0c853d0d",
          2909 => x"04dc3d0d",
          2910 => x"81578052",
          2911 => x"8287a008",
          2912 => x"5180e293",
          2913 => x"3f8287cc",
          2914 => x"0880d238",
          2915 => x"8287a008",
          2916 => x"5380f852",
          2917 => x"883d7052",
          2918 => x"56818ae1",
          2919 => x"3f8287cc",
          2920 => x"08802eb9",
          2921 => x"387551ff",
          2922 => x"b88d3f82",
          2923 => x"87cc0855",
          2924 => x"800b8287",
          2925 => x"cc08259c",
          2926 => x"388287cc",
          2927 => x"08ff0570",
          2928 => x"17555580",
          2929 => x"74347553",
          2930 => x"76528117",
          2931 => x"81ffc852",
          2932 => x"57f6b13f",
          2933 => x"74ff2e09",
          2934 => x"8106ffb0",
          2935 => x"38a63d0d",
          2936 => x"04d93d0d",
          2937 => x"aa3d08ad",
          2938 => x"3d085a5a",
          2939 => x"81705858",
          2940 => x"80528287",
          2941 => x"a0085180",
          2942 => x"e19d3f82",
          2943 => x"87cc0881",
          2944 => x"9438ff0b",
          2945 => x"8287a008",
          2946 => x"545580f8",
          2947 => x"528b3d70",
          2948 => x"52568189",
          2949 => x"e83f8287",
          2950 => x"cc08802e",
          2951 => x"a5387551",
          2952 => x"ffb7943f",
          2953 => x"8287cc08",
          2954 => x"81185855",
          2955 => x"800b8287",
          2956 => x"cc08258e",
          2957 => x"388287cc",
          2958 => x"08ff0570",
          2959 => x"17555580",
          2960 => x"74347409",
          2961 => x"70307072",
          2962 => x"079f2a51",
          2963 => x"55557877",
          2964 => x"2e853873",
          2965 => x"ffac3882",
          2966 => x"87a0088c",
          2967 => x"11085351",
          2968 => x"80e0b43f",
          2969 => x"8287cc08",
          2970 => x"802e8838",
          2971 => x"81ffd451",
          2972 => x"efae3f78",
          2973 => x"772e0981",
          2974 => x"069b3875",
          2975 => x"527951ff",
          2976 => x"b7a33f79",
          2977 => x"51ffb6af",
          2978 => x"3fab3d08",
          2979 => x"548287cc",
          2980 => x"08743480",
          2981 => x"58778287",
          2982 => x"cc0ca93d",
          2983 => x"0d04f63d",
          2984 => x"0d7c7e71",
          2985 => x"5c717233",
          2986 => x"57595a58",
          2987 => x"73a02e09",
          2988 => x"8106a238",
          2989 => x"78337805",
          2990 => x"56777627",
          2991 => x"98388117",
          2992 => x"705b7071",
          2993 => x"33565855",
          2994 => x"73a02e09",
          2995 => x"81068638",
          2996 => x"757526ea",
          2997 => x"38805473",
          2998 => x"88298287",
          2999 => x"a8057008",
          3000 => x"5255ffb5",
          3001 => x"d23f8287",
          3002 => x"cc085379",
          3003 => x"52740851",
          3004 => x"ffb8d13f",
          3005 => x"8287cc08",
          3006 => x"80c53884",
          3007 => x"15335574",
          3008 => x"812e8838",
          3009 => x"74822e88",
          3010 => x"38b539fc",
          3011 => x"e83fac39",
          3012 => x"811a5a8c",
          3013 => x"3dfc1153",
          3014 => x"f80551f5",
          3015 => x"dc3f8287",
          3016 => x"cc08802e",
          3017 => x"9a38ff1b",
          3018 => x"53785277",
          3019 => x"51fdb23f",
          3020 => x"8287cc08",
          3021 => x"81ff0655",
          3022 => x"74853874",
          3023 => x"54913981",
          3024 => x"147081ff",
          3025 => x"06515482",
          3026 => x"7427ff8b",
          3027 => x"38805473",
          3028 => x"8287cc0c",
          3029 => x"8c3d0d04",
          3030 => x"d33d0db0",
          3031 => x"3d08b23d",
          3032 => x"08b43d08",
          3033 => x"595f5a80",
          3034 => x"0baf3d34",
          3035 => x"8287a433",
          3036 => x"8287a008",
          3037 => x"555b7381",
          3038 => x"ca387382",
          3039 => x"879c3355",
          3040 => x"55738338",
          3041 => x"81557680",
          3042 => x"2e81bb38",
          3043 => x"81707606",
          3044 => x"55567380",
          3045 => x"2e81ac38",
          3046 => x"a8519b91",
          3047 => x"3f8287cc",
          3048 => x"088287a0",
          3049 => x"0c8287cc",
          3050 => x"08802e81",
          3051 => x"91389353",
          3052 => x"76528287",
          3053 => x"cc085180",
          3054 => x"cbdd3f82",
          3055 => x"87cc0880",
          3056 => x"2e8b3882",
          3057 => x"808051f2",
          3058 => x"bb3f80f7",
          3059 => x"398287cc",
          3060 => x"085b8287",
          3061 => x"a0085380",
          3062 => x"f852903d",
          3063 => x"70525481",
          3064 => x"869b3f82",
          3065 => x"87cc0856",
          3066 => x"8287cc08",
          3067 => x"742e0981",
          3068 => x"0680d038",
          3069 => x"8287cc08",
          3070 => x"51ffb3bb",
          3071 => x"3f8287cc",
          3072 => x"0855800b",
          3073 => x"8287cc08",
          3074 => x"25a93882",
          3075 => x"87cc08ff",
          3076 => x"05701755",
          3077 => x"55807434",
          3078 => x"80537481",
          3079 => x"ff065275",
          3080 => x"51f8c53f",
          3081 => x"811b7081",
          3082 => x"ff065c54",
          3083 => x"937b2783",
          3084 => x"38805b74",
          3085 => x"ff2e0981",
          3086 => x"06ff9738",
          3087 => x"86397582",
          3088 => x"879c3476",
          3089 => x"8c388287",
          3090 => x"a008802e",
          3091 => x"8438f9d9",
          3092 => x"3f8f3d5d",
          3093 => x"e0993f82",
          3094 => x"87cc0898",
          3095 => x"2b70982c",
          3096 => x"515978ff",
          3097 => x"2eee3878",
          3098 => x"81ff0682",
          3099 => x"9ee43370",
          3100 => x"982b7098",
          3101 => x"2c829ee0",
          3102 => x"3370982b",
          3103 => x"70972c71",
          3104 => x"982c0570",
          3105 => x"842981fc",
          3106 => x"d4057008",
          3107 => x"15703351",
          3108 => x"51515159",
          3109 => x"5951595d",
          3110 => x"58815673",
          3111 => x"782e80e9",
          3112 => x"38777427",
          3113 => x"b4387481",
          3114 => x"800a2981",
          3115 => x"ff0a0570",
          3116 => x"982c5155",
          3117 => x"80752480",
          3118 => x"ce387653",
          3119 => x"74527751",
          3120 => x"f69b3f82",
          3121 => x"87cc0881",
          3122 => x"ff065473",
          3123 => x"802ed738",
          3124 => x"74829ee0",
          3125 => x"348156b1",
          3126 => x"39748180",
          3127 => x"0a298180",
          3128 => x"0a057098",
          3129 => x"2c7081ff",
          3130 => x"06565155",
          3131 => x"73952697",
          3132 => x"38765374",
          3133 => x"527751f5",
          3134 => x"e43f8287",
          3135 => x"cc0881ff",
          3136 => x"065473cc",
          3137 => x"38d33980",
          3138 => x"5675802e",
          3139 => x"80ca3881",
          3140 => x"1c557482",
          3141 => x"9ee43474",
          3142 => x"982b7098",
          3143 => x"2c829ee0",
          3144 => x"3370982b",
          3145 => x"70982c70",
          3146 => x"10117082",
          3147 => x"2b81fcd8",
          3148 => x"11335e51",
          3149 => x"51515758",
          3150 => x"51557477",
          3151 => x"2e098106",
          3152 => x"fe923881",
          3153 => x"fcdc1408",
          3154 => x"7d0c800b",
          3155 => x"829ee434",
          3156 => x"800b829e",
          3157 => x"e0349239",
          3158 => x"75829ee4",
          3159 => x"3475829e",
          3160 => x"e03478af",
          3161 => x"3d34757d",
          3162 => x"0c7e5473",
          3163 => x"9526fde1",
          3164 => x"38738429",
          3165 => x"81e9a805",
          3166 => x"54730804",
          3167 => x"829eec33",
          3168 => x"54737e2e",
          3169 => x"fdcb3882",
          3170 => x"9ee83355",
          3171 => x"737527ab",
          3172 => x"3874982b",
          3173 => x"70982c51",
          3174 => x"55737524",
          3175 => x"9e38741a",
          3176 => x"54733381",
          3177 => x"15347481",
          3178 => x"800a2981",
          3179 => x"ff0a0570",
          3180 => x"982c829e",
          3181 => x"ec335651",
          3182 => x"55df3982",
          3183 => x"9eec3381",
          3184 => x"11565474",
          3185 => x"829eec34",
          3186 => x"731a54ae",
          3187 => x"3d337434",
          3188 => x"829ee833",
          3189 => x"54737e25",
          3190 => x"89388114",
          3191 => x"5473829e",
          3192 => x"e834829e",
          3193 => x"ec337081",
          3194 => x"800a2981",
          3195 => x"ff0a0570",
          3196 => x"982c829e",
          3197 => x"e8335a51",
          3198 => x"56567477",
          3199 => x"25a23874",
          3200 => x"1a703352",
          3201 => x"54e7bc3f",
          3202 => x"7481800a",
          3203 => x"2981800a",
          3204 => x"0570982c",
          3205 => x"829ee833",
          3206 => x"56515573",
          3207 => x"7524e038",
          3208 => x"829eec33",
          3209 => x"70982b70",
          3210 => x"982c829e",
          3211 => x"e8335a51",
          3212 => x"56567477",
          3213 => x"25fc9a38",
          3214 => x"8851e787",
          3215 => x"3f748180",
          3216 => x"0a298180",
          3217 => x"0a057098",
          3218 => x"2c829ee8",
          3219 => x"33565155",
          3220 => x"737524e4",
          3221 => x"38fbfa39",
          3222 => x"837a3480",
          3223 => x"0b811b34",
          3224 => x"829eec53",
          3225 => x"805281f5",
          3226 => x"b851f3be",
          3227 => x"3f81df39",
          3228 => x"829eec33",
          3229 => x"7081ff06",
          3230 => x"55557380",
          3231 => x"2efbd238",
          3232 => x"829ee833",
          3233 => x"ff055473",
          3234 => x"829ee834",
          3235 => x"ff155473",
          3236 => x"829eec34",
          3237 => x"8851e6ab",
          3238 => x"3f829eec",
          3239 => x"3370982b",
          3240 => x"70982c82",
          3241 => x"9ee83357",
          3242 => x"51565774",
          3243 => x"7425a738",
          3244 => x"741a5481",
          3245 => x"14337434",
          3246 => x"733351e6",
          3247 => x"863f7481",
          3248 => x"800a2981",
          3249 => x"800a0570",
          3250 => x"982c829e",
          3251 => x"e8335851",
          3252 => x"55757524",
          3253 => x"db38a051",
          3254 => x"e5e93f82",
          3255 => x"9eec3370",
          3256 => x"982b7098",
          3257 => x"2c829ee8",
          3258 => x"33575156",
          3259 => x"57747424",
          3260 => x"fadf3888",
          3261 => x"51e5cc3f",
          3262 => x"7481800a",
          3263 => x"2981800a",
          3264 => x"0570982c",
          3265 => x"829ee833",
          3266 => x"58515575",
          3267 => x"7525e438",
          3268 => x"fabf3982",
          3269 => x"9ee8337a",
          3270 => x"05548074",
          3271 => x"348a51e5",
          3272 => x"a23f829e",
          3273 => x"e8527951",
          3274 => x"f6f43f82",
          3275 => x"87cc0881",
          3276 => x"ff065473",
          3277 => x"9638829e",
          3278 => x"e8335473",
          3279 => x"802e8f38",
          3280 => x"81537352",
          3281 => x"7951f2a0",
          3282 => x"3f843980",
          3283 => x"7a34800b",
          3284 => x"829eec34",
          3285 => x"800b829e",
          3286 => x"e8347982",
          3287 => x"87cc0caf",
          3288 => x"3d0d0482",
          3289 => x"9eec3354",
          3290 => x"73802ef9",
          3291 => x"e4388851",
          3292 => x"e4d13f82",
          3293 => x"9eec33ff",
          3294 => x"05547382",
          3295 => x"9eec3473",
          3296 => x"81ff0654",
          3297 => x"e339829e",
          3298 => x"ec33829e",
          3299 => x"e8335555",
          3300 => x"73752ef9",
          3301 => x"bc38ff14",
          3302 => x"5473829e",
          3303 => x"e8347498",
          3304 => x"2b70982c",
          3305 => x"7581ff06",
          3306 => x"56515574",
          3307 => x"7425a738",
          3308 => x"741a5481",
          3309 => x"14337434",
          3310 => x"733351e4",
          3311 => x"863f7481",
          3312 => x"800a2981",
          3313 => x"800a0570",
          3314 => x"982c829e",
          3315 => x"e8335851",
          3316 => x"55757524",
          3317 => x"db38a051",
          3318 => x"e3e93f82",
          3319 => x"9eec3370",
          3320 => x"982b7098",
          3321 => x"2c829ee8",
          3322 => x"33575156",
          3323 => x"57747424",
          3324 => x"f8df3888",
          3325 => x"51e3cc3f",
          3326 => x"7481800a",
          3327 => x"2981800a",
          3328 => x"0570982c",
          3329 => x"829ee833",
          3330 => x"58515575",
          3331 => x"7525e438",
          3332 => x"f8bf3982",
          3333 => x"9eec3370",
          3334 => x"81ff0682",
          3335 => x"9ee83359",
          3336 => x"56547477",
          3337 => x"27f8aa38",
          3338 => x"81145473",
          3339 => x"829eec34",
          3340 => x"741a7033",
          3341 => x"5254e38b",
          3342 => x"3f829eec",
          3343 => x"337081ff",
          3344 => x"06829ee8",
          3345 => x"33585654",
          3346 => x"757526dc",
          3347 => x"38f88239",
          3348 => x"829eec53",
          3349 => x"805281f5",
          3350 => x"b851efce",
          3351 => x"3f800b82",
          3352 => x"9eec3480",
          3353 => x"0b829ee8",
          3354 => x"34f7e639",
          3355 => x"7ab03882",
          3356 => x"87980855",
          3357 => x"74802ea6",
          3358 => x"387451ff",
          3359 => x"aab93f82",
          3360 => x"87cc0882",
          3361 => x"9ee83482",
          3362 => x"87cc0881",
          3363 => x"ff068105",
          3364 => x"53745279",
          3365 => x"51ffabff",
          3366 => x"3f935b81",
          3367 => x"c0397a84",
          3368 => x"298286cc",
          3369 => x"05fc1108",
          3370 => x"56547480",
          3371 => x"2ea73874",
          3372 => x"51ffaa83",
          3373 => x"3f8287cc",
          3374 => x"08829ee8",
          3375 => x"348287cc",
          3376 => x"0881ff06",
          3377 => x"81055374",
          3378 => x"527951ff",
          3379 => x"abc93fff",
          3380 => x"1b5480fa",
          3381 => x"39730855",
          3382 => x"74802ef6",
          3383 => x"f4387451",
          3384 => x"ffa9d43f",
          3385 => x"99397a93",
          3386 => x"2e098106",
          3387 => x"ae388286",
          3388 => x"cc085574",
          3389 => x"802ea438",
          3390 => x"7451ffa9",
          3391 => x"ba3f8287",
          3392 => x"cc08829e",
          3393 => x"e8348287",
          3394 => x"cc0881ff",
          3395 => x"06810553",
          3396 => x"74527951",
          3397 => x"ffab803f",
          3398 => x"80c3397a",
          3399 => x"84298286",
          3400 => x"d0057008",
          3401 => x"56547480",
          3402 => x"2eab3874",
          3403 => x"51ffa987",
          3404 => x"3f8287cc",
          3405 => x"08829ee8",
          3406 => x"348287cc",
          3407 => x"0881ff06",
          3408 => x"81055374",
          3409 => x"527951ff",
          3410 => x"aacd3f81",
          3411 => x"1b547381",
          3412 => x"ff065b89",
          3413 => x"3974829e",
          3414 => x"e834747a",
          3415 => x"34829eec",
          3416 => x"53829ee8",
          3417 => x"33527951",
          3418 => x"edc03ff5",
          3419 => x"e439829e",
          3420 => x"ec337081",
          3421 => x"ff06829e",
          3422 => x"e8335956",
          3423 => x"54747727",
          3424 => x"f5cf3881",
          3425 => x"14547382",
          3426 => x"9eec3474",
          3427 => x"1a703352",
          3428 => x"54e0b03f",
          3429 => x"f5bb3982",
          3430 => x"9eec3354",
          3431 => x"73802ef5",
          3432 => x"b0388851",
          3433 => x"e09d3f82",
          3434 => x"9eec33ff",
          3435 => x"05547382",
          3436 => x"9eec34f5",
          3437 => x"9c39fb3d",
          3438 => x"0d779f2c",
          3439 => x"799f2c79",
          3440 => x"9f2c7a32",
          3441 => x"7073317c",
          3442 => x"9f2c7d32",
          3443 => x"74743271",
          3444 => x"75315855",
          3445 => x"59545557",
          3446 => x"54913f82",
          3447 => x"87cc0874",
          3448 => x"32743182",
          3449 => x"87cc0c87",
          3450 => x"3d0d04fa",
          3451 => x"3d0d787a",
          3452 => x"5855a052",
          3453 => x"76802e8b",
          3454 => x"38765180",
          3455 => x"f53f8287",
          3456 => x"cc0852e0",
          3457 => x"12537480",
          3458 => x"2e8d3874",
          3459 => x"5180e33f",
          3460 => x"718287cc",
          3461 => x"08315380",
          3462 => x"52729f26",
          3463 => x"80cb3874",
          3464 => x"52729f2e",
          3465 => x"80c33881",
          3466 => x"1375712a",
          3467 => x"a0723177",
          3468 => x"712b5854",
          3469 => x"55538056",
          3470 => x"72762ea8",
          3471 => x"38731075",
          3472 => x"9f2a0775",
          3473 => x"10770778",
          3474 => x"7231ff11",
          3475 => x"9f2c7081",
          3476 => x"067b7206",
          3477 => x"757131ff",
          3478 => x"1a5a5652",
          3479 => x"5a515456",
          3480 => x"5472da38",
          3481 => x"74107607",
          3482 => x"52718287",
          3483 => x"cc0c883d",
          3484 => x"0d04fd3d",
          3485 => x"0d7570fc",
          3486 => x"80800670",
          3487 => x"30707207",
          3488 => x"80257084",
          3489 => x"2b907131",
          3490 => x"75712a56",
          3491 => x"527483fe",
          3492 => x"80067030",
          3493 => x"70802583",
          3494 => x"2b887131",
          3495 => x"78712a59",
          3496 => x"52730577",
          3497 => x"81f00670",
          3498 => x"30708025",
          3499 => x"822b8471",
          3500 => x"317b712a",
          3501 => x"5c527305",
          3502 => x"7a8c0670",
          3503 => x"30708025",
          3504 => x"10827131",
          3505 => x"7e712a70",
          3506 => x"812a8132",
          3507 => x"70810670",
          3508 => x"30827431",
          3509 => x"06751905",
          3510 => x"8287cc0c",
          3511 => x"51525f52",
          3512 => x"41515253",
          3513 => x"51525351",
          3514 => x"52535153",
          3515 => x"5452853d",
          3516 => x"0d04fd3d",
          3517 => x"0d757770",
          3518 => x"54715354",
          3519 => x"54fdb73f",
          3520 => x"8287cc08",
          3521 => x"73297471",
          3522 => x"318287cc",
          3523 => x"0c53853d",
          3524 => x"0d04fa3d",
          3525 => x"0d787a57",
          3526 => x"55a05275",
          3527 => x"802e8b38",
          3528 => x"7551fece",
          3529 => x"3f8287cc",
          3530 => x"0852e012",
          3531 => x"5374802e",
          3532 => x"8d387451",
          3533 => x"febc3f71",
          3534 => x"8287cc08",
          3535 => x"31537452",
          3536 => x"729f2680",
          3537 => x"c8388052",
          3538 => x"729f2e80",
          3539 => x"c0388113",
          3540 => x"75712aa0",
          3541 => x"72317771",
          3542 => x"2b585455",
          3543 => x"53805772",
          3544 => x"772ea838",
          3545 => x"7310759f",
          3546 => x"2a077510",
          3547 => x"78077772",
          3548 => x"31ff119f",
          3549 => x"2c708106",
          3550 => x"7a720675",
          3551 => x"7131ff1a",
          3552 => x"5a56525b",
          3553 => x"51545654",
          3554 => x"72da3873",
          3555 => x"52718287",
          3556 => x"cc0c883d",
          3557 => x"0d04f93d",
          3558 => x"0d83c080",
          3559 => x"0b8287c4",
          3560 => x"0c84800b",
          3561 => x"8287c023",
          3562 => x"a0805380",
          3563 => x"5283c080",
          3564 => x"51ffa9b7",
          3565 => x"3f8287c4",
          3566 => x"08548058",
          3567 => x"77743481",
          3568 => x"57768115",
          3569 => x"348287c4",
          3570 => x"08547784",
          3571 => x"15347685",
          3572 => x"15348287",
          3573 => x"c4085477",
          3574 => x"86153476",
          3575 => x"87153482",
          3576 => x"87c40882",
          3577 => x"87c022ff",
          3578 => x"05fe8080",
          3579 => x"077083ff",
          3580 => x"ff067088",
          3581 => x"2a585155",
          3582 => x"56748817",
          3583 => x"34738917",
          3584 => x"348287c0",
          3585 => x"22708829",
          3586 => x"8287c408",
          3587 => x"05f81151",
          3588 => x"55557782",
          3589 => x"15347683",
          3590 => x"1534893d",
          3591 => x"0d04ff3d",
          3592 => x"0d735281",
          3593 => x"51847227",
          3594 => x"8f38fb12",
          3595 => x"832a8211",
          3596 => x"7083ffff",
          3597 => x"06515151",
          3598 => x"708287cc",
          3599 => x"0c833d0d",
          3600 => x"04f93d0d",
          3601 => x"02a60522",
          3602 => x"028405aa",
          3603 => x"05227105",
          3604 => x"8287c408",
          3605 => x"71832b71",
          3606 => x"1174832b",
          3607 => x"73117033",
          3608 => x"81123371",
          3609 => x"882b0702",
          3610 => x"a405ae05",
          3611 => x"227181ff",
          3612 => x"ff060770",
          3613 => x"882a5351",
          3614 => x"5259545b",
          3615 => x"5b575354",
          3616 => x"55717734",
          3617 => x"70811834",
          3618 => x"8287c408",
          3619 => x"1475882a",
          3620 => x"52547082",
          3621 => x"15347483",
          3622 => x"15348287",
          3623 => x"c4087017",
          3624 => x"70338112",
          3625 => x"3371882b",
          3626 => x"0770832b",
          3627 => x"8ffff806",
          3628 => x"51525652",
          3629 => x"71057383",
          3630 => x"ffff0670",
          3631 => x"882a5454",
          3632 => x"51718212",
          3633 => x"347281ff",
          3634 => x"06537283",
          3635 => x"12348287",
          3636 => x"c4081656",
          3637 => x"71763472",
          3638 => x"81173489",
          3639 => x"3d0d04fb",
          3640 => x"3d0d8287",
          3641 => x"c4080284",
          3642 => x"059e0522",
          3643 => x"70832b72",
          3644 => x"11861133",
          3645 => x"87123371",
          3646 => x"8b2b7183",
          3647 => x"2b07585b",
          3648 => x"59525552",
          3649 => x"72058412",
          3650 => x"33851333",
          3651 => x"71882b07",
          3652 => x"70882a54",
          3653 => x"56565270",
          3654 => x"84133473",
          3655 => x"85133482",
          3656 => x"87c40870",
          3657 => x"14841133",
          3658 => x"85123371",
          3659 => x"8b2b7183",
          3660 => x"2b075659",
          3661 => x"57527205",
          3662 => x"86123387",
          3663 => x"13337188",
          3664 => x"2b077088",
          3665 => x"2a545656",
          3666 => x"52708613",
          3667 => x"34738713",
          3668 => x"348287c4",
          3669 => x"08137033",
          3670 => x"81123371",
          3671 => x"882b0770",
          3672 => x"81ffff06",
          3673 => x"70882a53",
          3674 => x"51535353",
          3675 => x"71733470",
          3676 => x"81143487",
          3677 => x"3d0d04fa",
          3678 => x"3d0d02a2",
          3679 => x"05228287",
          3680 => x"c4087183",
          3681 => x"2b711170",
          3682 => x"33811233",
          3683 => x"71882b07",
          3684 => x"70882915",
          3685 => x"70338112",
          3686 => x"3371982b",
          3687 => x"71902b07",
          3688 => x"535f5355",
          3689 => x"525a5657",
          3690 => x"53547180",
          3691 => x"2580f638",
          3692 => x"7251feab",
          3693 => x"3f8287c4",
          3694 => x"08701670",
          3695 => x"33811233",
          3696 => x"718b2b71",
          3697 => x"832b0774",
          3698 => x"11703381",
          3699 => x"12337188",
          3700 => x"2b077083",
          3701 => x"2b8ffff8",
          3702 => x"06515254",
          3703 => x"51535a58",
          3704 => x"53720574",
          3705 => x"882a5452",
          3706 => x"72821334",
          3707 => x"73831334",
          3708 => x"8287c408",
          3709 => x"70167033",
          3710 => x"81123371",
          3711 => x"8b2b7183",
          3712 => x"2b075659",
          3713 => x"57557205",
          3714 => x"70338112",
          3715 => x"3371882b",
          3716 => x"077081ff",
          3717 => x"ff067088",
          3718 => x"2a575152",
          3719 => x"58527274",
          3720 => x"34718115",
          3721 => x"34883d0d",
          3722 => x"04fb3d0d",
          3723 => x"8287c408",
          3724 => x"0284059e",
          3725 => x"05227083",
          3726 => x"2b721182",
          3727 => x"11338312",
          3728 => x"33718b2b",
          3729 => x"71832b07",
          3730 => x"595b5952",
          3731 => x"56527305",
          3732 => x"71338113",
          3733 => x"3371882b",
          3734 => x"07028c05",
          3735 => x"a2052271",
          3736 => x"0770882a",
          3737 => x"53515353",
          3738 => x"53717334",
          3739 => x"70811434",
          3740 => x"8287c408",
          3741 => x"70157033",
          3742 => x"81123371",
          3743 => x"8b2b7183",
          3744 => x"2b075659",
          3745 => x"57527205",
          3746 => x"82123383",
          3747 => x"13337188",
          3748 => x"2b077088",
          3749 => x"2a545556",
          3750 => x"52708213",
          3751 => x"34728313",
          3752 => x"348287c4",
          3753 => x"08148211",
          3754 => x"33831233",
          3755 => x"71882b07",
          3756 => x"8287cc0c",
          3757 => x"5254873d",
          3758 => x"0d04f73d",
          3759 => x"0d7b8287",
          3760 => x"c4083183",
          3761 => x"2a7083ff",
          3762 => x"ff067053",
          3763 => x"5753fda7",
          3764 => x"3f8287c4",
          3765 => x"0876832b",
          3766 => x"71118211",
          3767 => x"33831233",
          3768 => x"718b2b71",
          3769 => x"832b0775",
          3770 => x"11703381",
          3771 => x"12337198",
          3772 => x"2b71902b",
          3773 => x"07534240",
          3774 => x"51535b58",
          3775 => x"55595472",
          3776 => x"80258d38",
          3777 => x"82808052",
          3778 => x"7551fe9d",
          3779 => x"3f818439",
          3780 => x"84143385",
          3781 => x"1533718b",
          3782 => x"2b71832b",
          3783 => x"07761179",
          3784 => x"882a5351",
          3785 => x"55585576",
          3786 => x"86143475",
          3787 => x"81ff0656",
          3788 => x"75871434",
          3789 => x"8287c408",
          3790 => x"70198412",
          3791 => x"33851333",
          3792 => x"71882b07",
          3793 => x"70882a54",
          3794 => x"575b5653",
          3795 => x"72841634",
          3796 => x"73851634",
          3797 => x"8287c408",
          3798 => x"1853800b",
          3799 => x"86143480",
          3800 => x"0b871434",
          3801 => x"8287c408",
          3802 => x"53768414",
          3803 => x"34758514",
          3804 => x"348287c4",
          3805 => x"08187033",
          3806 => x"81123371",
          3807 => x"882b0770",
          3808 => x"82808007",
          3809 => x"70882a53",
          3810 => x"51555654",
          3811 => x"74743472",
          3812 => x"8115348b",
          3813 => x"3d0d04ff",
          3814 => x"3d0d7352",
          3815 => x"8287c408",
          3816 => x"8438f7f2",
          3817 => x"3f71802e",
          3818 => x"86387151",
          3819 => x"fe8c3f83",
          3820 => x"3d0d04f5",
          3821 => x"3d0d807e",
          3822 => x"5258f8e2",
          3823 => x"3f8287cc",
          3824 => x"0883ffff",
          3825 => x"068287c4",
          3826 => x"08841133",
          3827 => x"85123371",
          3828 => x"882b0770",
          3829 => x"5f595658",
          3830 => x"5a81ffff",
          3831 => x"5975782e",
          3832 => x"80cb3875",
          3833 => x"88291770",
          3834 => x"33811233",
          3835 => x"71882b07",
          3836 => x"7081ffff",
          3837 => x"06793170",
          3838 => x"83ffff06",
          3839 => x"707f2752",
          3840 => x"53515659",
          3841 => x"55777927",
          3842 => x"8a387380",
          3843 => x"2e853875",
          3844 => x"785a5b84",
          3845 => x"15338516",
          3846 => x"3371882b",
          3847 => x"07575475",
          3848 => x"c2387881",
          3849 => x"ffff2e85",
          3850 => x"387a7959",
          3851 => x"56807683",
          3852 => x"2b8287c4",
          3853 => x"08117033",
          3854 => x"81123371",
          3855 => x"882b0770",
          3856 => x"81ffff06",
          3857 => x"51525a56",
          3858 => x"5c557375",
          3859 => x"2e833881",
          3860 => x"55805479",
          3861 => x"782681cc",
          3862 => x"38745474",
          3863 => x"802e81c4",
          3864 => x"38777a2e",
          3865 => x"09810689",
          3866 => x"387551f8",
          3867 => x"f23f81ac",
          3868 => x"39828080",
          3869 => x"53795275",
          3870 => x"51f7c63f",
          3871 => x"8287c408",
          3872 => x"701c8611",
          3873 => x"33871233",
          3874 => x"718b2b71",
          3875 => x"832b0753",
          3876 => x"5a5e5574",
          3877 => x"057a1770",
          3878 => x"83ffff06",
          3879 => x"70882a5c",
          3880 => x"59565478",
          3881 => x"84153476",
          3882 => x"81ff0657",
          3883 => x"76851534",
          3884 => x"8287c408",
          3885 => x"75832b71",
          3886 => x"11721e86",
          3887 => x"11338712",
          3888 => x"3371882b",
          3889 => x"0770882a",
          3890 => x"535b5e53",
          3891 => x"5a565473",
          3892 => x"86193475",
          3893 => x"87193482",
          3894 => x"87c40870",
          3895 => x"1c841133",
          3896 => x"85123371",
          3897 => x"8b2b7183",
          3898 => x"2b07535d",
          3899 => x"5a557405",
          3900 => x"54788615",
          3901 => x"34768715",
          3902 => x"348287c4",
          3903 => x"08701671",
          3904 => x"1d841133",
          3905 => x"85123371",
          3906 => x"882b0770",
          3907 => x"882a535a",
          3908 => x"5f525654",
          3909 => x"73841634",
          3910 => x"75851634",
          3911 => x"8287c408",
          3912 => x"1b840554",
          3913 => x"738287cc",
          3914 => x"0c8d3d0d",
          3915 => x"04fe3d0d",
          3916 => x"74528287",
          3917 => x"c4088438",
          3918 => x"f4dc3f71",
          3919 => x"5371802e",
          3920 => x"8b387151",
          3921 => x"fced3f82",
          3922 => x"87cc0853",
          3923 => x"728287cc",
          3924 => x"0c843d0d",
          3925 => x"04ff3d0d",
          3926 => x"028f0533",
          3927 => x"51815270",
          3928 => x"72268738",
          3929 => x"8287c811",
          3930 => x"33527182",
          3931 => x"87cc0c83",
          3932 => x"3d0d04fc",
          3933 => x"3d0d029b",
          3934 => x"05330284",
          3935 => x"059f0533",
          3936 => x"56538351",
          3937 => x"72812680",
          3938 => x"e0387284",
          3939 => x"2b87c092",
          3940 => x"8c115351",
          3941 => x"88547480",
          3942 => x"2e843881",
          3943 => x"88547372",
          3944 => x"0c87c092",
          3945 => x"8c115181",
          3946 => x"710c850b",
          3947 => x"87c0988c",
          3948 => x"0c705271",
          3949 => x"08708206",
          3950 => x"51517080",
          3951 => x"2e8a3887",
          3952 => x"c0988c08",
          3953 => x"5170ec38",
          3954 => x"7108fc80",
          3955 => x"80065271",
          3956 => x"923887c0",
          3957 => x"988c0851",
          3958 => x"70802e87",
          3959 => x"38718287",
          3960 => x"c8143482",
          3961 => x"87c81333",
          3962 => x"51708287",
          3963 => x"cc0c863d",
          3964 => x"0d04f33d",
          3965 => x"0d606264",
          3966 => x"028c05bf",
          3967 => x"05335740",
          3968 => x"585b8374",
          3969 => x"525afecd",
          3970 => x"3f8287cc",
          3971 => x"0881067a",
          3972 => x"54527181",
          3973 => x"be387172",
          3974 => x"75842b87",
          3975 => x"c0928011",
          3976 => x"87c0928c",
          3977 => x"1287c092",
          3978 => x"8413415a",
          3979 => x"40575a58",
          3980 => x"850b87c0",
          3981 => x"988c0c76",
          3982 => x"7d0c8476",
          3983 => x"0c750870",
          3984 => x"852a7081",
          3985 => x"06515354",
          3986 => x"71802e8e",
          3987 => x"387b0852",
          3988 => x"717b7081",
          3989 => x"055d3481",
          3990 => x"19598074",
          3991 => x"a2065353",
          3992 => x"71732e83",
          3993 => x"38815378",
          3994 => x"83ff268f",
          3995 => x"3872802e",
          3996 => x"8a3887c0",
          3997 => x"988c0852",
          3998 => x"71c33887",
          3999 => x"c0988c08",
          4000 => x"5271802e",
          4001 => x"87387884",
          4002 => x"802e9938",
          4003 => x"81760c87",
          4004 => x"c0928c15",
          4005 => x"53720870",
          4006 => x"82065152",
          4007 => x"71f738ff",
          4008 => x"1a5a8d39",
          4009 => x"84801781",
          4010 => x"197081ff",
          4011 => x"065a5357",
          4012 => x"79802e90",
          4013 => x"3873fc80",
          4014 => x"80065271",
          4015 => x"87387d78",
          4016 => x"26feed38",
          4017 => x"73fc8080",
          4018 => x"06527180",
          4019 => x"2e833881",
          4020 => x"52715372",
          4021 => x"8287cc0c",
          4022 => x"8f3d0d04",
          4023 => x"f33d0d60",
          4024 => x"6264028c",
          4025 => x"05bf0533",
          4026 => x"5740585b",
          4027 => x"83598074",
          4028 => x"5258fce1",
          4029 => x"3f8287cc",
          4030 => x"08810679",
          4031 => x"54527178",
          4032 => x"2e098106",
          4033 => x"81b13877",
          4034 => x"74842b87",
          4035 => x"c0928011",
          4036 => x"87c0928c",
          4037 => x"1287c092",
          4038 => x"84134059",
          4039 => x"5f565a85",
          4040 => x"0b87c098",
          4041 => x"8c0c767d",
          4042 => x"0c82760c",
          4043 => x"80587508",
          4044 => x"70842a70",
          4045 => x"81065153",
          4046 => x"5471802e",
          4047 => x"8c387a70",
          4048 => x"81055c33",
          4049 => x"7c0c8118",
          4050 => x"5873812a",
          4051 => x"70810651",
          4052 => x"5271802e",
          4053 => x"8a3887c0",
          4054 => x"988c0852",
          4055 => x"71d03887",
          4056 => x"c0988c08",
          4057 => x"5271802e",
          4058 => x"87387784",
          4059 => x"802e9938",
          4060 => x"81760c87",
          4061 => x"c0928c15",
          4062 => x"53720870",
          4063 => x"82065152",
          4064 => x"71f738ff",
          4065 => x"19598d39",
          4066 => x"811a7081",
          4067 => x"ff068480",
          4068 => x"19595b52",
          4069 => x"78802e90",
          4070 => x"3873fc80",
          4071 => x"80065271",
          4072 => x"87387d7a",
          4073 => x"26fef838",
          4074 => x"73fc8080",
          4075 => x"06527180",
          4076 => x"2e833881",
          4077 => x"52715372",
          4078 => x"8287cc0c",
          4079 => x"8f3d0d04",
          4080 => x"fa3d0d7a",
          4081 => x"028405a3",
          4082 => x"05330288",
          4083 => x"05a70533",
          4084 => x"71545456",
          4085 => x"57fafe3f",
          4086 => x"8287cc08",
          4087 => x"81065383",
          4088 => x"547280fe",
          4089 => x"38850b87",
          4090 => x"c0988c0c",
          4091 => x"81567176",
          4092 => x"2e80dc38",
          4093 => x"71762493",
          4094 => x"3874842b",
          4095 => x"87c0928c",
          4096 => x"11545471",
          4097 => x"802e8d38",
          4098 => x"80d43971",
          4099 => x"832e80c6",
          4100 => x"3880cb39",
          4101 => x"72087081",
          4102 => x"2a708106",
          4103 => x"51515271",
          4104 => x"802e8a38",
          4105 => x"87c0988c",
          4106 => x"085271e8",
          4107 => x"3887c098",
          4108 => x"8c085271",
          4109 => x"96388173",
          4110 => x"0c87c092",
          4111 => x"8c145372",
          4112 => x"08708206",
          4113 => x"515271f7",
          4114 => x"38963980",
          4115 => x"56923988",
          4116 => x"800a770c",
          4117 => x"85398180",
          4118 => x"770c7256",
          4119 => x"83398456",
          4120 => x"75547382",
          4121 => x"87cc0c88",
          4122 => x"3d0d04fe",
          4123 => x"3d0d7481",
          4124 => x"11337133",
          4125 => x"71882b07",
          4126 => x"8287cc0c",
          4127 => x"5351843d",
          4128 => x"0d04fd3d",
          4129 => x"0d758311",
          4130 => x"33821233",
          4131 => x"71902b71",
          4132 => x"882b0781",
          4133 => x"14337072",
          4134 => x"07882b75",
          4135 => x"33710782",
          4136 => x"87cc0c52",
          4137 => x"53545654",
          4138 => x"52853d0d",
          4139 => x"04ff3d0d",
          4140 => x"73028405",
          4141 => x"92052252",
          4142 => x"52707270",
          4143 => x"81055434",
          4144 => x"70882a51",
          4145 => x"70723483",
          4146 => x"3d0d04ff",
          4147 => x"3d0d7375",
          4148 => x"52527072",
          4149 => x"70810554",
          4150 => x"3470882a",
          4151 => x"51707270",
          4152 => x"81055434",
          4153 => x"70882a51",
          4154 => x"70727081",
          4155 => x"05543470",
          4156 => x"882a5170",
          4157 => x"7234833d",
          4158 => x"0d04fe3d",
          4159 => x"0d767577",
          4160 => x"54545170",
          4161 => x"802e9238",
          4162 => x"71708105",
          4163 => x"53337370",
          4164 => x"81055534",
          4165 => x"ff1151eb",
          4166 => x"39843d0d",
          4167 => x"04fe3d0d",
          4168 => x"75777654",
          4169 => x"52537272",
          4170 => x"70810554",
          4171 => x"34ff1151",
          4172 => x"70f43884",
          4173 => x"3d0d04fc",
          4174 => x"3d0d7877",
          4175 => x"79565653",
          4176 => x"74708105",
          4177 => x"56337470",
          4178 => x"81055633",
          4179 => x"717131ff",
          4180 => x"16565252",
          4181 => x"5272802e",
          4182 => x"86387180",
          4183 => x"2ee23871",
          4184 => x"8287cc0c",
          4185 => x"863d0d04",
          4186 => x"fe3d0d74",
          4187 => x"76545189",
          4188 => x"3971732e",
          4189 => x"8a388111",
          4190 => x"51703352",
          4191 => x"71f33870",
          4192 => x"338287cc",
          4193 => x"0c843d0d",
          4194 => x"04800b82",
          4195 => x"87cc0c04",
          4196 => x"800b8287",
          4197 => x"cc0c04f7",
          4198 => x"3d0d7b56",
          4199 => x"800b8317",
          4200 => x"33565a74",
          4201 => x"7a2e80d6",
          4202 => x"388154b0",
          4203 => x"160853b4",
          4204 => x"16705381",
          4205 => x"17335259",
          4206 => x"faa23f82",
          4207 => x"87cc087a",
          4208 => x"2e098106",
          4209 => x"b7388287",
          4210 => x"cc088317",
          4211 => x"34b01608",
          4212 => x"70a41808",
          4213 => x"319c1808",
          4214 => x"59565874",
          4215 => x"77279f38",
          4216 => x"82163355",
          4217 => x"74822e09",
          4218 => x"81069338",
          4219 => x"81547618",
          4220 => x"53785281",
          4221 => x"163351f9",
          4222 => x"e33f8339",
          4223 => x"815a7982",
          4224 => x"87cc0c8b",
          4225 => x"3d0d04fa",
          4226 => x"3d0d787a",
          4227 => x"56568057",
          4228 => x"74b01708",
          4229 => x"2eaf3875",
          4230 => x"51fefc3f",
          4231 => x"8287cc08",
          4232 => x"578287cc",
          4233 => x"089f3881",
          4234 => x"547453b4",
          4235 => x"16528116",
          4236 => x"3351f7be",
          4237 => x"3f8287cc",
          4238 => x"08802e85",
          4239 => x"38ff5581",
          4240 => x"5774b017",
          4241 => x"0c768287",
          4242 => x"cc0c883d",
          4243 => x"0d04f83d",
          4244 => x"0d7a7052",
          4245 => x"57fec03f",
          4246 => x"8287cc08",
          4247 => x"588287cc",
          4248 => x"08819138",
          4249 => x"76335574",
          4250 => x"832e0981",
          4251 => x"0680f038",
          4252 => x"84173359",
          4253 => x"78812e09",
          4254 => x"810680e3",
          4255 => x"38848053",
          4256 => x"8287cc08",
          4257 => x"52b41770",
          4258 => x"5256fd91",
          4259 => x"3f82d4d5",
          4260 => x"5284b217",
          4261 => x"51fc963f",
          4262 => x"848b85a4",
          4263 => x"d2527551",
          4264 => x"fca93f86",
          4265 => x"8a85e4f2",
          4266 => x"52849817",
          4267 => x"51fc9c3f",
          4268 => x"90170852",
          4269 => x"849c1751",
          4270 => x"fc913f8c",
          4271 => x"17085284",
          4272 => x"a01751fc",
          4273 => x"863fa017",
          4274 => x"08810570",
          4275 => x"b0190c79",
          4276 => x"55537552",
          4277 => x"81173351",
          4278 => x"f8823f77",
          4279 => x"84183480",
          4280 => x"53805281",
          4281 => x"173351f9",
          4282 => x"d73f8287",
          4283 => x"cc08802e",
          4284 => x"83388158",
          4285 => x"778287cc",
          4286 => x"0c8a3d0d",
          4287 => x"04fb3d0d",
          4288 => x"77fe1a98",
          4289 => x"1208fe05",
          4290 => x"55565480",
          4291 => x"56747327",
          4292 => x"8d388a14",
          4293 => x"22757129",
          4294 => x"ac160805",
          4295 => x"57537582",
          4296 => x"87cc0c87",
          4297 => x"3d0d04f9",
          4298 => x"3d0d7a7a",
          4299 => x"70085654",
          4300 => x"57817727",
          4301 => x"81df3876",
          4302 => x"98150827",
          4303 => x"81d738ff",
          4304 => x"74335458",
          4305 => x"72822e80",
          4306 => x"f5387282",
          4307 => x"24893872",
          4308 => x"812e8d38",
          4309 => x"81bf3972",
          4310 => x"832e818e",
          4311 => x"3881b639",
          4312 => x"76812a17",
          4313 => x"70892aa4",
          4314 => x"16080553",
          4315 => x"745255fd",
          4316 => x"963f8287",
          4317 => x"cc08819f",
          4318 => x"387483ff",
          4319 => x"0614b411",
          4320 => x"33811770",
          4321 => x"892aa418",
          4322 => x"08055576",
          4323 => x"54575753",
          4324 => x"fcf53f82",
          4325 => x"87cc0880",
          4326 => x"fe387483",
          4327 => x"ff0614b4",
          4328 => x"11337088",
          4329 => x"2b780779",
          4330 => x"81067184",
          4331 => x"2a5c5258",
          4332 => x"51537280",
          4333 => x"e238759f",
          4334 => x"ff065880",
          4335 => x"da397688",
          4336 => x"2aa41508",
          4337 => x"05527351",
          4338 => x"fcbd3f82",
          4339 => x"87cc0880",
          4340 => x"c6387610",
          4341 => x"83fe0674",
          4342 => x"05b40551",
          4343 => x"f98d3f82",
          4344 => x"87cc0883",
          4345 => x"ffff0658",
          4346 => x"ae397687",
          4347 => x"2aa41508",
          4348 => x"05527351",
          4349 => x"fc913f82",
          4350 => x"87cc089b",
          4351 => x"3876822b",
          4352 => x"83fc0674",
          4353 => x"05b40551",
          4354 => x"f8f83f82",
          4355 => x"87cc08f0",
          4356 => x"0a065883",
          4357 => x"39815877",
          4358 => x"8287cc0c",
          4359 => x"893d0d04",
          4360 => x"f83d0d7a",
          4361 => x"7c7e5a58",
          4362 => x"56825981",
          4363 => x"7727829e",
          4364 => x"38769817",
          4365 => x"08278296",
          4366 => x"38753353",
          4367 => x"72792e81",
          4368 => x"9d387279",
          4369 => x"24893872",
          4370 => x"812e8d38",
          4371 => x"82803972",
          4372 => x"832e81b8",
          4373 => x"3881f739",
          4374 => x"76812a17",
          4375 => x"70892aa4",
          4376 => x"18080553",
          4377 => x"765255fb",
          4378 => x"9e3f8287",
          4379 => x"cc085982",
          4380 => x"87cc0881",
          4381 => x"d9387483",
          4382 => x"ff0616b4",
          4383 => x"05811678",
          4384 => x"81065956",
          4385 => x"54775376",
          4386 => x"802e8f38",
          4387 => x"77842b9f",
          4388 => x"f0067433",
          4389 => x"8f067107",
          4390 => x"51537274",
          4391 => x"34810b83",
          4392 => x"17347489",
          4393 => x"2aa41708",
          4394 => x"05527551",
          4395 => x"fad93f82",
          4396 => x"87cc0859",
          4397 => x"8287cc08",
          4398 => x"81943874",
          4399 => x"83ff0616",
          4400 => x"b4057884",
          4401 => x"2a545476",
          4402 => x"8f387788",
          4403 => x"2a743381",
          4404 => x"f006718f",
          4405 => x"06075153",
          4406 => x"72743480",
          4407 => x"ec397688",
          4408 => x"2aa41708",
          4409 => x"05527551",
          4410 => x"fa9d3f82",
          4411 => x"87cc0859",
          4412 => x"8287cc08",
          4413 => x"80d83877",
          4414 => x"83ffff06",
          4415 => x"52761083",
          4416 => x"fe067605",
          4417 => x"b40551f7",
          4418 => x"a43fbe39",
          4419 => x"76872aa4",
          4420 => x"17080552",
          4421 => x"7551f9ef",
          4422 => x"3f8287cc",
          4423 => x"08598287",
          4424 => x"cc08ab38",
          4425 => x"77f00a06",
          4426 => x"77822b83",
          4427 => x"fc067018",
          4428 => x"b4057054",
          4429 => x"515454f6",
          4430 => x"c93f8287",
          4431 => x"cc088f0a",
          4432 => x"06740752",
          4433 => x"7251f783",
          4434 => x"3f810b83",
          4435 => x"17347882",
          4436 => x"87cc0c8a",
          4437 => x"3d0d04f8",
          4438 => x"3d0d7a7c",
          4439 => x"7e720859",
          4440 => x"56565981",
          4441 => x"7527a438",
          4442 => x"74981708",
          4443 => x"279d3873",
          4444 => x"802eaa38",
          4445 => x"ff537352",
          4446 => x"7551fda4",
          4447 => x"3f8287cc",
          4448 => x"08548287",
          4449 => x"cc0880f2",
          4450 => x"38933982",
          4451 => x"5480eb39",
          4452 => x"815480e6",
          4453 => x"398287cc",
          4454 => x"085480de",
          4455 => x"39745278",
          4456 => x"51fb843f",
          4457 => x"8287cc08",
          4458 => x"588287cc",
          4459 => x"08802e80",
          4460 => x"c7388287",
          4461 => x"cc08812e",
          4462 => x"d2388287",
          4463 => x"cc08ff2e",
          4464 => x"cf388053",
          4465 => x"74527551",
          4466 => x"fcd63f82",
          4467 => x"87cc08c5",
          4468 => x"38981608",
          4469 => x"fe119018",
          4470 => x"08575557",
          4471 => x"74742790",
          4472 => x"38811590",
          4473 => x"170c8416",
          4474 => x"33810754",
          4475 => x"73841734",
          4476 => x"77557678",
          4477 => x"26ffa638",
          4478 => x"80547382",
          4479 => x"87cc0c8a",
          4480 => x"3d0d04f6",
          4481 => x"3d0d7c7e",
          4482 => x"7108595b",
          4483 => x"5b799538",
          4484 => x"8c170858",
          4485 => x"77802e88",
          4486 => x"38981708",
          4487 => x"7826b238",
          4488 => x"8158ae39",
          4489 => x"79527a51",
          4490 => x"f9fd3f81",
          4491 => x"55748287",
          4492 => x"cc082782",
          4493 => x"e0388287",
          4494 => x"cc085582",
          4495 => x"87cc08ff",
          4496 => x"2e82d238",
          4497 => x"98170882",
          4498 => x"87cc0826",
          4499 => x"82c73879",
          4500 => x"58901708",
          4501 => x"70565473",
          4502 => x"802e82b9",
          4503 => x"38777a2e",
          4504 => x"09810680",
          4505 => x"e238811a",
          4506 => x"56981708",
          4507 => x"76268338",
          4508 => x"82567552",
          4509 => x"7a51f9af",
          4510 => x"3f805982",
          4511 => x"87cc0881",
          4512 => x"2e098106",
          4513 => x"86388287",
          4514 => x"cc085982",
          4515 => x"87cc0809",
          4516 => x"70307072",
          4517 => x"07802570",
          4518 => x"7c078287",
          4519 => x"cc085451",
          4520 => x"51555573",
          4521 => x"81ef3882",
          4522 => x"87cc0880",
          4523 => x"2e95388c",
          4524 => x"17085481",
          4525 => x"74279038",
          4526 => x"73981808",
          4527 => x"27893873",
          4528 => x"58853975",
          4529 => x"80db3877",
          4530 => x"56811656",
          4531 => x"98170876",
          4532 => x"26893882",
          4533 => x"56757826",
          4534 => x"81ac3875",
          4535 => x"527a51f8",
          4536 => x"c63f8287",
          4537 => x"cc08802e",
          4538 => x"b8388059",
          4539 => x"8287cc08",
          4540 => x"812e0981",
          4541 => x"06863882",
          4542 => x"87cc0859",
          4543 => x"8287cc08",
          4544 => x"09703070",
          4545 => x"72078025",
          4546 => x"707c0751",
          4547 => x"51555573",
          4548 => x"80f83875",
          4549 => x"782e0981",
          4550 => x"06ffae38",
          4551 => x"735580f5",
          4552 => x"39ff5375",
          4553 => x"527651f9",
          4554 => x"f73f8287",
          4555 => x"cc088287",
          4556 => x"cc083070",
          4557 => x"8287cc08",
          4558 => x"07802551",
          4559 => x"55557980",
          4560 => x"2e943873",
          4561 => x"802e8f38",
          4562 => x"75537952",
          4563 => x"7651f9d0",
          4564 => x"3f8287cc",
          4565 => x"085574a5",
          4566 => x"38758c18",
          4567 => x"0c981708",
          4568 => x"fe059018",
          4569 => x"08565474",
          4570 => x"74268638",
          4571 => x"ff159018",
          4572 => x"0c841733",
          4573 => x"81075473",
          4574 => x"84183497",
          4575 => x"39ff5674",
          4576 => x"812e9038",
          4577 => x"8c398055",
          4578 => x"8c398287",
          4579 => x"cc085585",
          4580 => x"39815675",
          4581 => x"55748287",
          4582 => x"cc0c8c3d",
          4583 => x"0d04f83d",
          4584 => x"0d7a7052",
          4585 => x"55f3f03f",
          4586 => x"8287cc08",
          4587 => x"58815682",
          4588 => x"87cc0880",
          4589 => x"d8387b52",
          4590 => x"7451f6c1",
          4591 => x"3f8287cc",
          4592 => x"088287cc",
          4593 => x"08b0170c",
          4594 => x"59848053",
          4595 => x"7752b415",
          4596 => x"705257f2",
          4597 => x"c83f7756",
          4598 => x"84398116",
          4599 => x"568a1522",
          4600 => x"58757827",
          4601 => x"97388154",
          4602 => x"75195376",
          4603 => x"52811533",
          4604 => x"51ede93f",
          4605 => x"8287cc08",
          4606 => x"802edf38",
          4607 => x"8a152276",
          4608 => x"32703070",
          4609 => x"7207709f",
          4610 => x"2a535156",
          4611 => x"56758287",
          4612 => x"cc0c8a3d",
          4613 => x"0d04f83d",
          4614 => x"0d7a7c71",
          4615 => x"08585657",
          4616 => x"74f0800a",
          4617 => x"2680f138",
          4618 => x"749f0653",
          4619 => x"7280e938",
          4620 => x"7490180c",
          4621 => x"88170854",
          4622 => x"73aa3875",
          4623 => x"33538273",
          4624 => x"278838a8",
          4625 => x"16085473",
          4626 => x"9b387485",
          4627 => x"2a53820b",
          4628 => x"8817225a",
          4629 => x"58727927",
          4630 => x"80fe38a8",
          4631 => x"16089818",
          4632 => x"0c80cd39",
          4633 => x"8a162270",
          4634 => x"892b5458",
          4635 => x"727526b2",
          4636 => x"38735276",
          4637 => x"51f5b03f",
          4638 => x"8287cc08",
          4639 => x"548287cc",
          4640 => x"08ff2ebd",
          4641 => x"38810b82",
          4642 => x"87cc0827",
          4643 => x"8b389816",
          4644 => x"088287cc",
          4645 => x"08268538",
          4646 => x"8258bd39",
          4647 => x"74733155",
          4648 => x"cb397352",
          4649 => x"7551f4d5",
          4650 => x"3f8287cc",
          4651 => x"0898180c",
          4652 => x"7394180c",
          4653 => x"98170853",
          4654 => x"82587280",
          4655 => x"2e9a3885",
          4656 => x"39815894",
          4657 => x"3974892a",
          4658 => x"1398180c",
          4659 => x"7483ff06",
          4660 => x"16b4059c",
          4661 => x"180c8058",
          4662 => x"778287cc",
          4663 => x"0c8a3d0d",
          4664 => x"04f83d0d",
          4665 => x"7a700890",
          4666 => x"1208a005",
          4667 => x"595754f0",
          4668 => x"800a7727",
          4669 => x"8638800b",
          4670 => x"98150c98",
          4671 => x"14085384",
          4672 => x"5572802e",
          4673 => x"81cb3876",
          4674 => x"83ff0658",
          4675 => x"7781b538",
          4676 => x"81139815",
          4677 => x"0c941408",
          4678 => x"55749238",
          4679 => x"76852a88",
          4680 => x"17225653",
          4681 => x"74732681",
          4682 => x"9b3880c0",
          4683 => x"398a1622",
          4684 => x"ff057789",
          4685 => x"2a065372",
          4686 => x"818a3874",
          4687 => x"527351f3",
          4688 => x"e63f8287",
          4689 => x"cc085382",
          4690 => x"55810b82",
          4691 => x"87cc0827",
          4692 => x"80ff3881",
          4693 => x"558287cc",
          4694 => x"08ff2e80",
          4695 => x"f4389816",
          4696 => x"088287cc",
          4697 => x"082680ca",
          4698 => x"387b8a38",
          4699 => x"7798150c",
          4700 => x"845580dd",
          4701 => x"39941408",
          4702 => x"527351f9",
          4703 => x"863f8287",
          4704 => x"cc085387",
          4705 => x"558287cc",
          4706 => x"08802e80",
          4707 => x"c4388255",
          4708 => x"8287cc08",
          4709 => x"812eba38",
          4710 => x"81558287",
          4711 => x"cc08ff2e",
          4712 => x"b0388287",
          4713 => x"cc085275",
          4714 => x"51fbf33f",
          4715 => x"8287cc08",
          4716 => x"a0387294",
          4717 => x"150c7252",
          4718 => x"7551f2c1",
          4719 => x"3f8287cc",
          4720 => x"0898150c",
          4721 => x"7690150c",
          4722 => x"7716b405",
          4723 => x"9c150c80",
          4724 => x"55748287",
          4725 => x"cc0c8a3d",
          4726 => x"0d04f73d",
          4727 => x"0d7b7d71",
          4728 => x"085b5b57",
          4729 => x"80527651",
          4730 => x"fcac3f82",
          4731 => x"87cc0854",
          4732 => x"8287cc08",
          4733 => x"80ec3882",
          4734 => x"87cc0856",
          4735 => x"98170852",
          4736 => x"7851f083",
          4737 => x"3f8287cc",
          4738 => x"08548287",
          4739 => x"cc0880d2",
          4740 => x"388287cc",
          4741 => x"089c1808",
          4742 => x"70335154",
          4743 => x"587281e5",
          4744 => x"2e098106",
          4745 => x"83388158",
          4746 => x"8287cc08",
          4747 => x"55728338",
          4748 => x"81557775",
          4749 => x"07537280",
          4750 => x"2e8e3881",
          4751 => x"1656757a",
          4752 => x"2e098106",
          4753 => x"8838a539",
          4754 => x"8287cc08",
          4755 => x"56815276",
          4756 => x"51fd8e3f",
          4757 => x"8287cc08",
          4758 => x"548287cc",
          4759 => x"08802eff",
          4760 => x"9b387384",
          4761 => x"2e098106",
          4762 => x"83388754",
          4763 => x"738287cc",
          4764 => x"0c8b3d0d",
          4765 => x"04fd3d0d",
          4766 => x"769a1152",
          4767 => x"54ebec3f",
          4768 => x"8287cc08",
          4769 => x"83ffff06",
          4770 => x"76703351",
          4771 => x"53537183",
          4772 => x"2e098106",
          4773 => x"90389414",
          4774 => x"51ebd03f",
          4775 => x"8287cc08",
          4776 => x"902b7307",
          4777 => x"53728287",
          4778 => x"cc0c853d",
          4779 => x"0d04fc3d",
          4780 => x"0d777970",
          4781 => x"83ffff06",
          4782 => x"549a1253",
          4783 => x"5555ebed",
          4784 => x"3f767033",
          4785 => x"51537283",
          4786 => x"2e098106",
          4787 => x"8b387390",
          4788 => x"2a529415",
          4789 => x"51ebd63f",
          4790 => x"863d0d04",
          4791 => x"f73d0d7b",
          4792 => x"7d5b5584",
          4793 => x"75085a58",
          4794 => x"98150880",
          4795 => x"2e818a38",
          4796 => x"98150852",
          4797 => x"7851ee8f",
          4798 => x"3f8287cc",
          4799 => x"08588287",
          4800 => x"cc0880f5",
          4801 => x"389c1508",
          4802 => x"70335553",
          4803 => x"73863884",
          4804 => x"5880e639",
          4805 => x"8b133370",
          4806 => x"bf067081",
          4807 => x"ff065851",
          4808 => x"53728616",
          4809 => x"348287cc",
          4810 => x"08537381",
          4811 => x"e52e8338",
          4812 => x"815373ae",
          4813 => x"2ea93881",
          4814 => x"70740654",
          4815 => x"5772802e",
          4816 => x"9e38758f",
          4817 => x"2e993882",
          4818 => x"87cc0876",
          4819 => x"df065454",
          4820 => x"72882e09",
          4821 => x"81068338",
          4822 => x"7654737a",
          4823 => x"2ea03880",
          4824 => x"527451fa",
          4825 => x"fc3f8287",
          4826 => x"cc085882",
          4827 => x"87cc0889",
          4828 => x"38981508",
          4829 => x"fefa3886",
          4830 => x"39800b98",
          4831 => x"160c7782",
          4832 => x"87cc0c8b",
          4833 => x"3d0d04fb",
          4834 => x"3d0d7770",
          4835 => x"08575481",
          4836 => x"527351fc",
          4837 => x"c53f8287",
          4838 => x"cc085582",
          4839 => x"87cc08b4",
          4840 => x"38981408",
          4841 => x"527551ec",
          4842 => x"de3f8287",
          4843 => x"cc085582",
          4844 => x"87cc08a0",
          4845 => x"38a05382",
          4846 => x"87cc0852",
          4847 => x"9c140851",
          4848 => x"eadb3f8b",
          4849 => x"53a01452",
          4850 => x"9c140851",
          4851 => x"eaac3f81",
          4852 => x"0b831734",
          4853 => x"748287cc",
          4854 => x"0c873d0d",
          4855 => x"04fd3d0d",
          4856 => x"75700898",
          4857 => x"12085470",
          4858 => x"535553ec",
          4859 => x"9a3f8287",
          4860 => x"cc088d38",
          4861 => x"9c130853",
          4862 => x"e5733481",
          4863 => x"0b831534",
          4864 => x"853d0d04",
          4865 => x"fa3d0d78",
          4866 => x"7a575780",
          4867 => x"0b891734",
          4868 => x"98170880",
          4869 => x"2e818238",
          4870 => x"80708918",
          4871 => x"5555559c",
          4872 => x"17081470",
          4873 => x"33811656",
          4874 => x"515271a0",
          4875 => x"2ea83871",
          4876 => x"852e0981",
          4877 => x"06843881",
          4878 => x"e5527389",
          4879 => x"2e098106",
          4880 => x"8b38ae73",
          4881 => x"70810555",
          4882 => x"34811555",
          4883 => x"71737081",
          4884 => x"05553481",
          4885 => x"15558a74",
          4886 => x"27c53875",
          4887 => x"15880552",
          4888 => x"800b8113",
          4889 => x"349c1708",
          4890 => x"528b1233",
          4891 => x"8817349c",
          4892 => x"17089c11",
          4893 => x"5252e88a",
          4894 => x"3f8287cc",
          4895 => x"08760c96",
          4896 => x"1251e7e7",
          4897 => x"3f8287cc",
          4898 => x"08861723",
          4899 => x"981251e7",
          4900 => x"da3f8287",
          4901 => x"cc088417",
          4902 => x"23883d0d",
          4903 => x"04f33d0d",
          4904 => x"7f70085e",
          4905 => x"5b806170",
          4906 => x"33515555",
          4907 => x"73af2e83",
          4908 => x"38815573",
          4909 => x"80dc2e91",
          4910 => x"3874802e",
          4911 => x"8c38941d",
          4912 => x"08881c0c",
          4913 => x"aa398115",
          4914 => x"41806170",
          4915 => x"33565656",
          4916 => x"73af2e09",
          4917 => x"81068338",
          4918 => x"81567380",
          4919 => x"dc327030",
          4920 => x"70802578",
          4921 => x"07515154",
          4922 => x"73dc3873",
          4923 => x"881c0c60",
          4924 => x"70335154",
          4925 => x"739f2696",
          4926 => x"38ff800b",
          4927 => x"ab1c3480",
          4928 => x"527a51f6",
          4929 => x"913f8287",
          4930 => x"cc085585",
          4931 => x"9839913d",
          4932 => x"61a01d5c",
          4933 => x"5a5e8b53",
          4934 => x"a0527951",
          4935 => x"e7ff3f80",
          4936 => x"70595788",
          4937 => x"7933555c",
          4938 => x"73ae2e09",
          4939 => x"810680d4",
          4940 => x"38781870",
          4941 => x"33811a71",
          4942 => x"ae327030",
          4943 => x"709f2a73",
          4944 => x"82260751",
          4945 => x"51535a57",
          4946 => x"54738c38",
          4947 => x"79175475",
          4948 => x"74348117",
          4949 => x"57db3975",
          4950 => x"af327030",
          4951 => x"709f2a51",
          4952 => x"51547580",
          4953 => x"dc2e8c38",
          4954 => x"73802e87",
          4955 => x"3875a026",
          4956 => x"82bd3877",
          4957 => x"197e0ca4",
          4958 => x"54a07627",
          4959 => x"82bd38a0",
          4960 => x"5482b839",
          4961 => x"78187033",
          4962 => x"811a5a57",
          4963 => x"54a07627",
          4964 => x"81fc3875",
          4965 => x"af327030",
          4966 => x"7780dc32",
          4967 => x"70307280",
          4968 => x"25718025",
          4969 => x"07515156",
          4970 => x"51557380",
          4971 => x"2eac3884",
          4972 => x"39811858",
          4973 => x"80781a70",
          4974 => x"33515555",
          4975 => x"73af2e09",
          4976 => x"81068338",
          4977 => x"81557380",
          4978 => x"dc327030",
          4979 => x"70802577",
          4980 => x"07515154",
          4981 => x"73db3881",
          4982 => x"b53975ae",
          4983 => x"2e098106",
          4984 => x"83388154",
          4985 => x"767c2774",
          4986 => x"07547380",
          4987 => x"2ea2387b",
          4988 => x"8b327030",
          4989 => x"77ae3270",
          4990 => x"30728025",
          4991 => x"719f2a07",
          4992 => x"53515651",
          4993 => x"557481a7",
          4994 => x"3888578b",
          4995 => x"5cfef539",
          4996 => x"75982b54",
          4997 => x"7380258c",
          4998 => x"387580ff",
          4999 => x"06828194",
          5000 => x"11335754",
          5001 => x"7551e6e1",
          5002 => x"3f8287cc",
          5003 => x"08802eb2",
          5004 => x"38781870",
          5005 => x"33811a71",
          5006 => x"545a5654",
          5007 => x"e6d23f82",
          5008 => x"87cc0880",
          5009 => x"2e80e838",
          5010 => x"ff1c5476",
          5011 => x"742780df",
          5012 => x"38791754",
          5013 => x"75743481",
          5014 => x"177a1155",
          5015 => x"57747434",
          5016 => x"a7397552",
          5017 => x"8280b451",
          5018 => x"e5fe3f82",
          5019 => x"87cc08bf",
          5020 => x"38ff9f16",
          5021 => x"54739926",
          5022 => x"8938e016",
          5023 => x"7081ff06",
          5024 => x"57547917",
          5025 => x"54757434",
          5026 => x"811757fd",
          5027 => x"f7397719",
          5028 => x"7e0c7680",
          5029 => x"2e993879",
          5030 => x"33547381",
          5031 => x"e52e0981",
          5032 => x"06843885",
          5033 => x"7a348454",
          5034 => x"a076278f",
          5035 => x"388b3986",
          5036 => x"5581f239",
          5037 => x"845680f3",
          5038 => x"39805473",
          5039 => x"8b1b3480",
          5040 => x"7b085852",
          5041 => x"7a51f2ce",
          5042 => x"3f8287cc",
          5043 => x"08568287",
          5044 => x"cc0880d7",
          5045 => x"38981b08",
          5046 => x"527651e6",
          5047 => x"aa3f8287",
          5048 => x"cc085682",
          5049 => x"87cc0880",
          5050 => x"c2389c1b",
          5051 => x"08703355",
          5052 => x"5573802e",
          5053 => x"ffbe388b",
          5054 => x"1533bf06",
          5055 => x"5473861c",
          5056 => x"348b1533",
          5057 => x"70832a70",
          5058 => x"81065155",
          5059 => x"58739238",
          5060 => x"8b537952",
          5061 => x"7451e49f",
          5062 => x"3f8287cc",
          5063 => x"08802e8b",
          5064 => x"3875527a",
          5065 => x"51f3ba3f",
          5066 => x"ff9f3975",
          5067 => x"ab1c3357",
          5068 => x"5574802e",
          5069 => x"bb387484",
          5070 => x"2e098106",
          5071 => x"80e73875",
          5072 => x"852a7081",
          5073 => x"0677822a",
          5074 => x"58515473",
          5075 => x"802e9638",
          5076 => x"75810654",
          5077 => x"73802efb",
          5078 => x"b538ff80",
          5079 => x"0bab1c34",
          5080 => x"805580c1",
          5081 => x"39758106",
          5082 => x"5473ba38",
          5083 => x"8555b639",
          5084 => x"75822a70",
          5085 => x"81065154",
          5086 => x"73ab3886",
          5087 => x"1b337084",
          5088 => x"2a708106",
          5089 => x"51555573",
          5090 => x"802ee138",
          5091 => x"901b0883",
          5092 => x"ff061db4",
          5093 => x"05527c51",
          5094 => x"f5db3f82",
          5095 => x"87cc0888",
          5096 => x"1c0cfaea",
          5097 => x"39748287",
          5098 => x"cc0c8f3d",
          5099 => x"0d04f63d",
          5100 => x"0d7c5bff",
          5101 => x"7b087071",
          5102 => x"7355595c",
          5103 => x"55597380",
          5104 => x"2e81c638",
          5105 => x"75708105",
          5106 => x"573370a0",
          5107 => x"26525271",
          5108 => x"ba2e8d38",
          5109 => x"70ee3871",
          5110 => x"ba2e0981",
          5111 => x"0681a538",
          5112 => x"7333d011",
          5113 => x"7081ff06",
          5114 => x"51525370",
          5115 => x"89269138",
          5116 => x"82147381",
          5117 => x"ff06d005",
          5118 => x"56527176",
          5119 => x"2e80f738",
          5120 => x"800b8281",
          5121 => x"84595577",
          5122 => x"087a5557",
          5123 => x"76708105",
          5124 => x"58337470",
          5125 => x"81055633",
          5126 => x"ff9f1253",
          5127 => x"53537099",
          5128 => x"268938e0",
          5129 => x"137081ff",
          5130 => x"065451ff",
          5131 => x"9f125170",
          5132 => x"99268938",
          5133 => x"e0127081",
          5134 => x"ff065351",
          5135 => x"7230709f",
          5136 => x"2a515172",
          5137 => x"722e0981",
          5138 => x"06853870",
          5139 => x"ffbe3872",
          5140 => x"30747732",
          5141 => x"70307072",
          5142 => x"079f2a73",
          5143 => x"9f2a0753",
          5144 => x"54545170",
          5145 => x"802e8f38",
          5146 => x"81158419",
          5147 => x"59558375",
          5148 => x"25ff9438",
          5149 => x"8b397483",
          5150 => x"24863874",
          5151 => x"767c0c59",
          5152 => x"78518639",
          5153 => x"829f8433",
          5154 => x"51708287",
          5155 => x"cc0c8c3d",
          5156 => x"0d04fa3d",
          5157 => x"0d785680",
          5158 => x"0b831734",
          5159 => x"ff0bb017",
          5160 => x"0c795275",
          5161 => x"51e2e03f",
          5162 => x"84558287",
          5163 => x"cc088180",
          5164 => x"3884b216",
          5165 => x"51dfb43f",
          5166 => x"8287cc08",
          5167 => x"83ffff06",
          5168 => x"54835573",
          5169 => x"82d4d52e",
          5170 => x"09810680",
          5171 => x"e338800b",
          5172 => x"b4173356",
          5173 => x"577481e9",
          5174 => x"2e098106",
          5175 => x"83388157",
          5176 => x"7481eb32",
          5177 => x"70307080",
          5178 => x"25790751",
          5179 => x"5154738a",
          5180 => x"387481e8",
          5181 => x"2e098106",
          5182 => x"b5388353",
          5183 => x"8280c452",
          5184 => x"80ea1651",
          5185 => x"e0b13f82",
          5186 => x"87cc0855",
          5187 => x"8287cc08",
          5188 => x"802e9d38",
          5189 => x"85538280",
          5190 => x"c8528186",
          5191 => x"1651e097",
          5192 => x"3f8287cc",
          5193 => x"08558287",
          5194 => x"cc08802e",
          5195 => x"83388255",
          5196 => x"748287cc",
          5197 => x"0c883d0d",
          5198 => x"04f23d0d",
          5199 => x"61028405",
          5200 => x"80cb0533",
          5201 => x"58558075",
          5202 => x"0c6051fc",
          5203 => x"e13f8287",
          5204 => x"cc08588b",
          5205 => x"56800b82",
          5206 => x"87cc0824",
          5207 => x"86fb3882",
          5208 => x"87cc0884",
          5209 => x"29829ef0",
          5210 => x"05700855",
          5211 => x"538c5673",
          5212 => x"802e86e5",
          5213 => x"3873750c",
          5214 => x"7681fe06",
          5215 => x"74335457",
          5216 => x"72802eae",
          5217 => x"38811433",
          5218 => x"51d7ca3f",
          5219 => x"8287cc08",
          5220 => x"81ff0670",
          5221 => x"81065455",
          5222 => x"72983876",
          5223 => x"802e86b7",
          5224 => x"3874822a",
          5225 => x"70810651",
          5226 => x"538a5672",
          5227 => x"86ab3886",
          5228 => x"a6398074",
          5229 => x"34778115",
          5230 => x"34815281",
          5231 => x"143351d7",
          5232 => x"b23f8287",
          5233 => x"cc0881ff",
          5234 => x"06708106",
          5235 => x"54558356",
          5236 => x"72868638",
          5237 => x"76802e8f",
          5238 => x"3874822a",
          5239 => x"70810651",
          5240 => x"538a5672",
          5241 => x"85f33880",
          5242 => x"70537452",
          5243 => x"5bfda33f",
          5244 => x"8287cc08",
          5245 => x"81ff0657",
          5246 => x"76822e09",
          5247 => x"810680e2",
          5248 => x"388c3d74",
          5249 => x"56588356",
          5250 => x"83f61533",
          5251 => x"70585372",
          5252 => x"802e8d38",
          5253 => x"83fa1551",
          5254 => x"dce83f82",
          5255 => x"87cc0857",
          5256 => x"76787084",
          5257 => x"055a0cff",
          5258 => x"16901656",
          5259 => x"56758025",
          5260 => x"d738800b",
          5261 => x"8d3d5456",
          5262 => x"72708405",
          5263 => x"54085b83",
          5264 => x"577a802e",
          5265 => x"95387a52",
          5266 => x"7351fcc6",
          5267 => x"3f8287cc",
          5268 => x"0881ff06",
          5269 => x"57817727",
          5270 => x"89388116",
          5271 => x"56837627",
          5272 => x"d7388156",
          5273 => x"76842e84",
          5274 => x"f0388d56",
          5275 => x"76812684",
          5276 => x"e838bf14",
          5277 => x"51dbf43f",
          5278 => x"8287cc08",
          5279 => x"83ffff06",
          5280 => x"53728480",
          5281 => x"2e098106",
          5282 => x"84cf3880",
          5283 => x"ca1451db",
          5284 => x"da3f8287",
          5285 => x"cc0883ff",
          5286 => x"ff065877",
          5287 => x"8d3880d8",
          5288 => x"1451dbde",
          5289 => x"3f8287cc",
          5290 => x"0858779c",
          5291 => x"150c80c4",
          5292 => x"14338215",
          5293 => x"3480c414",
          5294 => x"33ff1170",
          5295 => x"81ff0651",
          5296 => x"54558d56",
          5297 => x"72812684",
          5298 => x"90387481",
          5299 => x"ff067871",
          5300 => x"2980c116",
          5301 => x"33525953",
          5302 => x"728a1523",
          5303 => x"72802e8b",
          5304 => x"38ff1373",
          5305 => x"06537280",
          5306 => x"2e86388d",
          5307 => x"5683ea39",
          5308 => x"80c51451",
          5309 => x"daf53f82",
          5310 => x"87cc0853",
          5311 => x"8287cc08",
          5312 => x"88152372",
          5313 => x"8f06578d",
          5314 => x"567683cd",
          5315 => x"3880c714",
          5316 => x"51dad83f",
          5317 => x"8287cc08",
          5318 => x"83ffff06",
          5319 => x"55748d38",
          5320 => x"80d41451",
          5321 => x"dadc3f82",
          5322 => x"87cc0855",
          5323 => x"80c21451",
          5324 => x"dab93f82",
          5325 => x"87cc0883",
          5326 => x"ffff0653",
          5327 => x"8d567280",
          5328 => x"2e839638",
          5329 => x"88142278",
          5330 => x"1471842a",
          5331 => x"055a5a78",
          5332 => x"75268385",
          5333 => x"388a1422",
          5334 => x"52747931",
          5335 => x"51c58c3f",
          5336 => x"8287cc08",
          5337 => x"558287cc",
          5338 => x"08802e82",
          5339 => x"ec388287",
          5340 => x"cc0880ff",
          5341 => x"fffff526",
          5342 => x"83388357",
          5343 => x"7483fff5",
          5344 => x"26833882",
          5345 => x"57749ff5",
          5346 => x"26853881",
          5347 => x"5789398d",
          5348 => x"5676802e",
          5349 => x"82c33882",
          5350 => x"15709816",
          5351 => x"0c7ba016",
          5352 => x"0c731c70",
          5353 => x"a4170c7a",
          5354 => x"1dac170c",
          5355 => x"54557683",
          5356 => x"2e098106",
          5357 => x"af3880de",
          5358 => x"1451d9af",
          5359 => x"3f8287cc",
          5360 => x"0883ffff",
          5361 => x"06538d56",
          5362 => x"72828e38",
          5363 => x"79828a38",
          5364 => x"80e01451",
          5365 => x"d9ac3f82",
          5366 => x"87cc08a8",
          5367 => x"150c7482",
          5368 => x"2b53a239",
          5369 => x"8d567980",
          5370 => x"2e81ee38",
          5371 => x"7713a815",
          5372 => x"0c741553",
          5373 => x"76822e8d",
          5374 => x"38741015",
          5375 => x"70812a76",
          5376 => x"81060551",
          5377 => x"5383ff13",
          5378 => x"892a538d",
          5379 => x"56729c15",
          5380 => x"082681c5",
          5381 => x"38ff0b90",
          5382 => x"150cff0b",
          5383 => x"8c150cff",
          5384 => x"800b8415",
          5385 => x"3476832e",
          5386 => x"09810681",
          5387 => x"923880e4",
          5388 => x"1451d8b7",
          5389 => x"3f8287cc",
          5390 => x"0883ffff",
          5391 => x"06537281",
          5392 => x"2e098106",
          5393 => x"80f93881",
          5394 => x"1b527351",
          5395 => x"dbb93f82",
          5396 => x"87cc0880",
          5397 => x"ea388287",
          5398 => x"cc088415",
          5399 => x"3484b214",
          5400 => x"51d8883f",
          5401 => x"8287cc08",
          5402 => x"83ffff06",
          5403 => x"537282d4",
          5404 => x"d52e0981",
          5405 => x"0680c838",
          5406 => x"b41451d8",
          5407 => x"853f8287",
          5408 => x"cc08848b",
          5409 => x"85a4d22e",
          5410 => x"098106b3",
          5411 => x"38849814",
          5412 => x"51d7ef3f",
          5413 => x"8287cc08",
          5414 => x"868a85e4",
          5415 => x"f22e0981",
          5416 => x"069d3884",
          5417 => x"9c1451d7",
          5418 => x"d93f8287",
          5419 => x"cc089015",
          5420 => x"0c84a014",
          5421 => x"51d7cb3f",
          5422 => x"8287cc08",
          5423 => x"8c150c76",
          5424 => x"7434829f",
          5425 => x"80228105",
          5426 => x"5372829f",
          5427 => x"80237286",
          5428 => x"1523800b",
          5429 => x"94150c80",
          5430 => x"56758287",
          5431 => x"cc0c903d",
          5432 => x"0d04fb3d",
          5433 => x"0d775489",
          5434 => x"5573802e",
          5435 => x"b9387308",
          5436 => x"5372802e",
          5437 => x"b1387233",
          5438 => x"5271802e",
          5439 => x"a9388613",
          5440 => x"22841522",
          5441 => x"57527176",
          5442 => x"2e098106",
          5443 => x"99388113",
          5444 => x"3351d0c1",
          5445 => x"3f8287cc",
          5446 => x"08810652",
          5447 => x"71883871",
          5448 => x"74085455",
          5449 => x"83398053",
          5450 => x"7873710c",
          5451 => x"52748287",
          5452 => x"cc0c873d",
          5453 => x"0d04fa3d",
          5454 => x"0d02ab05",
          5455 => x"337a5889",
          5456 => x"3dfc0552",
          5457 => x"56f4e73f",
          5458 => x"8b54800b",
          5459 => x"8287cc08",
          5460 => x"24bc3882",
          5461 => x"87cc0884",
          5462 => x"29829ef0",
          5463 => x"05700855",
          5464 => x"5573802e",
          5465 => x"84388074",
          5466 => x"34785473",
          5467 => x"802e8438",
          5468 => x"80743478",
          5469 => x"750c7554",
          5470 => x"75802e92",
          5471 => x"38805389",
          5472 => x"3d705384",
          5473 => x"0551f7b1",
          5474 => x"3f8287cc",
          5475 => x"08547382",
          5476 => x"87cc0c88",
          5477 => x"3d0d04eb",
          5478 => x"3d0d6702",
          5479 => x"840580e7",
          5480 => x"05335959",
          5481 => x"89547880",
          5482 => x"2e84c838",
          5483 => x"77bf0670",
          5484 => x"54983dd0",
          5485 => x"0553993d",
          5486 => x"84055258",
          5487 => x"f6fb3f82",
          5488 => x"87cc0855",
          5489 => x"8287cc08",
          5490 => x"84a4387a",
          5491 => x"5c68528c",
          5492 => x"3d705256",
          5493 => x"edc73f82",
          5494 => x"87cc0855",
          5495 => x"8287cc08",
          5496 => x"92380280",
          5497 => x"d7053370",
          5498 => x"982b5557",
          5499 => x"73802583",
          5500 => x"38865577",
          5501 => x"9c065473",
          5502 => x"802e81ab",
          5503 => x"3874802e",
          5504 => x"95387484",
          5505 => x"2e098106",
          5506 => x"aa387551",
          5507 => x"eaf93f82",
          5508 => x"87cc0855",
          5509 => x"9e3902b2",
          5510 => x"05339106",
          5511 => x"547381b8",
          5512 => x"3877822a",
          5513 => x"70810651",
          5514 => x"5473802e",
          5515 => x"8e388855",
          5516 => x"83bc3977",
          5517 => x"88075874",
          5518 => x"83b43877",
          5519 => x"832a7081",
          5520 => x"06515473",
          5521 => x"802e81af",
          5522 => x"3862527a",
          5523 => x"51e8a63f",
          5524 => x"8287cc08",
          5525 => x"568288b2",
          5526 => x"0a52628e",
          5527 => x"0551d4eb",
          5528 => x"3f6254a0",
          5529 => x"0b8b1534",
          5530 => x"80536252",
          5531 => x"7a51e8be",
          5532 => x"3f805262",
          5533 => x"9c0551d4",
          5534 => x"d23f7a54",
          5535 => x"810b8315",
          5536 => x"3475802e",
          5537 => x"80f1387a",
          5538 => x"b0110851",
          5539 => x"54805375",
          5540 => x"52973dd4",
          5541 => x"0551ddbf",
          5542 => x"3f8287cc",
          5543 => x"08558287",
          5544 => x"cc0882ca",
          5545 => x"38b73974",
          5546 => x"82c43802",
          5547 => x"b2053370",
          5548 => x"842a7081",
          5549 => x"06515556",
          5550 => x"73802e86",
          5551 => x"38845582",
          5552 => x"ad397781",
          5553 => x"2a708106",
          5554 => x"51547380",
          5555 => x"2ea93875",
          5556 => x"81065473",
          5557 => x"802ea038",
          5558 => x"87558292",
          5559 => x"3973527a",
          5560 => x"51d6a43f",
          5561 => x"8287cc08",
          5562 => x"7bff188c",
          5563 => x"120c5555",
          5564 => x"8287cc08",
          5565 => x"81f83877",
          5566 => x"832a7081",
          5567 => x"06515473",
          5568 => x"802e8638",
          5569 => x"7780c007",
          5570 => x"587ab011",
          5571 => x"08a01b0c",
          5572 => x"63a41b0c",
          5573 => x"63537052",
          5574 => x"57e6da3f",
          5575 => x"8287cc08",
          5576 => x"8287cc08",
          5577 => x"881b0c63",
          5578 => x"9c05525a",
          5579 => x"d2d43f82",
          5580 => x"87cc0882",
          5581 => x"87cc088c",
          5582 => x"1b0c777a",
          5583 => x"0c568617",
          5584 => x"22841a23",
          5585 => x"77901a34",
          5586 => x"800b911a",
          5587 => x"34800b9c",
          5588 => x"1a0c800b",
          5589 => x"941a0c77",
          5590 => x"852a7081",
          5591 => x"06515473",
          5592 => x"802e818d",
          5593 => x"388287cc",
          5594 => x"08802e81",
          5595 => x"84388287",
          5596 => x"cc08941a",
          5597 => x"0c8a1722",
          5598 => x"70892b7b",
          5599 => x"525957a8",
          5600 => x"39765278",
          5601 => x"51d7a03f",
          5602 => x"8287cc08",
          5603 => x"578287cc",
          5604 => x"08812683",
          5605 => x"38825582",
          5606 => x"87cc08ff",
          5607 => x"2e098106",
          5608 => x"83387955",
          5609 => x"75783156",
          5610 => x"74307076",
          5611 => x"07802551",
          5612 => x"54777627",
          5613 => x"8a388170",
          5614 => x"7506555a",
          5615 => x"73c33876",
          5616 => x"981a0c74",
          5617 => x"a9387583",
          5618 => x"ff065473",
          5619 => x"802ea238",
          5620 => x"76527a51",
          5621 => x"d6a73f82",
          5622 => x"87cc0885",
          5623 => x"3882558e",
          5624 => x"3975892a",
          5625 => x"8287cc08",
          5626 => x"059c1a0c",
          5627 => x"84398079",
          5628 => x"0c745473",
          5629 => x"8287cc0c",
          5630 => x"973d0d04",
          5631 => x"f23d0d60",
          5632 => x"63656440",
          5633 => x"405d5980",
          5634 => x"7e0c903d",
          5635 => x"fc055278",
          5636 => x"51f9cf3f",
          5637 => x"8287cc08",
          5638 => x"558287cc",
          5639 => x"088a3891",
          5640 => x"19335574",
          5641 => x"802e8638",
          5642 => x"745682c4",
          5643 => x"39901933",
          5644 => x"81065587",
          5645 => x"5674802e",
          5646 => x"82b63895",
          5647 => x"39820b91",
          5648 => x"1a348256",
          5649 => x"82aa3981",
          5650 => x"0b911a34",
          5651 => x"815682a0",
          5652 => x"398c1908",
          5653 => x"941a0831",
          5654 => x"55747c27",
          5655 => x"8338745c",
          5656 => x"7b802e82",
          5657 => x"89389419",
          5658 => x"087083ff",
          5659 => x"06565674",
          5660 => x"81b2387e",
          5661 => x"8a1122ff",
          5662 => x"0577892a",
          5663 => x"065b5579",
          5664 => x"a8387587",
          5665 => x"38881908",
          5666 => x"558f3998",
          5667 => x"19085278",
          5668 => x"51d5943f",
          5669 => x"8287cc08",
          5670 => x"55817527",
          5671 => x"ff9f3874",
          5672 => x"ff2effa3",
          5673 => x"3874981a",
          5674 => x"0c981908",
          5675 => x"527e51d4",
          5676 => x"cc3f8287",
          5677 => x"cc08802e",
          5678 => x"ff833882",
          5679 => x"87cc081a",
          5680 => x"7c892a59",
          5681 => x"5777802e",
          5682 => x"80d63877",
          5683 => x"1a7f8a11",
          5684 => x"22585c55",
          5685 => x"75752785",
          5686 => x"38757a31",
          5687 => x"58775476",
          5688 => x"537c5281",
          5689 => x"1b3351ca",
          5690 => x"893f8287",
          5691 => x"cc08fed7",
          5692 => x"387e8311",
          5693 => x"33565674",
          5694 => x"802e9f38",
          5695 => x"b0160877",
          5696 => x"31557478",
          5697 => x"27943884",
          5698 => x"8053b416",
          5699 => x"52b01608",
          5700 => x"7731892b",
          5701 => x"7d0551cf",
          5702 => x"e13f7789",
          5703 => x"2b56b939",
          5704 => x"769c1a0c",
          5705 => x"94190883",
          5706 => x"ff068480",
          5707 => x"71315755",
          5708 => x"7b762783",
          5709 => x"387b569c",
          5710 => x"1908527e",
          5711 => x"51d1c83f",
          5712 => x"8287cc08",
          5713 => x"fe813875",
          5714 => x"53941908",
          5715 => x"83ff061f",
          5716 => x"b405527c",
          5717 => x"51cfa33f",
          5718 => x"7b76317e",
          5719 => x"08177f0c",
          5720 => x"761e941b",
          5721 => x"0818941c",
          5722 => x"0c5e5cfd",
          5723 => x"f3398056",
          5724 => x"758287cc",
          5725 => x"0c903d0d",
          5726 => x"04f23d0d",
          5727 => x"60636564",
          5728 => x"40405d58",
          5729 => x"807e0c90",
          5730 => x"3dfc0552",
          5731 => x"7751f6d2",
          5732 => x"3f8287cc",
          5733 => x"08558287",
          5734 => x"cc088a38",
          5735 => x"91183355",
          5736 => x"74802e86",
          5737 => x"38745683",
          5738 => x"b8399018",
          5739 => x"3370812a",
          5740 => x"70810651",
          5741 => x"56568756",
          5742 => x"74802e83",
          5743 => x"a4389539",
          5744 => x"820b9119",
          5745 => x"34825683",
          5746 => x"9839810b",
          5747 => x"91193481",
          5748 => x"56838e39",
          5749 => x"9418087c",
          5750 => x"11565674",
          5751 => x"76278438",
          5752 => x"75095c7b",
          5753 => x"802e82ec",
          5754 => x"38941808",
          5755 => x"7083ff06",
          5756 => x"56567481",
          5757 => x"fd387e8a",
          5758 => x"1122ff05",
          5759 => x"77892a06",
          5760 => x"5c557abf",
          5761 => x"38758c38",
          5762 => x"88180855",
          5763 => x"749c387a",
          5764 => x"52853998",
          5765 => x"18085277",
          5766 => x"51d7e83f",
          5767 => x"8287cc08",
          5768 => x"558287cc",
          5769 => x"08802e82",
          5770 => x"ab387481",
          5771 => x"2eff9138",
          5772 => x"74ff2eff",
          5773 => x"95387498",
          5774 => x"190c8818",
          5775 => x"08853874",
          5776 => x"88190c7e",
          5777 => x"55b01508",
          5778 => x"9c19082e",
          5779 => x"0981068d",
          5780 => x"387451ce",
          5781 => x"c23f8287",
          5782 => x"cc08feee",
          5783 => x"38981808",
          5784 => x"527e51d1",
          5785 => x"983f8287",
          5786 => x"cc08802e",
          5787 => x"fed23882",
          5788 => x"87cc081b",
          5789 => x"7c892a5a",
          5790 => x"5778802e",
          5791 => x"80d53878",
          5792 => x"1b7f8a11",
          5793 => x"22585b55",
          5794 => x"75752785",
          5795 => x"38757b31",
          5796 => x"59785476",
          5797 => x"537c5281",
          5798 => x"1a3351c8",
          5799 => x"bf3f8287",
          5800 => x"cc08fea6",
          5801 => x"387eb011",
          5802 => x"08783156",
          5803 => x"56747927",
          5804 => x"9b388480",
          5805 => x"53b01608",
          5806 => x"7731892b",
          5807 => x"7d0552b4",
          5808 => x"1651ccb6",
          5809 => x"3f7e5580",
          5810 => x"0b831634",
          5811 => x"78892b56",
          5812 => x"80db398c",
          5813 => x"18089419",
          5814 => x"08269338",
          5815 => x"7e51cdb7",
          5816 => x"3f8287cc",
          5817 => x"08fde338",
          5818 => x"7e77b012",
          5819 => x"0c55769c",
          5820 => x"190c9418",
          5821 => x"0883ff06",
          5822 => x"84807131",
          5823 => x"57557b76",
          5824 => x"2783387b",
          5825 => x"569c1808",
          5826 => x"527e51cd",
          5827 => x"fa3f8287",
          5828 => x"cc08fdb6",
          5829 => x"3875537c",
          5830 => x"52941808",
          5831 => x"83ff061f",
          5832 => x"b40551cb",
          5833 => x"d53f7e55",
          5834 => x"810b8316",
          5835 => x"347b7631",
          5836 => x"7e08177f",
          5837 => x"0c761e94",
          5838 => x"1a081870",
          5839 => x"941c0c8c",
          5840 => x"1b085858",
          5841 => x"5e5c7476",
          5842 => x"27833875",
          5843 => x"55748c19",
          5844 => x"0cfd9039",
          5845 => x"90183380",
          5846 => x"c0075574",
          5847 => x"90193480",
          5848 => x"56758287",
          5849 => x"cc0c903d",
          5850 => x"0d04f83d",
          5851 => x"0d7a8b3d",
          5852 => x"fc055370",
          5853 => x"5256f2ea",
          5854 => x"3f8287cc",
          5855 => x"08578287",
          5856 => x"cc0880fb",
          5857 => x"38901633",
          5858 => x"70862a70",
          5859 => x"81065155",
          5860 => x"5573802e",
          5861 => x"80e938a0",
          5862 => x"16085278",
          5863 => x"51cce83f",
          5864 => x"8287cc08",
          5865 => x"578287cc",
          5866 => x"0880d438",
          5867 => x"a416088b",
          5868 => x"1133a007",
          5869 => x"5555738b",
          5870 => x"16348816",
          5871 => x"08537452",
          5872 => x"750851dd",
          5873 => x"e93f8c16",
          5874 => x"08529c15",
          5875 => x"51c9fc3f",
          5876 => x"8288b20a",
          5877 => x"52961551",
          5878 => x"c9f13f76",
          5879 => x"52921551",
          5880 => x"c9cb3f78",
          5881 => x"54810b83",
          5882 => x"15347851",
          5883 => x"cce03f82",
          5884 => x"87cc0890",
          5885 => x"173381bf",
          5886 => x"06555773",
          5887 => x"90173476",
          5888 => x"8287cc0c",
          5889 => x"8a3d0d04",
          5890 => x"fc3d0d76",
          5891 => x"705254fe",
          5892 => x"d93f8287",
          5893 => x"cc085382",
          5894 => x"87cc089c",
          5895 => x"38863dfc",
          5896 => x"05527351",
          5897 => x"f1bc3f82",
          5898 => x"87cc0853",
          5899 => x"8287cc08",
          5900 => x"87388287",
          5901 => x"cc08740c",
          5902 => x"728287cc",
          5903 => x"0c863d0d",
          5904 => x"04ff3d0d",
          5905 => x"843d51e6",
          5906 => x"e53f8b52",
          5907 => x"800b8287",
          5908 => x"cc08248b",
          5909 => x"388287cc",
          5910 => x"08829f84",
          5911 => x"34805271",
          5912 => x"8287cc0c",
          5913 => x"833d0d04",
          5914 => x"ef3d0d80",
          5915 => x"53933dd0",
          5916 => x"0552943d",
          5917 => x"51e9c23f",
          5918 => x"8287cc08",
          5919 => x"558287cc",
          5920 => x"0880e038",
          5921 => x"76586352",
          5922 => x"933dd405",
          5923 => x"51e08e3f",
          5924 => x"8287cc08",
          5925 => x"558287cc",
          5926 => x"08bc3802",
          5927 => x"80c70533",
          5928 => x"70982b55",
          5929 => x"56738025",
          5930 => x"8938767a",
          5931 => x"94120c54",
          5932 => x"b23902a2",
          5933 => x"05337084",
          5934 => x"2a708106",
          5935 => x"51555673",
          5936 => x"802e9e38",
          5937 => x"767f5370",
          5938 => x"5254dba9",
          5939 => x"3f8287cc",
          5940 => x"0894150c",
          5941 => x"8e398287",
          5942 => x"cc08842e",
          5943 => x"09810683",
          5944 => x"38855574",
          5945 => x"8287cc0c",
          5946 => x"933d0d04",
          5947 => x"e43d0d6f",
          5948 => x"6f5b5b80",
          5949 => x"7a348053",
          5950 => x"9e3dffb8",
          5951 => x"05529f3d",
          5952 => x"51e8b63f",
          5953 => x"8287cc08",
          5954 => x"578287cc",
          5955 => x"0882fc38",
          5956 => x"7b437a7c",
          5957 => x"94110847",
          5958 => x"55586454",
          5959 => x"73802e81",
          5960 => x"ed38a052",
          5961 => x"933d7052",
          5962 => x"55d5eb3f",
          5963 => x"8287cc08",
          5964 => x"578287cc",
          5965 => x"0882d438",
          5966 => x"68527b51",
          5967 => x"c9c93f82",
          5968 => x"87cc0857",
          5969 => x"8287cc08",
          5970 => x"82c13869",
          5971 => x"527b51da",
          5972 => x"a43f8287",
          5973 => x"cc084576",
          5974 => x"527451d5",
          5975 => x"b93f8287",
          5976 => x"cc085782",
          5977 => x"87cc0882",
          5978 => x"a2388052",
          5979 => x"7451daec",
          5980 => x"3f8287cc",
          5981 => x"08578287",
          5982 => x"cc08a438",
          5983 => x"69527b51",
          5984 => x"d9f33f73",
          5985 => x"8287cc08",
          5986 => x"2ea63876",
          5987 => x"527451d6",
          5988 => x"d03f8287",
          5989 => x"cc085782",
          5990 => x"87cc0880",
          5991 => x"2ecc3876",
          5992 => x"842e0981",
          5993 => x"06863882",
          5994 => x"5781e039",
          5995 => x"7681dc38",
          5996 => x"9e3dffbc",
          5997 => x"05527451",
          5998 => x"dcca3f76",
          5999 => x"903d7811",
          6000 => x"81113351",
          6001 => x"565a5673",
          6002 => x"802e9138",
          6003 => x"02b90555",
          6004 => x"81168116",
          6005 => x"70335656",
          6006 => x"5673f538",
          6007 => x"81165473",
          6008 => x"78268190",
          6009 => x"3875802e",
          6010 => x"99387816",
          6011 => x"810555ff",
          6012 => x"186f11ff",
          6013 => x"18ff1858",
          6014 => x"58555874",
          6015 => x"33743475",
          6016 => x"ee38ff18",
          6017 => x"6f115558",
          6018 => x"af7434fe",
          6019 => x"8d39777b",
          6020 => x"2e098106",
          6021 => x"8a38ff18",
          6022 => x"6f115558",
          6023 => x"af743480",
          6024 => x"0b829f84",
          6025 => x"33708429",
          6026 => x"82818405",
          6027 => x"70087033",
          6028 => x"525c5656",
          6029 => x"5673762e",
          6030 => x"8d388116",
          6031 => x"701a7033",
          6032 => x"51555673",
          6033 => x"f5388216",
          6034 => x"54737826",
          6035 => x"a7388055",
          6036 => x"74762791",
          6037 => x"38741954",
          6038 => x"73337a70",
          6039 => x"81055c34",
          6040 => x"811555ec",
          6041 => x"39ba7a70",
          6042 => x"81055c34",
          6043 => x"74ff2e09",
          6044 => x"81068538",
          6045 => x"91579439",
          6046 => x"6e188119",
          6047 => x"59547333",
          6048 => x"7a708105",
          6049 => x"5c347a78",
          6050 => x"26ee3880",
          6051 => x"7a347682",
          6052 => x"87cc0c9e",
          6053 => x"3d0d04f7",
          6054 => x"3d0d7b7d",
          6055 => x"8d3dfc05",
          6056 => x"54715357",
          6057 => x"55ecbb3f",
          6058 => x"8287cc08",
          6059 => x"538287cc",
          6060 => x"0882fa38",
          6061 => x"91153353",
          6062 => x"7282f238",
          6063 => x"8c150854",
          6064 => x"73762792",
          6065 => x"38901533",
          6066 => x"70812a70",
          6067 => x"81065154",
          6068 => x"57728338",
          6069 => x"73569415",
          6070 => x"08548070",
          6071 => x"94170c58",
          6072 => x"75782e82",
          6073 => x"9738798a",
          6074 => x"11227089",
          6075 => x"2b595153",
          6076 => x"73782eb7",
          6077 => x"387652ff",
          6078 => x"1651ffad",
          6079 => x"ee3f8287",
          6080 => x"cc08ff15",
          6081 => x"78547053",
          6082 => x"5553ffad",
          6083 => x"de3f8287",
          6084 => x"cc087326",
          6085 => x"96387630",
          6086 => x"70750670",
          6087 => x"94180c77",
          6088 => x"71319818",
          6089 => x"08575851",
          6090 => x"53b13988",
          6091 => x"15085473",
          6092 => x"a6387352",
          6093 => x"7451cdcb",
          6094 => x"3f8287cc",
          6095 => x"08548287",
          6096 => x"cc08812e",
          6097 => x"819a3882",
          6098 => x"87cc08ff",
          6099 => x"2e819b38",
          6100 => x"8287cc08",
          6101 => x"88160c73",
          6102 => x"98160c73",
          6103 => x"802e819c",
          6104 => x"38767627",
          6105 => x"80dc3875",
          6106 => x"77319416",
          6107 => x"08189417",
          6108 => x"0c901633",
          6109 => x"70812a70",
          6110 => x"81065155",
          6111 => x"5a567280",
          6112 => x"2e9a3873",
          6113 => x"527451cc",
          6114 => x"fa3f8287",
          6115 => x"cc085482",
          6116 => x"87cc0894",
          6117 => x"388287cc",
          6118 => x"0856a739",
          6119 => x"73527451",
          6120 => x"c7853f82",
          6121 => x"87cc0854",
          6122 => x"73ff2ebe",
          6123 => x"38817427",
          6124 => x"af387953",
          6125 => x"73981408",
          6126 => x"27a63873",
          6127 => x"98160cff",
          6128 => x"a0399415",
          6129 => x"08169416",
          6130 => x"0c7583ff",
          6131 => x"06537280",
          6132 => x"2eaa3873",
          6133 => x"527951c6",
          6134 => x"a43f8287",
          6135 => x"cc089438",
          6136 => x"820b9116",
          6137 => x"34825380",
          6138 => x"c439810b",
          6139 => x"91163481",
          6140 => x"53bb3975",
          6141 => x"892a8287",
          6142 => x"cc080558",
          6143 => x"94150854",
          6144 => x"8c150874",
          6145 => x"27903873",
          6146 => x"8c160c90",
          6147 => x"153380c0",
          6148 => x"07537290",
          6149 => x"16347383",
          6150 => x"ff065372",
          6151 => x"802e8c38",
          6152 => x"779c1608",
          6153 => x"2e853877",
          6154 => x"9c160c80",
          6155 => x"53728287",
          6156 => x"cc0c8b3d",
          6157 => x"0d04f93d",
          6158 => x"0d795689",
          6159 => x"5475802e",
          6160 => x"818a3880",
          6161 => x"53893dfc",
          6162 => x"05528a3d",
          6163 => x"840551e1",
          6164 => x"e83f8287",
          6165 => x"cc085582",
          6166 => x"87cc0880",
          6167 => x"ea387776",
          6168 => x"0c7a5275",
          6169 => x"51d8b63f",
          6170 => x"8287cc08",
          6171 => x"558287cc",
          6172 => x"0880c338",
          6173 => x"ab163370",
          6174 => x"982b5557",
          6175 => x"807424a2",
          6176 => x"38861633",
          6177 => x"70842a70",
          6178 => x"81065155",
          6179 => x"5773802e",
          6180 => x"ad389c16",
          6181 => x"08527751",
          6182 => x"d3db3f82",
          6183 => x"87cc0888",
          6184 => x"170c7754",
          6185 => x"86142284",
          6186 => x"17237452",
          6187 => x"7551cee6",
          6188 => x"3f8287cc",
          6189 => x"08557484",
          6190 => x"2e098106",
          6191 => x"85388555",
          6192 => x"86397480",
          6193 => x"2e843880",
          6194 => x"760c7454",
          6195 => x"738287cc",
          6196 => x"0c893d0d",
          6197 => x"04fc3d0d",
          6198 => x"76873dfc",
          6199 => x"05537052",
          6200 => x"53e7ff3f",
          6201 => x"8287cc08",
          6202 => x"87388287",
          6203 => x"cc08730c",
          6204 => x"863d0d04",
          6205 => x"fb3d0d77",
          6206 => x"79893dfc",
          6207 => x"05547153",
          6208 => x"5654e7de",
          6209 => x"3f8287cc",
          6210 => x"08538287",
          6211 => x"cc0880df",
          6212 => x"38749338",
          6213 => x"8287cc08",
          6214 => x"527351cd",
          6215 => x"f93f8287",
          6216 => x"cc085380",
          6217 => x"ca398287",
          6218 => x"cc085273",
          6219 => x"51d3ad3f",
          6220 => x"8287cc08",
          6221 => x"538287cc",
          6222 => x"08842e09",
          6223 => x"81068538",
          6224 => x"80538739",
          6225 => x"8287cc08",
          6226 => x"a6387452",
          6227 => x"7351d5b4",
          6228 => x"3f725273",
          6229 => x"51cf8a3f",
          6230 => x"8287cc08",
          6231 => x"84327030",
          6232 => x"7072079f",
          6233 => x"2c708287",
          6234 => x"cc080651",
          6235 => x"51545472",
          6236 => x"8287cc0c",
          6237 => x"873d0d04",
          6238 => x"ee3d0d65",
          6239 => x"57805389",
          6240 => x"3d705396",
          6241 => x"3d5256df",
          6242 => x"b03f8287",
          6243 => x"cc085582",
          6244 => x"87cc08b2",
          6245 => x"38645275",
          6246 => x"51d6823f",
          6247 => x"8287cc08",
          6248 => x"558287cc",
          6249 => x"08a03802",
          6250 => x"80cb0533",
          6251 => x"70982b55",
          6252 => x"58738025",
          6253 => x"85388655",
          6254 => x"8d397680",
          6255 => x"2e883876",
          6256 => x"527551d4",
          6257 => x"bf3f7482",
          6258 => x"87cc0c94",
          6259 => x"3d0d04f0",
          6260 => x"3d0d6365",
          6261 => x"555c8053",
          6262 => x"923dec05",
          6263 => x"52933d51",
          6264 => x"ded73f82",
          6265 => x"87cc085b",
          6266 => x"8287cc08",
          6267 => x"8280387c",
          6268 => x"740c7308",
          6269 => x"981108fe",
          6270 => x"11901308",
          6271 => x"59565855",
          6272 => x"75742691",
          6273 => x"38757c0c",
          6274 => x"81e43981",
          6275 => x"5b81cc39",
          6276 => x"825b81c7",
          6277 => x"398287cc",
          6278 => x"08753355",
          6279 => x"5973812e",
          6280 => x"098106bf",
          6281 => x"3882755f",
          6282 => x"57765292",
          6283 => x"3df00551",
          6284 => x"c1f53f82",
          6285 => x"87cc08ff",
          6286 => x"2ed13882",
          6287 => x"87cc0881",
          6288 => x"2ece3882",
          6289 => x"87cc0830",
          6290 => x"708287cc",
          6291 => x"08078025",
          6292 => x"7a058119",
          6293 => x"7f53595a",
          6294 => x"54981408",
          6295 => x"7726ca38",
          6296 => x"80f939a4",
          6297 => x"15088287",
          6298 => x"cc085758",
          6299 => x"75983877",
          6300 => x"5281187d",
          6301 => x"5258ffbf",
          6302 => x"8e3f8287",
          6303 => x"cc085b82",
          6304 => x"87cc0880",
          6305 => x"d6387c70",
          6306 => x"337712ff",
          6307 => x"1a5d5256",
          6308 => x"5474822e",
          6309 => x"0981069e",
          6310 => x"38b41451",
          6311 => x"ffbbcc3f",
          6312 => x"8287cc08",
          6313 => x"83ffff06",
          6314 => x"70307080",
          6315 => x"251b8219",
          6316 => x"595b5154",
          6317 => x"9b39b414",
          6318 => x"51ffbbc6",
          6319 => x"3f8287cc",
          6320 => x"08f00a06",
          6321 => x"70307080",
          6322 => x"251b8419",
          6323 => x"595b5154",
          6324 => x"7583ff06",
          6325 => x"7a585679",
          6326 => x"ff923878",
          6327 => x"7c0c7c79",
          6328 => x"90120c84",
          6329 => x"11338107",
          6330 => x"56547484",
          6331 => x"15347a82",
          6332 => x"87cc0c92",
          6333 => x"3d0d04f9",
          6334 => x"3d0d798a",
          6335 => x"3dfc0553",
          6336 => x"705257e3",
          6337 => x"dd3f8287",
          6338 => x"cc085682",
          6339 => x"87cc0881",
          6340 => x"a8389117",
          6341 => x"33567581",
          6342 => x"a0389017",
          6343 => x"3370812a",
          6344 => x"70810651",
          6345 => x"55558755",
          6346 => x"73802e81",
          6347 => x"8e389417",
          6348 => x"0854738c",
          6349 => x"18082781",
          6350 => x"8038739b",
          6351 => x"388287cc",
          6352 => x"08538817",
          6353 => x"08527651",
          6354 => x"c48d3f82",
          6355 => x"87cc0874",
          6356 => x"88190c56",
          6357 => x"80c93998",
          6358 => x"17085276",
          6359 => x"51ffbfc7",
          6360 => x"3f8287cc",
          6361 => x"08ff2e09",
          6362 => x"81068338",
          6363 => x"81568287",
          6364 => x"cc08812e",
          6365 => x"09810685",
          6366 => x"388256a3",
          6367 => x"3975a038",
          6368 => x"77548287",
          6369 => x"cc089815",
          6370 => x"08279438",
          6371 => x"98170853",
          6372 => x"8287cc08",
          6373 => x"527651c3",
          6374 => x"be3f8287",
          6375 => x"cc085694",
          6376 => x"17088c18",
          6377 => x"0c901733",
          6378 => x"80c00754",
          6379 => x"73901834",
          6380 => x"75802e85",
          6381 => x"38759118",
          6382 => x"34755574",
          6383 => x"8287cc0c",
          6384 => x"893d0d04",
          6385 => x"e23d0d82",
          6386 => x"53a03dff",
          6387 => x"a40552a1",
          6388 => x"3d51dae5",
          6389 => x"3f8287cc",
          6390 => x"08558287",
          6391 => x"cc0881f5",
          6392 => x"387845a1",
          6393 => x"3d085295",
          6394 => x"3d705258",
          6395 => x"d1af3f82",
          6396 => x"87cc0855",
          6397 => x"8287cc08",
          6398 => x"81db3802",
          6399 => x"80fb0533",
          6400 => x"70852a70",
          6401 => x"81065155",
          6402 => x"56865573",
          6403 => x"81c73875",
          6404 => x"982b5480",
          6405 => x"742481bd",
          6406 => x"380280d6",
          6407 => x"05337081",
          6408 => x"06585487",
          6409 => x"557681ad",
          6410 => x"386b5278",
          6411 => x"51ccc63f",
          6412 => x"8287cc08",
          6413 => x"74842a70",
          6414 => x"81065155",
          6415 => x"5673802e",
          6416 => x"80d43878",
          6417 => x"548287cc",
          6418 => x"08941508",
          6419 => x"2e818638",
          6420 => x"735a8287",
          6421 => x"cc085c76",
          6422 => x"528a3d70",
          6423 => x"5254c7b6",
          6424 => x"3f8287cc",
          6425 => x"08558287",
          6426 => x"cc0880e9",
          6427 => x"388287cc",
          6428 => x"08527351",
          6429 => x"cce63f82",
          6430 => x"87cc0855",
          6431 => x"8287cc08",
          6432 => x"86388755",
          6433 => x"80cf3982",
          6434 => x"87cc0884",
          6435 => x"2e883882",
          6436 => x"87cc0880",
          6437 => x"c0387751",
          6438 => x"cec33f82",
          6439 => x"87cc0882",
          6440 => x"87cc0830",
          6441 => x"708287cc",
          6442 => x"08078025",
          6443 => x"51555575",
          6444 => x"802e9438",
          6445 => x"73802e8f",
          6446 => x"38805375",
          6447 => x"527751c1",
          6448 => x"963f8287",
          6449 => x"cc085574",
          6450 => x"8c387851",
          6451 => x"ffbaff3f",
          6452 => x"8287cc08",
          6453 => x"55748287",
          6454 => x"cc0ca03d",
          6455 => x"0d04e93d",
          6456 => x"0d825399",
          6457 => x"3dc00552",
          6458 => x"9a3d51d8",
          6459 => x"cc3f8287",
          6460 => x"cc085482",
          6461 => x"87cc0882",
          6462 => x"b038785e",
          6463 => x"69528e3d",
          6464 => x"705258cf",
          6465 => x"983f8287",
          6466 => x"cc085482",
          6467 => x"87cc0886",
          6468 => x"38885482",
          6469 => x"94398287",
          6470 => x"cc08842e",
          6471 => x"09810682",
          6472 => x"88380280",
          6473 => x"df053370",
          6474 => x"852a8106",
          6475 => x"51558654",
          6476 => x"7481f638",
          6477 => x"785a7452",
          6478 => x"8a3d7052",
          6479 => x"57c1c43f",
          6480 => x"8287cc08",
          6481 => x"75555682",
          6482 => x"87cc0883",
          6483 => x"38875482",
          6484 => x"87cc0881",
          6485 => x"2e098106",
          6486 => x"83388254",
          6487 => x"8287cc08",
          6488 => x"ff2e0981",
          6489 => x"06863881",
          6490 => x"5481b439",
          6491 => x"7381b038",
          6492 => x"8287cc08",
          6493 => x"527851c4",
          6494 => x"a53f8287",
          6495 => x"cc085482",
          6496 => x"87cc0881",
          6497 => x"9a388b53",
          6498 => x"a052b419",
          6499 => x"51ffb78d",
          6500 => x"3f7854ae",
          6501 => x"0bb41534",
          6502 => x"7854900b",
          6503 => x"bf153482",
          6504 => x"88b20a52",
          6505 => x"80ca1951",
          6506 => x"ffb6a03f",
          6507 => x"755378b4",
          6508 => x"115351c9",
          6509 => x"f93fa053",
          6510 => x"78b41153",
          6511 => x"80d40551",
          6512 => x"ffb6b73f",
          6513 => x"7854ae0b",
          6514 => x"80d51534",
          6515 => x"7f537880",
          6516 => x"d4115351",
          6517 => x"c9d83f78",
          6518 => x"54810b83",
          6519 => x"15347751",
          6520 => x"cba53f82",
          6521 => x"87cc0854",
          6522 => x"8287cc08",
          6523 => x"b2388288",
          6524 => x"b20a5264",
          6525 => x"960551ff",
          6526 => x"b5d13f75",
          6527 => x"53645278",
          6528 => x"51c9ab3f",
          6529 => x"6454900b",
          6530 => x"8b153478",
          6531 => x"54810b83",
          6532 => x"15347851",
          6533 => x"ffb8b73f",
          6534 => x"8287cc08",
          6535 => x"548b3980",
          6536 => x"53755276",
          6537 => x"51ffbeaf",
          6538 => x"3f738287",
          6539 => x"cc0c993d",
          6540 => x"0d04da3d",
          6541 => x"0da93d84",
          6542 => x"0551d2f2",
          6543 => x"3f8253a8",
          6544 => x"3dff8405",
          6545 => x"52a93d51",
          6546 => x"d5ef3f82",
          6547 => x"87cc0855",
          6548 => x"8287cc08",
          6549 => x"82d33878",
          6550 => x"4da93d08",
          6551 => x"529d3d70",
          6552 => x"5258ccb9",
          6553 => x"3f8287cc",
          6554 => x"08558287",
          6555 => x"cc0882b9",
          6556 => x"3802819b",
          6557 => x"053381a0",
          6558 => x"06548655",
          6559 => x"7382aa38",
          6560 => x"a053a43d",
          6561 => x"0852a83d",
          6562 => x"ff880551",
          6563 => x"ffb4eb3f",
          6564 => x"ac537752",
          6565 => x"923d7052",
          6566 => x"54ffb4de",
          6567 => x"3faa3d08",
          6568 => x"527351cb",
          6569 => x"f83f8287",
          6570 => x"cc085582",
          6571 => x"87cc0895",
          6572 => x"38636f2e",
          6573 => x"09810688",
          6574 => x"3865a23d",
          6575 => x"082e9238",
          6576 => x"885581e5",
          6577 => x"398287cc",
          6578 => x"08842e09",
          6579 => x"810681b8",
          6580 => x"387351c9",
          6581 => x"b23f8287",
          6582 => x"cc085582",
          6583 => x"87cc0881",
          6584 => x"c8386856",
          6585 => x"9353a83d",
          6586 => x"ff950552",
          6587 => x"8d1651ff",
          6588 => x"b4883f02",
          6589 => x"af05338b",
          6590 => x"17348b16",
          6591 => x"3370842a",
          6592 => x"70810651",
          6593 => x"55557389",
          6594 => x"3874a007",
          6595 => x"54738b17",
          6596 => x"34785481",
          6597 => x"0b831534",
          6598 => x"8b163370",
          6599 => x"842a7081",
          6600 => x"06515555",
          6601 => x"73802e80",
          6602 => x"e5386e64",
          6603 => x"2e80df38",
          6604 => x"75527851",
          6605 => x"c6bf3f82",
          6606 => x"87cc0852",
          6607 => x"7851ffb7",
          6608 => x"bc3f8255",
          6609 => x"8287cc08",
          6610 => x"802e80dd",
          6611 => x"388287cc",
          6612 => x"08527851",
          6613 => x"ffb5b03f",
          6614 => x"8287cc08",
          6615 => x"7980d411",
          6616 => x"58585582",
          6617 => x"87cc0880",
          6618 => x"c0388116",
          6619 => x"335473ae",
          6620 => x"2e098106",
          6621 => x"99386353",
          6622 => x"75527651",
          6623 => x"c6b03f78",
          6624 => x"54810b83",
          6625 => x"15348739",
          6626 => x"8287cc08",
          6627 => x"9c387751",
          6628 => x"c8cb3f82",
          6629 => x"87cc0855",
          6630 => x"8287cc08",
          6631 => x"8c387851",
          6632 => x"ffb5ab3f",
          6633 => x"8287cc08",
          6634 => x"55748287",
          6635 => x"cc0ca83d",
          6636 => x"0d04ed3d",
          6637 => x"0d0280db",
          6638 => x"05330284",
          6639 => x"0580df05",
          6640 => x"33575782",
          6641 => x"53953dd0",
          6642 => x"0552963d",
          6643 => x"51d2ea3f",
          6644 => x"8287cc08",
          6645 => x"558287cc",
          6646 => x"0880cf38",
          6647 => x"785a6552",
          6648 => x"953dd405",
          6649 => x"51c9b63f",
          6650 => x"8287cc08",
          6651 => x"558287cc",
          6652 => x"08b83802",
          6653 => x"80cf0533",
          6654 => x"81a00654",
          6655 => x"865573aa",
          6656 => x"3875a706",
          6657 => x"6171098b",
          6658 => x"12337106",
          6659 => x"7a740607",
          6660 => x"51575556",
          6661 => x"748b1534",
          6662 => x"7854810b",
          6663 => x"83153478",
          6664 => x"51ffb4aa",
          6665 => x"3f8287cc",
          6666 => x"08557482",
          6667 => x"87cc0c95",
          6668 => x"3d0d04ef",
          6669 => x"3d0d6456",
          6670 => x"8253933d",
          6671 => x"d0055294",
          6672 => x"3d51d1f5",
          6673 => x"3f8287cc",
          6674 => x"08558287",
          6675 => x"cc0880cb",
          6676 => x"38765863",
          6677 => x"52933dd4",
          6678 => x"0551c8c1",
          6679 => x"3f8287cc",
          6680 => x"08558287",
          6681 => x"cc08b438",
          6682 => x"0280c705",
          6683 => x"3381a006",
          6684 => x"54865573",
          6685 => x"a6388416",
          6686 => x"22861722",
          6687 => x"71902b07",
          6688 => x"5354961f",
          6689 => x"51ffb0c3",
          6690 => x"3f765481",
          6691 => x"0b831534",
          6692 => x"7651ffb3",
          6693 => x"b93f8287",
          6694 => x"cc085574",
          6695 => x"8287cc0c",
          6696 => x"933d0d04",
          6697 => x"ea3d0d69",
          6698 => x"6b5c5a80",
          6699 => x"53983dd0",
          6700 => x"0552993d",
          6701 => x"51d1823f",
          6702 => x"8287cc08",
          6703 => x"8287cc08",
          6704 => x"30708287",
          6705 => x"cc080780",
          6706 => x"25515557",
          6707 => x"79802e81",
          6708 => x"85388170",
          6709 => x"75065555",
          6710 => x"73802e80",
          6711 => x"f9387b5d",
          6712 => x"805f8052",
          6713 => x"8d3d7052",
          6714 => x"54ffbeaa",
          6715 => x"3f8287cc",
          6716 => x"08578287",
          6717 => x"cc0880d1",
          6718 => x"38745273",
          6719 => x"51c3dd3f",
          6720 => x"8287cc08",
          6721 => x"578287cc",
          6722 => x"08bf3882",
          6723 => x"87cc0882",
          6724 => x"87cc0865",
          6725 => x"5b595678",
          6726 => x"1881197b",
          6727 => x"18565955",
          6728 => x"74337434",
          6729 => x"8116568a",
          6730 => x"7827ec38",
          6731 => x"8b56751a",
          6732 => x"54807434",
          6733 => x"75802e9e",
          6734 => x"38ff1670",
          6735 => x"1b703351",
          6736 => x"555673a0",
          6737 => x"2ee8388e",
          6738 => x"3976842e",
          6739 => x"09810686",
          6740 => x"38807a34",
          6741 => x"80577630",
          6742 => x"70780780",
          6743 => x"2551547a",
          6744 => x"802e80c1",
          6745 => x"3873802e",
          6746 => x"bc387ba0",
          6747 => x"11085351",
          6748 => x"ffb1943f",
          6749 => x"8287cc08",
          6750 => x"578287cc",
          6751 => x"08a7387b",
          6752 => x"70335555",
          6753 => x"80c35673",
          6754 => x"832e8b38",
          6755 => x"80e45673",
          6756 => x"842e8338",
          6757 => x"a7567515",
          6758 => x"b40551ff",
          6759 => x"ade43f82",
          6760 => x"87cc087b",
          6761 => x"0c768287",
          6762 => x"cc0c983d",
          6763 => x"0d04e63d",
          6764 => x"0d82539c",
          6765 => x"3dffb805",
          6766 => x"529d3d51",
          6767 => x"cefb3f82",
          6768 => x"87cc0882",
          6769 => x"87cc0856",
          6770 => x"548287cc",
          6771 => x"08839838",
          6772 => x"8b53a052",
          6773 => x"8b3d7052",
          6774 => x"59ffaec1",
          6775 => x"3f736d70",
          6776 => x"337081ff",
          6777 => x"06525755",
          6778 => x"579f7427",
          6779 => x"81bc3878",
          6780 => x"587481ff",
          6781 => x"066d8105",
          6782 => x"4e705255",
          6783 => x"ffaf8a3f",
          6784 => x"8287cc08",
          6785 => x"802ea538",
          6786 => x"6c703370",
          6787 => x"535754ff",
          6788 => x"aefe3f82",
          6789 => x"87cc0880",
          6790 => x"2e8d3874",
          6791 => x"882b7607",
          6792 => x"6d81054e",
          6793 => x"55863982",
          6794 => x"87cc0855",
          6795 => x"ff9f1570",
          6796 => x"83ffff06",
          6797 => x"51547399",
          6798 => x"268a38e0",
          6799 => x"157083ff",
          6800 => x"ff065654",
          6801 => x"80ff7527",
          6802 => x"87388280",
          6803 => x"94153355",
          6804 => x"74802ea3",
          6805 => x"38745282",
          6806 => x"829451ff",
          6807 => x"ae8a3f82",
          6808 => x"87cc0893",
          6809 => x"3881ff75",
          6810 => x"27883876",
          6811 => x"89268838",
          6812 => x"8b398a77",
          6813 => x"27863886",
          6814 => x"5581ec39",
          6815 => x"81ff7527",
          6816 => x"8f387488",
          6817 => x"2a547378",
          6818 => x"7081055a",
          6819 => x"34811757",
          6820 => x"74787081",
          6821 => x"055a3481",
          6822 => x"176d7033",
          6823 => x"7081ff06",
          6824 => x"52575557",
          6825 => x"739f26fe",
          6826 => x"c8388b3d",
          6827 => x"33548655",
          6828 => x"7381e52e",
          6829 => x"81b13876",
          6830 => x"802e9938",
          6831 => x"02a70555",
          6832 => x"76157033",
          6833 => x"515473a0",
          6834 => x"2e098106",
          6835 => x"8738ff17",
          6836 => x"5776ed38",
          6837 => x"79418043",
          6838 => x"8052913d",
          6839 => x"705255ff",
          6840 => x"bab43f82",
          6841 => x"87cc0854",
          6842 => x"8287cc08",
          6843 => x"80f73881",
          6844 => x"527451ff",
          6845 => x"bfe63f82",
          6846 => x"87cc0854",
          6847 => x"8287cc08",
          6848 => x"8d387680",
          6849 => x"c4386754",
          6850 => x"e5743480",
          6851 => x"c6398287",
          6852 => x"cc08842e",
          6853 => x"09810680",
          6854 => x"cc388054",
          6855 => x"76742e80",
          6856 => x"c4388152",
          6857 => x"7451ffbd",
          6858 => x"b13f8287",
          6859 => x"cc085482",
          6860 => x"87cc08b1",
          6861 => x"38a05382",
          6862 => x"87cc0852",
          6863 => x"6751ffab",
          6864 => x"dc3f6754",
          6865 => x"880b8b15",
          6866 => x"348b5378",
          6867 => x"526751ff",
          6868 => x"aba83f79",
          6869 => x"54810b83",
          6870 => x"15347951",
          6871 => x"ffadef3f",
          6872 => x"8287cc08",
          6873 => x"54735574",
          6874 => x"8287cc0c",
          6875 => x"9c3d0d04",
          6876 => x"f23d0d60",
          6877 => x"62028805",
          6878 => x"80cb0533",
          6879 => x"933dfc05",
          6880 => x"55725440",
          6881 => x"5e5ad2da",
          6882 => x"3f8287cc",
          6883 => x"08588287",
          6884 => x"cc0882bd",
          6885 => x"38911a33",
          6886 => x"587782b5",
          6887 => x"387c802e",
          6888 => x"97388c1a",
          6889 => x"08597890",
          6890 => x"38901a33",
          6891 => x"70812a70",
          6892 => x"81065155",
          6893 => x"55739038",
          6894 => x"87548297",
          6895 => x"39825882",
          6896 => x"90398158",
          6897 => x"828b397e",
          6898 => x"8a112270",
          6899 => x"892b7055",
          6900 => x"7f545656",
          6901 => x"56ff9493",
          6902 => x"3fff147d",
          6903 => x"06703070",
          6904 => x"72079f2a",
          6905 => x"8287cc08",
          6906 => x"058c1908",
          6907 => x"7c405a5d",
          6908 => x"55558177",
          6909 => x"27883898",
          6910 => x"16087726",
          6911 => x"83388257",
          6912 => x"76775659",
          6913 => x"80567452",
          6914 => x"7951ffae",
          6915 => x"9a3f8115",
          6916 => x"7f555598",
          6917 => x"14087526",
          6918 => x"83388255",
          6919 => x"8287cc08",
          6920 => x"812eff99",
          6921 => x"388287cc",
          6922 => x"08ff2eff",
          6923 => x"95388287",
          6924 => x"cc088e38",
          6925 => x"81165675",
          6926 => x"7b2e0981",
          6927 => x"06873893",
          6928 => x"39745980",
          6929 => x"5674772e",
          6930 => x"098106ff",
          6931 => x"b9388758",
          6932 => x"80ff397d",
          6933 => x"802eba38",
          6934 => x"787b5555",
          6935 => x"7a802eb4",
          6936 => x"38811556",
          6937 => x"73812e09",
          6938 => x"81068338",
          6939 => x"ff567553",
          6940 => x"74527e51",
          6941 => x"ffafa93f",
          6942 => x"8287cc08",
          6943 => x"588287cc",
          6944 => x"0880ce38",
          6945 => x"748116ff",
          6946 => x"1656565c",
          6947 => x"73d33884",
          6948 => x"39ff195c",
          6949 => x"7e7c8c12",
          6950 => x"0c557d80",
          6951 => x"2eb33878",
          6952 => x"881b0c7c",
          6953 => x"8c1b0c90",
          6954 => x"1a3380c0",
          6955 => x"07547390",
          6956 => x"1b349815",
          6957 => x"08fe0590",
          6958 => x"16085754",
          6959 => x"75742691",
          6960 => x"38757b31",
          6961 => x"90160c84",
          6962 => x"15338107",
          6963 => x"54738416",
          6964 => x"34775473",
          6965 => x"8287cc0c",
          6966 => x"903d0d04",
          6967 => x"e93d0d6b",
          6968 => x"6d028805",
          6969 => x"80eb0533",
          6970 => x"9d3d545a",
          6971 => x"5c59c5be",
          6972 => x"3f8b5680",
          6973 => x"0b8287cc",
          6974 => x"08248bf8",
          6975 => x"388287cc",
          6976 => x"08842982",
          6977 => x"9ef00570",
          6978 => x"08515574",
          6979 => x"802e8438",
          6980 => x"80753482",
          6981 => x"87cc0881",
          6982 => x"ff065f81",
          6983 => x"527e51ff",
          6984 => x"a0d13f82",
          6985 => x"87cc0881",
          6986 => x"ff067081",
          6987 => x"06565783",
          6988 => x"56748bc0",
          6989 => x"3876822a",
          6990 => x"70810651",
          6991 => x"558a5674",
          6992 => x"8bb23899",
          6993 => x"3dfc0553",
          6994 => x"83527e51",
          6995 => x"ffa4f13f",
          6996 => x"8287cc08",
          6997 => x"99386755",
          6998 => x"74802e92",
          6999 => x"38748280",
          7000 => x"80268b38",
          7001 => x"ff157506",
          7002 => x"5574802e",
          7003 => x"83388148",
          7004 => x"78802e87",
          7005 => x"38848079",
          7006 => x"26923878",
          7007 => x"81800a26",
          7008 => x"8b38ff19",
          7009 => x"79065574",
          7010 => x"802e8638",
          7011 => x"93568ae4",
          7012 => x"3978892a",
          7013 => x"6e892a70",
          7014 => x"892b7759",
          7015 => x"4843597a",
          7016 => x"83388156",
          7017 => x"61307080",
          7018 => x"25770751",
          7019 => x"55915674",
          7020 => x"8ac23899",
          7021 => x"3df80553",
          7022 => x"81527e51",
          7023 => x"ffa4813f",
          7024 => x"81568287",
          7025 => x"cc088aac",
          7026 => x"3877832a",
          7027 => x"70770682",
          7028 => x"87cc0843",
          7029 => x"56457483",
          7030 => x"38bf4166",
          7031 => x"558e5660",
          7032 => x"75268a90",
          7033 => x"38746131",
          7034 => x"70485580",
          7035 => x"ff75278a",
          7036 => x"83389356",
          7037 => x"78818026",
          7038 => x"89fa3877",
          7039 => x"812a7081",
          7040 => x"06564374",
          7041 => x"802e9538",
          7042 => x"77870655",
          7043 => x"74822e83",
          7044 => x"8d387781",
          7045 => x"06557480",
          7046 => x"2e838338",
          7047 => x"77810655",
          7048 => x"9356825e",
          7049 => x"74802e89",
          7050 => x"cb38785a",
          7051 => x"7d832e09",
          7052 => x"810680e1",
          7053 => x"3878ae38",
          7054 => x"66912a57",
          7055 => x"810b8282",
          7056 => x"b822565a",
          7057 => x"74802e9d",
          7058 => x"38747726",
          7059 => x"98388282",
          7060 => x"b8567910",
          7061 => x"82177022",
          7062 => x"57575a74",
          7063 => x"802e8638",
          7064 => x"767527ee",
          7065 => x"38795266",
          7066 => x"51ff8eff",
          7067 => x"3f8287cc",
          7068 => x"08842984",
          7069 => x"87057089",
          7070 => x"2a5e55a0",
          7071 => x"5c800b82",
          7072 => x"87cc08fc",
          7073 => x"808a0556",
          7074 => x"44fdfff0",
          7075 => x"0a752780",
          7076 => x"ec3888d3",
          7077 => x"3978ae38",
          7078 => x"668c2a57",
          7079 => x"810b8282",
          7080 => x"a822565a",
          7081 => x"74802e9d",
          7082 => x"38747726",
          7083 => x"98388282",
          7084 => x"a8567910",
          7085 => x"82177022",
          7086 => x"57575a74",
          7087 => x"802e8638",
          7088 => x"767527ee",
          7089 => x"38795266",
          7090 => x"51ff8e9f",
          7091 => x"3f8287cc",
          7092 => x"08108405",
          7093 => x"578287cc",
          7094 => x"089ff526",
          7095 => x"9638810b",
          7096 => x"8287cc08",
          7097 => x"108287cc",
          7098 => x"08057111",
          7099 => x"722a8305",
          7100 => x"59565e83",
          7101 => x"ff17892a",
          7102 => x"5d815ca0",
          7103 => x"44601c7d",
          7104 => x"11650569",
          7105 => x"7012ff05",
          7106 => x"71307072",
          7107 => x"0674315c",
          7108 => x"52595759",
          7109 => x"407d832e",
          7110 => x"09810689",
          7111 => x"38761c60",
          7112 => x"18415c84",
          7113 => x"39761d5d",
          7114 => x"79902918",
          7115 => x"70623168",
          7116 => x"58515574",
          7117 => x"762687af",
          7118 => x"38757c31",
          7119 => x"7d317a53",
          7120 => x"70653152",
          7121 => x"55ff8da3",
          7122 => x"3f8287cc",
          7123 => x"08587d83",
          7124 => x"2e098106",
          7125 => x"9b388287",
          7126 => x"cc0883ff",
          7127 => x"f52680dd",
          7128 => x"38788783",
          7129 => x"3879812a",
          7130 => x"5978fdbe",
          7131 => x"3886f839",
          7132 => x"7d822e09",
          7133 => x"810680c5",
          7134 => x"3883fff5",
          7135 => x"0b8287cc",
          7136 => x"0827a038",
          7137 => x"788f3879",
          7138 => x"1a557480",
          7139 => x"c0268638",
          7140 => x"7459fd96",
          7141 => x"39628106",
          7142 => x"5574802e",
          7143 => x"8f38835e",
          7144 => x"fd883982",
          7145 => x"87cc089f",
          7146 => x"f5269238",
          7147 => x"7886b838",
          7148 => x"791a5981",
          7149 => x"807927fc",
          7150 => x"f13886ab",
          7151 => x"3980557d",
          7152 => x"812e0981",
          7153 => x"0683387d",
          7154 => x"559ff578",
          7155 => x"278b3874",
          7156 => x"8106558e",
          7157 => x"5674869c",
          7158 => x"38848053",
          7159 => x"80527a51",
          7160 => x"ffa2ba3f",
          7161 => x"8b538280",
          7162 => x"d0527a51",
          7163 => x"ffa28b3f",
          7164 => x"8480528b",
          7165 => x"1b51ffa1",
          7166 => x"b43f798d",
          7167 => x"1c347b83",
          7168 => x"ffff0652",
          7169 => x"8e1b51ff",
          7170 => x"a1a33f81",
          7171 => x"0b901c34",
          7172 => x"7d833270",
          7173 => x"3070962a",
          7174 => x"84800654",
          7175 => x"5155911b",
          7176 => x"51ffa189",
          7177 => x"3f665574",
          7178 => x"83ffff26",
          7179 => x"90387483",
          7180 => x"ffff0652",
          7181 => x"931b51ff",
          7182 => x"a0f33f8a",
          7183 => x"397452a0",
          7184 => x"1b51ffa1",
          7185 => x"863ff80b",
          7186 => x"951c34bf",
          7187 => x"52981b51",
          7188 => x"ffa0da3f",
          7189 => x"81ff529a",
          7190 => x"1b51ffa0",
          7191 => x"d03f6052",
          7192 => x"9c1b51ff",
          7193 => x"a0e53f7d",
          7194 => x"832e0981",
          7195 => x"0680cb38",
          7196 => x"8288b20a",
          7197 => x"5280c31b",
          7198 => x"51ffa0cf",
          7199 => x"3f7c52a4",
          7200 => x"1b51ffa0",
          7201 => x"c63f8252",
          7202 => x"ac1b51ff",
          7203 => x"a0bd3f81",
          7204 => x"52b01b51",
          7205 => x"ffa0963f",
          7206 => x"8652b21b",
          7207 => x"51ffa08d",
          7208 => x"3fff800b",
          7209 => x"80c01c34",
          7210 => x"a90b80c2",
          7211 => x"1c349353",
          7212 => x"8280dc52",
          7213 => x"80c71b51",
          7214 => x"ae398288",
          7215 => x"b20a52a7",
          7216 => x"1b51ffa0",
          7217 => x"863f7c83",
          7218 => x"ffff0652",
          7219 => x"961b51ff",
          7220 => x"9fdb3fff",
          7221 => x"800ba41c",
          7222 => x"34a90ba6",
          7223 => x"1c349353",
          7224 => x"8280f052",
          7225 => x"ab1b51ff",
          7226 => x"a0903f82",
          7227 => x"d4d55283",
          7228 => x"fe1b7052",
          7229 => x"59ff9fb5",
          7230 => x"3f815460",
          7231 => x"537a527e",
          7232 => x"51ff9bd8",
          7233 => x"3f815682",
          7234 => x"87cc0883",
          7235 => x"e7387d83",
          7236 => x"2e098106",
          7237 => x"80ee3875",
          7238 => x"54608605",
          7239 => x"537a527e",
          7240 => x"51ff9bb8",
          7241 => x"3f848053",
          7242 => x"80527a51",
          7243 => x"ff9fee3f",
          7244 => x"848b85a4",
          7245 => x"d2527a51",
          7246 => x"ff9f903f",
          7247 => x"868a85e4",
          7248 => x"f25283e4",
          7249 => x"1b51ff9f",
          7250 => x"823fff18",
          7251 => x"5283e81b",
          7252 => x"51ff9ef7",
          7253 => x"3f825283",
          7254 => x"ec1b51ff",
          7255 => x"9eed3f82",
          7256 => x"d4d55278",
          7257 => x"51ff9ec5",
          7258 => x"3f755460",
          7259 => x"8705537a",
          7260 => x"527e51ff",
          7261 => x"9ae63f75",
          7262 => x"54601653",
          7263 => x"7a527e51",
          7264 => x"ff9ad93f",
          7265 => x"65538052",
          7266 => x"7a51ff9f",
          7267 => x"903f7f56",
          7268 => x"80587d83",
          7269 => x"2e098106",
          7270 => x"9a38f852",
          7271 => x"7a51ff9e",
          7272 => x"aa3fff52",
          7273 => x"841b51ff",
          7274 => x"9ea13ff0",
          7275 => x"0a52881b",
          7276 => x"51913987",
          7277 => x"fffff855",
          7278 => x"7d812e83",
          7279 => x"38f85574",
          7280 => x"527a51ff",
          7281 => x"9e853f7c",
          7282 => x"55615774",
          7283 => x"62268338",
          7284 => x"74577654",
          7285 => x"75537a52",
          7286 => x"7e51ff99",
          7287 => x"ff3f8287",
          7288 => x"cc088287",
          7289 => x"38848053",
          7290 => x"8287cc08",
          7291 => x"527a51ff",
          7292 => x"9eab3f76",
          7293 => x"16757831",
          7294 => x"565674cd",
          7295 => x"38811858",
          7296 => x"77802eff",
          7297 => x"8d387955",
          7298 => x"7d832e83",
          7299 => x"38635561",
          7300 => x"57746226",
          7301 => x"83387457",
          7302 => x"76547553",
          7303 => x"7a527e51",
          7304 => x"ff99b93f",
          7305 => x"8287cc08",
          7306 => x"81c13876",
          7307 => x"16757831",
          7308 => x"565674db",
          7309 => x"388c567d",
          7310 => x"832e9338",
          7311 => x"86566683",
          7312 => x"ffff268a",
          7313 => x"3884567d",
          7314 => x"822e8338",
          7315 => x"81566481",
          7316 => x"06587780",
          7317 => x"fe388480",
          7318 => x"5377527a",
          7319 => x"51ff9dbd",
          7320 => x"3f82d4d5",
          7321 => x"527851ff",
          7322 => x"9cc33f83",
          7323 => x"be1b5577",
          7324 => x"7534810b",
          7325 => x"81163481",
          7326 => x"0b821634",
          7327 => x"77831634",
          7328 => x"75841634",
          7329 => x"60670556",
          7330 => x"80fdc152",
          7331 => x"7551ff86",
          7332 => x"da3ffe0b",
          7333 => x"85163482",
          7334 => x"87cc0882",
          7335 => x"2abf0756",
          7336 => x"75861634",
          7337 => x"8287cc08",
          7338 => x"87163460",
          7339 => x"5283c61b",
          7340 => x"51ff9c97",
          7341 => x"3f665283",
          7342 => x"ca1b51ff",
          7343 => x"9c8d3f81",
          7344 => x"5477537a",
          7345 => x"527e51ff",
          7346 => x"98923f81",
          7347 => x"568287cc",
          7348 => x"08a23880",
          7349 => x"5380527e",
          7350 => x"51ff99e4",
          7351 => x"3f815682",
          7352 => x"87cc0890",
          7353 => x"3889398e",
          7354 => x"568a3981",
          7355 => x"56863982",
          7356 => x"87cc0856",
          7357 => x"758287cc",
          7358 => x"0c993d0d",
          7359 => x"04f53d0d",
          7360 => x"7d605b59",
          7361 => x"807960ff",
          7362 => x"055a5757",
          7363 => x"767825b4",
          7364 => x"388d3df8",
          7365 => x"11555581",
          7366 => x"53fc1552",
          7367 => x"7951c9dc",
          7368 => x"3f7a812e",
          7369 => x"0981069c",
          7370 => x"388c3d33",
          7371 => x"55748d2e",
          7372 => x"db387476",
          7373 => x"70810558",
          7374 => x"34811757",
          7375 => x"748a2e09",
          7376 => x"8106c938",
          7377 => x"80763478",
          7378 => x"55768338",
          7379 => x"76557482",
          7380 => x"87cc0c8d",
          7381 => x"3d0d04f7",
          7382 => x"3d0d7b02",
          7383 => x"8405b305",
          7384 => x"33595777",
          7385 => x"8a2e0981",
          7386 => x"0687388d",
          7387 => x"527651e7",
          7388 => x"3f841708",
          7389 => x"56807624",
          7390 => x"be388817",
          7391 => x"0877178c",
          7392 => x"05565977",
          7393 => x"75348116",
          7394 => x"56bb7625",
          7395 => x"a1388b3d",
          7396 => x"fc055475",
          7397 => x"538c1752",
          7398 => x"760851cb",
          7399 => x"dc3f7976",
          7400 => x"32703070",
          7401 => x"72079f2a",
          7402 => x"70305351",
          7403 => x"56567584",
          7404 => x"180c8119",
          7405 => x"88180c8b",
          7406 => x"3d0d04f9",
          7407 => x"3d0d7984",
          7408 => x"11085656",
          7409 => x"807524a7",
          7410 => x"38893dfc",
          7411 => x"05547453",
          7412 => x"8c165275",
          7413 => x"0851cba1",
          7414 => x"3f8287cc",
          7415 => x"08913884",
          7416 => x"1608782e",
          7417 => x"09810687",
          7418 => x"38881608",
          7419 => x"558339ff",
          7420 => x"55748287",
          7421 => x"cc0c893d",
          7422 => x"0d04fd3d",
          7423 => x"0d755480",
          7424 => x"cc538052",
          7425 => x"7351ff9a",
          7426 => x"943f7674",
          7427 => x"0c853d0d",
          7428 => x"04ea3d0d",
          7429 => x"0280e305",
          7430 => x"336a5386",
          7431 => x"3d705354",
          7432 => x"54d83f73",
          7433 => x"527251fe",
          7434 => x"ae3f7251",
          7435 => x"ff8d3f98",
          7436 => x"3d0d0400",
          7437 => x"00ffffff",
          7438 => x"ff00ffff",
          7439 => x"ffff00ff",
          7440 => x"ffffff00",
          7441 => x"00000e06",
          7442 => x"00000d8a",
          7443 => x"00000d91",
          7444 => x"00000d98",
          7445 => x"00000d9f",
          7446 => x"00000da6",
          7447 => x"00000dad",
          7448 => x"00000db4",
          7449 => x"00000dbb",
          7450 => x"00000dc2",
          7451 => x"00000dc9",
          7452 => x"00000dd0",
          7453 => x"00000dd6",
          7454 => x"00000ddc",
          7455 => x"00000de2",
          7456 => x"00000de8",
          7457 => x"00000dee",
          7458 => x"00000df4",
          7459 => x"00000dfa",
          7460 => x"00000e00",
          7461 => x"00002542",
          7462 => x"00002548",
          7463 => x"0000254e",
          7464 => x"00002554",
          7465 => x"0000255a",
          7466 => x"0000317c",
          7467 => x"00003270",
          7468 => x"00003363",
          7469 => x"00003597",
          7470 => x"00003258",
          7471 => x"00003051",
          7472 => x"00003413",
          7473 => x"0000356e",
          7474 => x"00003450",
          7475 => x"000034e6",
          7476 => x"0000346c",
          7477 => x"00003313",
          7478 => x"00003051",
          7479 => x"00003363",
          7480 => x"00003386",
          7481 => x"00003413",
          7482 => x"00003051",
          7483 => x"00003051",
          7484 => x"0000346c",
          7485 => x"000034e6",
          7486 => x"0000356e",
          7487 => x"00003597",
          7488 => x"64696e69",
          7489 => x"74000000",
          7490 => x"64696f63",
          7491 => x"746c0000",
          7492 => x"66696e69",
          7493 => x"74000000",
          7494 => x"666c6f61",
          7495 => x"64000000",
          7496 => x"66657865",
          7497 => x"63000000",
          7498 => x"6d636c65",
          7499 => x"61720000",
          7500 => x"6d636f70",
          7501 => x"79000000",
          7502 => x"6d646966",
          7503 => x"66000000",
          7504 => x"6d64756d",
          7505 => x"70000000",
          7506 => x"6d656200",
          7507 => x"6d656800",
          7508 => x"6d657700",
          7509 => x"68696400",
          7510 => x"68696500",
          7511 => x"68666400",
          7512 => x"68666500",
          7513 => x"63616c6c",
          7514 => x"00000000",
          7515 => x"6a6d7000",
          7516 => x"72657374",
          7517 => x"61727400",
          7518 => x"72657365",
          7519 => x"74000000",
          7520 => x"696e666f",
          7521 => x"00000000",
          7522 => x"74657374",
          7523 => x"00000000",
          7524 => x"74626173",
          7525 => x"69630000",
          7526 => x"6d626173",
          7527 => x"69630000",
          7528 => x"6b696c6f",
          7529 => x"00000000",
          7530 => x"65640000",
          7531 => x"4469736b",
          7532 => x"20457272",
          7533 => x"6f720a00",
          7534 => x"496e7465",
          7535 => x"726e616c",
          7536 => x"20657272",
          7537 => x"6f722e0a",
          7538 => x"00000000",
          7539 => x"4469736b",
          7540 => x"206e6f74",
          7541 => x"20726561",
          7542 => x"64792e0a",
          7543 => x"00000000",
          7544 => x"4e6f2066",
          7545 => x"696c6520",
          7546 => x"666f756e",
          7547 => x"642e0a00",
          7548 => x"4e6f2070",
          7549 => x"61746820",
          7550 => x"666f756e",
          7551 => x"642e0a00",
          7552 => x"496e7661",
          7553 => x"6c696420",
          7554 => x"66696c65",
          7555 => x"6e616d65",
          7556 => x"2e0a0000",
          7557 => x"41636365",
          7558 => x"73732064",
          7559 => x"656e6965",
          7560 => x"642e0a00",
          7561 => x"46696c65",
          7562 => x"20616c72",
          7563 => x"65616479",
          7564 => x"20657869",
          7565 => x"7374732e",
          7566 => x"0a000000",
          7567 => x"46696c65",
          7568 => x"2068616e",
          7569 => x"646c6520",
          7570 => x"696e7661",
          7571 => x"6c69642e",
          7572 => x"0a000000",
          7573 => x"53442069",
          7574 => x"73207772",
          7575 => x"69746520",
          7576 => x"70726f74",
          7577 => x"65637465",
          7578 => x"642e0a00",
          7579 => x"44726976",
          7580 => x"65206e75",
          7581 => x"6d626572",
          7582 => x"20697320",
          7583 => x"696e7661",
          7584 => x"6c69642e",
          7585 => x"0a000000",
          7586 => x"4469736b",
          7587 => x"206e6f74",
          7588 => x"20656e61",
          7589 => x"626c6564",
          7590 => x"2e0a0000",
          7591 => x"4e6f2063",
          7592 => x"6f6d7061",
          7593 => x"7469626c",
          7594 => x"65206669",
          7595 => x"6c657379",
          7596 => x"7374656d",
          7597 => x"20666f75",
          7598 => x"6e64206f",
          7599 => x"6e206469",
          7600 => x"736b2e0a",
          7601 => x"00000000",
          7602 => x"466f726d",
          7603 => x"61742061",
          7604 => x"626f7274",
          7605 => x"65642e0a",
          7606 => x"00000000",
          7607 => x"54696d65",
          7608 => x"6f75742c",
          7609 => x"206f7065",
          7610 => x"72617469",
          7611 => x"6f6e2063",
          7612 => x"616e6365",
          7613 => x"6c6c6564",
          7614 => x"2e0a0000",
          7615 => x"46696c65",
          7616 => x"20697320",
          7617 => x"6c6f636b",
          7618 => x"65642e0a",
          7619 => x"00000000",
          7620 => x"496e7375",
          7621 => x"66666963",
          7622 => x"69656e74",
          7623 => x"206d656d",
          7624 => x"6f72792e",
          7625 => x"0a000000",
          7626 => x"546f6f20",
          7627 => x"6d616e79",
          7628 => x"206f7065",
          7629 => x"6e206669",
          7630 => x"6c65732e",
          7631 => x"0a000000",
          7632 => x"50617261",
          7633 => x"6d657465",
          7634 => x"72732069",
          7635 => x"6e636f72",
          7636 => x"72656374",
          7637 => x"2e0a0000",
          7638 => x"53756363",
          7639 => x"6573732e",
          7640 => x"0a000000",
          7641 => x"556e6b6e",
          7642 => x"6f776e20",
          7643 => x"6572726f",
          7644 => x"722e0a00",
          7645 => x"0a256c75",
          7646 => x"20627974",
          7647 => x"65732025",
          7648 => x"73206174",
          7649 => x"20256c75",
          7650 => x"20627974",
          7651 => x"65732f73",
          7652 => x"65632e0a",
          7653 => x"00000000",
          7654 => x"72656164",
          7655 => x"00000000",
          7656 => x"25303858",
          7657 => x"00000000",
          7658 => x"3a202000",
          7659 => x"25303458",
          7660 => x"00000000",
          7661 => x"20202020",
          7662 => x"20202020",
          7663 => x"00000000",
          7664 => x"25303258",
          7665 => x"00000000",
          7666 => x"20200000",
          7667 => x"207c0000",
          7668 => x"7c0d0a00",
          7669 => x"5a505554",
          7670 => x"41000000",
          7671 => x"0a2a2a20",
          7672 => x"25732028",
          7673 => x"00000000",
          7674 => x"30322f30",
          7675 => x"352f3230",
          7676 => x"32300000",
          7677 => x"76312e35",
          7678 => x"32000000",
          7679 => x"205a5055",
          7680 => x"2c207265",
          7681 => x"76202530",
          7682 => x"32782920",
          7683 => x"25732025",
          7684 => x"73202a2a",
          7685 => x"0a0a0000",
          7686 => x"5a505554",
          7687 => x"4120496e",
          7688 => x"74657272",
          7689 => x"75707420",
          7690 => x"48616e64",
          7691 => x"6c65720a",
          7692 => x"00000000",
          7693 => x"54696d65",
          7694 => x"7220696e",
          7695 => x"74657272",
          7696 => x"7570740a",
          7697 => x"00000000",
          7698 => x"50533220",
          7699 => x"696e7465",
          7700 => x"72727570",
          7701 => x"740a0000",
          7702 => x"494f4354",
          7703 => x"4c205244",
          7704 => x"20696e74",
          7705 => x"65727275",
          7706 => x"70740a00",
          7707 => x"494f4354",
          7708 => x"4c205752",
          7709 => x"20696e74",
          7710 => x"65727275",
          7711 => x"70740a00",
          7712 => x"55415254",
          7713 => x"30205258",
          7714 => x"20696e74",
          7715 => x"65727275",
          7716 => x"70740a00",
          7717 => x"55415254",
          7718 => x"30205458",
          7719 => x"20696e74",
          7720 => x"65727275",
          7721 => x"70740a00",
          7722 => x"55415254",
          7723 => x"31205258",
          7724 => x"20696e74",
          7725 => x"65727275",
          7726 => x"70740a00",
          7727 => x"55415254",
          7728 => x"31205458",
          7729 => x"20696e74",
          7730 => x"65727275",
          7731 => x"70740a00",
          7732 => x"53657474",
          7733 => x"696e6720",
          7734 => x"75702074",
          7735 => x"696d6572",
          7736 => x"2e2e2e0a",
          7737 => x"00000000",
          7738 => x"456e6162",
          7739 => x"6c696e67",
          7740 => x"2074696d",
          7741 => x"65722e2e",
          7742 => x"2e0a0000",
          7743 => x"6175746f",
          7744 => x"65786563",
          7745 => x"2e626174",
          7746 => x"00000000",
          7747 => x"7a707574",
          7748 => x"612e6873",
          7749 => x"74000000",
          7750 => x"303a0000",
          7751 => x"4661696c",
          7752 => x"65642074",
          7753 => x"6f20696e",
          7754 => x"69746961",
          7755 => x"6c697365",
          7756 => x"20736420",
          7757 => x"63617264",
          7758 => x"20302c20",
          7759 => x"706c6561",
          7760 => x"73652069",
          7761 => x"6e697420",
          7762 => x"6d616e75",
          7763 => x"616c6c79",
          7764 => x"2e0a0000",
          7765 => x"2a200000",
          7766 => x"42616420",
          7767 => x"6469736b",
          7768 => x"20696421",
          7769 => x"0a000000",
          7770 => x"496e6974",
          7771 => x"69616c69",
          7772 => x"7365642e",
          7773 => x"0a000000",
          7774 => x"4661696c",
          7775 => x"65642074",
          7776 => x"6f20696e",
          7777 => x"69746961",
          7778 => x"6c697365",
          7779 => x"2e0a0000",
          7780 => x"72633d25",
          7781 => x"640a0000",
          7782 => x"25753a00",
          7783 => x"436c6561",
          7784 => x"72696e67",
          7785 => x"2e2e2e2e",
          7786 => x"00000000",
          7787 => x"436f7079",
          7788 => x"696e672e",
          7789 => x"2e2e0000",
          7790 => x"436f6d70",
          7791 => x"6172696e",
          7792 => x"672e2e2e",
          7793 => x"00000000",
          7794 => x"2530386c",
          7795 => x"78282530",
          7796 => x"3878292d",
          7797 => x"3e253038",
          7798 => x"6c782825",
          7799 => x"30387829",
          7800 => x"0a000000",
          7801 => x"44756d70",
          7802 => x"204d656d",
          7803 => x"6f72790a",
          7804 => x"00000000",
          7805 => x"0a436f6d",
          7806 => x"706c6574",
          7807 => x"652e0a00",
          7808 => x"25303858",
          7809 => x"20253032",
          7810 => x"582d0000",
          7811 => x"3f3f3f0a",
          7812 => x"00000000",
          7813 => x"25303858",
          7814 => x"20253034",
          7815 => x"582d0000",
          7816 => x"25303858",
          7817 => x"20253038",
          7818 => x"582d0000",
          7819 => x"44697361",
          7820 => x"626c696e",
          7821 => x"6720696e",
          7822 => x"74657272",
          7823 => x"75707473",
          7824 => x"0a000000",
          7825 => x"456e6162",
          7826 => x"6c696e67",
          7827 => x"20696e74",
          7828 => x"65727275",
          7829 => x"7074730a",
          7830 => x"00000000",
          7831 => x"44697361",
          7832 => x"626c6564",
          7833 => x"20756172",
          7834 => x"74206669",
          7835 => x"666f0a00",
          7836 => x"456e6162",
          7837 => x"6c696e67",
          7838 => x"20756172",
          7839 => x"74206669",
          7840 => x"666f0a00",
          7841 => x"45786563",
          7842 => x"7574696e",
          7843 => x"6720636f",
          7844 => x"64652040",
          7845 => x"20253038",
          7846 => x"78202e2e",
          7847 => x"2e0a0000",
          7848 => x"43616c6c",
          7849 => x"696e6720",
          7850 => x"636f6465",
          7851 => x"20402025",
          7852 => x"30387820",
          7853 => x"2e2e2e0a",
          7854 => x"00000000",
          7855 => x"43616c6c",
          7856 => x"20726574",
          7857 => x"75726e65",
          7858 => x"6420636f",
          7859 => x"64652028",
          7860 => x"2564292e",
          7861 => x"0a000000",
          7862 => x"52657374",
          7863 => x"61727469",
          7864 => x"6e672061",
          7865 => x"70706c69",
          7866 => x"63617469",
          7867 => x"6f6e2e2e",
          7868 => x"2e0a0000",
          7869 => x"436f6c64",
          7870 => x"20726562",
          7871 => x"6f6f7469",
          7872 => x"6e672e2e",
          7873 => x"2e0a0000",
          7874 => x"5a505500",
          7875 => x"62696e00",
          7876 => x"25643a5c",
          7877 => x"25735c25",
          7878 => x"732e2573",
          7879 => x"00000000",
          7880 => x"25643a5c",
          7881 => x"25735c25",
          7882 => x"73000000",
          7883 => x"25643a5c",
          7884 => x"25730000",
          7885 => x"42616420",
          7886 => x"636f6d6d",
          7887 => x"616e642e",
          7888 => x"0a000000",
          7889 => x"52756e6e",
          7890 => x"696e672e",
          7891 => x"2e2e0a00",
          7892 => x"456e6162",
          7893 => x"6c696e67",
          7894 => x"20696e74",
          7895 => x"65727275",
          7896 => x"7074732e",
          7897 => x"2e2e0a00",
          7898 => x"25642f25",
          7899 => x"642f2564",
          7900 => x"2025643a",
          7901 => x"25643a25",
          7902 => x"642e2564",
          7903 => x"25640a00",
          7904 => x"536f4320",
          7905 => x"436f6e66",
          7906 => x"69677572",
          7907 => x"6174696f",
          7908 => x"6e000000",
          7909 => x"20286672",
          7910 => x"6f6d2053",
          7911 => x"6f432063",
          7912 => x"6f6e6669",
          7913 => x"67290000",
          7914 => x"3a0a4465",
          7915 => x"76696365",
          7916 => x"7320696d",
          7917 => x"706c656d",
          7918 => x"656e7465",
          7919 => x"643a0a00",
          7920 => x"20202020",
          7921 => x"57422053",
          7922 => x"4452414d",
          7923 => x"20202825",
          7924 => x"3038583a",
          7925 => x"25303858",
          7926 => x"292e0a00",
          7927 => x"20202020",
          7928 => x"53445241",
          7929 => x"4d202020",
          7930 => x"20202825",
          7931 => x"3038583a",
          7932 => x"25303858",
          7933 => x"292e0a00",
          7934 => x"20202020",
          7935 => x"494e534e",
          7936 => x"20425241",
          7937 => x"4d202825",
          7938 => x"3038583a",
          7939 => x"25303858",
          7940 => x"292e0a00",
          7941 => x"20202020",
          7942 => x"4252414d",
          7943 => x"20202020",
          7944 => x"20202825",
          7945 => x"3038583a",
          7946 => x"25303858",
          7947 => x"292e0a00",
          7948 => x"20202020",
          7949 => x"52414d20",
          7950 => x"20202020",
          7951 => x"20202825",
          7952 => x"3038583a",
          7953 => x"25303858",
          7954 => x"292e0a00",
          7955 => x"20202020",
          7956 => x"53442043",
          7957 => x"41524420",
          7958 => x"20202844",
          7959 => x"65766963",
          7960 => x"6573203d",
          7961 => x"25303264",
          7962 => x"292e0a00",
          7963 => x"20202020",
          7964 => x"54494d45",
          7965 => x"52312020",
          7966 => x"20202854",
          7967 => x"696d6572",
          7968 => x"7320203d",
          7969 => x"25303264",
          7970 => x"292e0a00",
          7971 => x"20202020",
          7972 => x"494e5452",
          7973 => x"20435452",
          7974 => x"4c202843",
          7975 => x"68616e6e",
          7976 => x"656c733d",
          7977 => x"25303264",
          7978 => x"292e0a00",
          7979 => x"20202020",
          7980 => x"57495348",
          7981 => x"424f4e45",
          7982 => x"20425553",
          7983 => x"0a000000",
          7984 => x"20202020",
          7985 => x"57422049",
          7986 => x"32430a00",
          7987 => x"20202020",
          7988 => x"494f4354",
          7989 => x"4c0a0000",
          7990 => x"20202020",
          7991 => x"5053320a",
          7992 => x"00000000",
          7993 => x"20202020",
          7994 => x"5350490a",
          7995 => x"00000000",
          7996 => x"41646472",
          7997 => x"65737365",
          7998 => x"733a0a00",
          7999 => x"20202020",
          8000 => x"43505520",
          8001 => x"52657365",
          8002 => x"74205665",
          8003 => x"63746f72",
          8004 => x"20416464",
          8005 => x"72657373",
          8006 => x"203d2025",
          8007 => x"3038580a",
          8008 => x"00000000",
          8009 => x"20202020",
          8010 => x"43505520",
          8011 => x"4d656d6f",
          8012 => x"72792053",
          8013 => x"74617274",
          8014 => x"20416464",
          8015 => x"72657373",
          8016 => x"203d2025",
          8017 => x"3038580a",
          8018 => x"00000000",
          8019 => x"20202020",
          8020 => x"53746163",
          8021 => x"6b205374",
          8022 => x"61727420",
          8023 => x"41646472",
          8024 => x"65737320",
          8025 => x"20202020",
          8026 => x"203d2025",
          8027 => x"3038580a",
          8028 => x"00000000",
          8029 => x"4d697363",
          8030 => x"3a0a0000",
          8031 => x"20202020",
          8032 => x"5a505520",
          8033 => x"49642020",
          8034 => x"20202020",
          8035 => x"20202020",
          8036 => x"20202020",
          8037 => x"20202020",
          8038 => x"203d2025",
          8039 => x"3034580a",
          8040 => x"00000000",
          8041 => x"20202020",
          8042 => x"53797374",
          8043 => x"656d2043",
          8044 => x"6c6f636b",
          8045 => x"20467265",
          8046 => x"71202020",
          8047 => x"20202020",
          8048 => x"203d2025",
          8049 => x"642e2530",
          8050 => x"34644d48",
          8051 => x"7a0a0000",
          8052 => x"20202020",
          8053 => x"53445241",
          8054 => x"4d20436c",
          8055 => x"6f636b20",
          8056 => x"46726571",
          8057 => x"20202020",
          8058 => x"20202020",
          8059 => x"203d2025",
          8060 => x"642e2530",
          8061 => x"34644d48",
          8062 => x"7a0a0000",
          8063 => x"20202020",
          8064 => x"57697368",
          8065 => x"626f6e65",
          8066 => x"20534452",
          8067 => x"414d2043",
          8068 => x"6c6f636b",
          8069 => x"20467265",
          8070 => x"713d2025",
          8071 => x"642e2530",
          8072 => x"34644d48",
          8073 => x"7a0a0000",
          8074 => x"536d616c",
          8075 => x"6c000000",
          8076 => x"4d656469",
          8077 => x"756d0000",
          8078 => x"466c6578",
          8079 => x"00000000",
          8080 => x"45564f00",
          8081 => x"45564f6d",
          8082 => x"696e0000",
          8083 => x"556e6b6e",
          8084 => x"6f776e00",
          8085 => x"00007fb0",
          8086 => x"01000000",
          8087 => x"00000002",
          8088 => x"00007fac",
          8089 => x"01000000",
          8090 => x"00000003",
          8091 => x"00007fa8",
          8092 => x"01000000",
          8093 => x"00000004",
          8094 => x"00007fa4",
          8095 => x"01000000",
          8096 => x"00000005",
          8097 => x"00007fa0",
          8098 => x"01000000",
          8099 => x"00000006",
          8100 => x"00007f9c",
          8101 => x"01000000",
          8102 => x"00000007",
          8103 => x"00007f98",
          8104 => x"01000000",
          8105 => x"00000001",
          8106 => x"00007f94",
          8107 => x"01000000",
          8108 => x"00000008",
          8109 => x"00007f90",
          8110 => x"01000000",
          8111 => x"0000000b",
          8112 => x"00007f8c",
          8113 => x"01000000",
          8114 => x"00000009",
          8115 => x"00007f88",
          8116 => x"01000000",
          8117 => x"0000000a",
          8118 => x"00007f84",
          8119 => x"04000000",
          8120 => x"0000000d",
          8121 => x"00007f80",
          8122 => x"04000000",
          8123 => x"0000000c",
          8124 => x"00007f7c",
          8125 => x"04000000",
          8126 => x"0000000e",
          8127 => x"00007f78",
          8128 => x"03000000",
          8129 => x"0000000f",
          8130 => x"00007f74",
          8131 => x"04000000",
          8132 => x"0000000f",
          8133 => x"00007f70",
          8134 => x"04000000",
          8135 => x"00000010",
          8136 => x"00007f6c",
          8137 => x"04000000",
          8138 => x"00000011",
          8139 => x"00007f68",
          8140 => x"03000000",
          8141 => x"00000012",
          8142 => x"00007f64",
          8143 => x"03000000",
          8144 => x"00000013",
          8145 => x"00007f60",
          8146 => x"03000000",
          8147 => x"00000014",
          8148 => x"00007f5c",
          8149 => x"03000000",
          8150 => x"00000015",
          8151 => x"1b5b4400",
          8152 => x"1b5b4300",
          8153 => x"1b5b4200",
          8154 => x"1b5b4100",
          8155 => x"1b5b367e",
          8156 => x"1b5b357e",
          8157 => x"1b5b347e",
          8158 => x"1b304600",
          8159 => x"1b5b337e",
          8160 => x"1b5b327e",
          8161 => x"1b5b317e",
          8162 => x"10000000",
          8163 => x"0e000000",
          8164 => x"0d000000",
          8165 => x"0b000000",
          8166 => x"08000000",
          8167 => x"06000000",
          8168 => x"05000000",
          8169 => x"04000000",
          8170 => x"03000000",
          8171 => x"02000000",
          8172 => x"01000000",
          8173 => x"68697374",
          8174 => x"6f727900",
          8175 => x"68697374",
          8176 => x"00000000",
          8177 => x"21000000",
          8178 => x"25303464",
          8179 => x"20202573",
          8180 => x"0a000000",
          8181 => x"4661696c",
          8182 => x"65642074",
          8183 => x"6f207265",
          8184 => x"73657420",
          8185 => x"74686520",
          8186 => x"68697374",
          8187 => x"6f727920",
          8188 => x"66696c65",
          8189 => x"20746f20",
          8190 => x"454f462e",
          8191 => x"0a000000",
          8192 => x"43616e6e",
          8193 => x"6f74206f",
          8194 => x"70656e2f",
          8195 => x"63726561",
          8196 => x"74652068",
          8197 => x"6973746f",
          8198 => x"72792066",
          8199 => x"696c652c",
          8200 => x"20646973",
          8201 => x"61626c69",
          8202 => x"6e672e0a",
          8203 => x"00000000",
          8204 => x"53440000",
          8205 => x"222a2b2c",
          8206 => x"3a3b3c3d",
          8207 => x"3e3f5b5d",
          8208 => x"7c7f0000",
          8209 => x"46415400",
          8210 => x"46415433",
          8211 => x"32000000",
          8212 => x"ebfe904d",
          8213 => x"53444f53",
          8214 => x"352e3000",
          8215 => x"4e4f204e",
          8216 => x"414d4520",
          8217 => x"20202046",
          8218 => x"41543332",
          8219 => x"20202000",
          8220 => x"4e4f204e",
          8221 => x"414d4520",
          8222 => x"20202046",
          8223 => x"41542020",
          8224 => x"20202000",
          8225 => x"00008030",
          8226 => x"00000000",
          8227 => x"00000000",
          8228 => x"00000000",
          8229 => x"809a4541",
          8230 => x"8e418f80",
          8231 => x"45454549",
          8232 => x"49498e8f",
          8233 => x"9092924f",
          8234 => x"994f5555",
          8235 => x"59999a9b",
          8236 => x"9c9d9e9f",
          8237 => x"41494f55",
          8238 => x"a5a5a6a7",
          8239 => x"a8a9aaab",
          8240 => x"acadaeaf",
          8241 => x"b0b1b2b3",
          8242 => x"b4b5b6b7",
          8243 => x"b8b9babb",
          8244 => x"bcbdbebf",
          8245 => x"c0c1c2c3",
          8246 => x"c4c5c6c7",
          8247 => x"c8c9cacb",
          8248 => x"cccdcecf",
          8249 => x"d0d1d2d3",
          8250 => x"d4d5d6d7",
          8251 => x"d8d9dadb",
          8252 => x"dcdddedf",
          8253 => x"e0e1e2e3",
          8254 => x"e4e5e6e7",
          8255 => x"e8e9eaeb",
          8256 => x"ecedeeef",
          8257 => x"f0f1f2f3",
          8258 => x"f4f5f6f7",
          8259 => x"f8f9fafb",
          8260 => x"fcfdfeff",
          8261 => x"2b2e2c3b",
          8262 => x"3d5b5d2f",
          8263 => x"5c222a3a",
          8264 => x"3c3e3f7c",
          8265 => x"7f000000",
          8266 => x"00010004",
          8267 => x"00100040",
          8268 => x"01000200",
          8269 => x"00000000",
          8270 => x"00010002",
          8271 => x"00040008",
          8272 => x"00100020",
          8273 => x"00000000",
          8274 => x"00000000",
          8275 => x"00007500",
          8276 => x"01020100",
          8277 => x"00000000",
          8278 => x"00000000",
          8279 => x"00007508",
          8280 => x"01040100",
          8281 => x"00000000",
          8282 => x"00000000",
          8283 => x"00007510",
          8284 => x"01140300",
          8285 => x"00000000",
          8286 => x"00000000",
          8287 => x"00007518",
          8288 => x"012b0300",
          8289 => x"00000000",
          8290 => x"00000000",
          8291 => x"00007520",
          8292 => x"01300300",
          8293 => x"00000000",
          8294 => x"00000000",
          8295 => x"00007528",
          8296 => x"013c0400",
          8297 => x"00000000",
          8298 => x"00000000",
          8299 => x"00007530",
          8300 => x"013d0400",
          8301 => x"00000000",
          8302 => x"00000000",
          8303 => x"00007538",
          8304 => x"013f0400",
          8305 => x"00000000",
          8306 => x"00000000",
          8307 => x"00007540",
          8308 => x"01400400",
          8309 => x"00000000",
          8310 => x"00000000",
          8311 => x"00007548",
          8312 => x"01410400",
          8313 => x"00000000",
          8314 => x"00000000",
          8315 => x"0000754c",
          8316 => x"01420400",
          8317 => x"00000000",
          8318 => x"00000000",
          8319 => x"00007550",
          8320 => x"01430400",
          8321 => x"00000000",
          8322 => x"00000000",
          8323 => x"00007554",
          8324 => x"01500500",
          8325 => x"00000000",
          8326 => x"00000000",
          8327 => x"00007558",
          8328 => x"01510500",
          8329 => x"00000000",
          8330 => x"00000000",
          8331 => x"0000755c",
          8332 => x"01540500",
          8333 => x"00000000",
          8334 => x"00000000",
          8335 => x"00007560",
          8336 => x"01550500",
          8337 => x"00000000",
          8338 => x"00000000",
          8339 => x"00007564",
          8340 => x"01790700",
          8341 => x"00000000",
          8342 => x"00000000",
          8343 => x"0000756c",
          8344 => x"01780700",
          8345 => x"00000000",
          8346 => x"00000000",
          8347 => x"00007570",
          8348 => x"01820800",
          8349 => x"00000000",
          8350 => x"00000000",
          8351 => x"00007578",
          8352 => x"01830800",
          8353 => x"00000000",
          8354 => x"00000000",
          8355 => x"00007580",
          8356 => x"01850800",
          8357 => x"00000000",
          8358 => x"00000000",
          8359 => x"00007588",
          8360 => x"01870800",
          8361 => x"00000000",
          8362 => x"00000000",
          8363 => x"00007590",
          8364 => x"018c0900",
          8365 => x"00000000",
          8366 => x"00000000",
          8367 => x"00007598",
          8368 => x"018d0900",
          8369 => x"00000000",
          8370 => x"00000000",
          8371 => x"000075a0",
          8372 => x"018e0900",
          8373 => x"00000000",
          8374 => x"00000000",
          8375 => x"000075a8",
          8376 => x"018f0900",
          8377 => x"00000000",
          8378 => x"00000000",
          8379 => x"00000000",
          8380 => x"00000000",
          8381 => x"00007fff",
          8382 => x"00000000",
          8383 => x"00007fff",
          8384 => x"00010000",
          8385 => x"00007fff",
          8386 => x"00010000",
          8387 => x"00810000",
          8388 => x"01000000",
          8389 => x"017fffff",
          8390 => x"00000000",
          8391 => x"00000000",
          8392 => x"00007800",
          8393 => x"00000000",
          8394 => x"05f5e100",
          8395 => x"05f5e100",
          8396 => x"05f5e100",
          8397 => x"00000000",
          8398 => x"01010101",
          8399 => x"01010101",
          8400 => x"01011001",
          8401 => x"01000000",
          8402 => x"00000000",
          8403 => x"00000000",
          8404 => x"00000000",
          8405 => x"00000000",
          8406 => x"00000000",
          8407 => x"00000000",
          8408 => x"00000000",
          8409 => x"00000000",
          8410 => x"00000000",
          8411 => x"00000000",
          8412 => x"00000000",
          8413 => x"00000000",
          8414 => x"00000000",
          8415 => x"00000000",
          8416 => x"00000000",
          8417 => x"00000000",
          8418 => x"00000000",
          8419 => x"00000000",
          8420 => x"00000000",
          8421 => x"00000000",
          8422 => x"00000000",
          8423 => x"00000000",
          8424 => x"00000000",
          8425 => x"00000000",
          8426 => x"00007fb4",
          8427 => x"01000000",
          8428 => x"00007fbc",
          8429 => x"01000000",
          8430 => x"00007fc4",
          8431 => x"02000000",
          8432 => x"00000000",
          8433 => x"00000000",
          8434 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

